module bsg_mem_1rw_sync_mask_write_bit_synth_width_p7_els_p64
(
  clk_i,
  reset_i,
  data_i,
  addr_i,
  v_i,
  w_mask_i,
  w_i,
  data_o
);

  input [6:0] data_i;
  input [5:0] addr_i;
  input [6:0] w_mask_i;
  output [6:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input w_i;
  wire [6:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140;
  wire [5:0] addr_r;
  wire [447:0] mem;
  reg addr_r_5_sv2v_reg,addr_r_4_sv2v_reg,addr_r_3_sv2v_reg,addr_r_2_sv2v_reg,
  addr_r_1_sv2v_reg,addr_r_0_sv2v_reg,mem_447_sv2v_reg,mem_446_sv2v_reg,mem_445_sv2v_reg,
  mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,mem_441_sv2v_reg,
  mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,mem_436_sv2v_reg,
  mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,mem_431_sv2v_reg,
  mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,mem_427_sv2v_reg,
  mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,mem_422_sv2v_reg,
  mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,mem_417_sv2v_reg,
  mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,mem_413_sv2v_reg,mem_412_sv2v_reg,
  mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,mem_408_sv2v_reg,
  mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,mem_403_sv2v_reg,
  mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,mem_399_sv2v_reg,mem_398_sv2v_reg,
  mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,mem_394_sv2v_reg,
  mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,mem_389_sv2v_reg,
  mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,mem_384_sv2v_reg,
  mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,mem_380_sv2v_reg,
  mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,mem_375_sv2v_reg,
  mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,mem_370_sv2v_reg,
  mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,mem_366_sv2v_reg,mem_365_sv2v_reg,
  mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,mem_361_sv2v_reg,
  mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,mem_356_sv2v_reg,
  mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,mem_351_sv2v_reg,
  mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,mem_347_sv2v_reg,
  mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,mem_342_sv2v_reg,
  mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,mem_337_sv2v_reg,
  mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,mem_333_sv2v_reg,mem_332_sv2v_reg,
  mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,mem_328_sv2v_reg,
  mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,mem_323_sv2v_reg,
  mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,mem_319_sv2v_reg,mem_318_sv2v_reg,
  mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,mem_314_sv2v_reg,
  mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,mem_309_sv2v_reg,
  mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,mem_304_sv2v_reg,
  mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,mem_300_sv2v_reg,
  mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,mem_295_sv2v_reg,
  mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,mem_290_sv2v_reg,
  mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,mem_286_sv2v_reg,mem_285_sv2v_reg,
  mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,mem_281_sv2v_reg,
  mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,mem_276_sv2v_reg,
  mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,mem_271_sv2v_reg,
  mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,mem_267_sv2v_reg,
  mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,mem_262_sv2v_reg,
  mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,mem_257_sv2v_reg,
  mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,mem_253_sv2v_reg,mem_252_sv2v_reg,
  mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,mem_248_sv2v_reg,
  mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,mem_243_sv2v_reg,
  mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,mem_239_sv2v_reg,mem_238_sv2v_reg,
  mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,mem_234_sv2v_reg,
  mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,mem_229_sv2v_reg,
  mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,mem_224_sv2v_reg,
  mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,mem_220_sv2v_reg,
  mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,mem_215_sv2v_reg,
  mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,mem_210_sv2v_reg,
  mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,mem_206_sv2v_reg,mem_205_sv2v_reg,
  mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,mem_201_sv2v_reg,
  mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,mem_196_sv2v_reg,
  mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,mem_191_sv2v_reg,
  mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,mem_187_sv2v_reg,
  mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,mem_182_sv2v_reg,
  mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,mem_177_sv2v_reg,
  mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,mem_173_sv2v_reg,mem_172_sv2v_reg,
  mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,mem_168_sv2v_reg,
  mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,mem_163_sv2v_reg,
  mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,mem_159_sv2v_reg,mem_158_sv2v_reg,
  mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,mem_154_sv2v_reg,
  mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,mem_149_sv2v_reg,
  mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,mem_144_sv2v_reg,
  mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,mem_140_sv2v_reg,
  mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,mem_135_sv2v_reg,
  mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,mem_130_sv2v_reg,
  mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,mem_126_sv2v_reg,mem_125_sv2v_reg,
  mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,mem_121_sv2v_reg,
  mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,mem_116_sv2v_reg,
  mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,mem_111_sv2v_reg,
  mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,mem_107_sv2v_reg,
  mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,mem_102_sv2v_reg,
  mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,mem_97_sv2v_reg,
  mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,mem_92_sv2v_reg,
  mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,mem_87_sv2v_reg,
  mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,mem_82_sv2v_reg,
  mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,mem_77_sv2v_reg,
  mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,mem_72_sv2v_reg,
  mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,mem_67_sv2v_reg,
  mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,mem_62_sv2v_reg,
  mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,mem_57_sv2v_reg,
  mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,mem_52_sv2v_reg,
  mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,mem_47_sv2v_reg,
  mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,mem_42_sv2v_reg,
  mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,mem_37_sv2v_reg,
  mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,mem_32_sv2v_reg,
  mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,mem_27_sv2v_reg,
  mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,mem_22_sv2v_reg,
  mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,mem_17_sv2v_reg,
  mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,mem_12_sv2v_reg,
  mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,mem_7_sv2v_reg,
  mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,mem_2_sv2v_reg,mem_1_sv2v_reg,
  mem_0_sv2v_reg;
  assign addr_r[5] = addr_r_5_sv2v_reg;
  assign addr_r[4] = addr_r_4_sv2v_reg;
  assign addr_r[3] = addr_r_3_sv2v_reg;
  assign addr_r[2] = addr_r_2_sv2v_reg;
  assign addr_r[1] = addr_r_1_sv2v_reg;
  assign addr_r[0] = addr_r_0_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_5_sv2v_reg <= addr_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_4_sv2v_reg <= addr_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_3_sv2v_reg <= addr_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_2_sv2v_reg <= addr_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_1_sv2v_reg <= addr_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      addr_r_0_sv2v_reg <= addr_i[0];
    end 
  end

  assign data_o[6] = (N82)? mem[6] : 
                     (N84)? mem[13] : 
                     (N86)? mem[20] : 
                     (N88)? mem[27] : 
                     (N90)? mem[34] : 
                     (N92)? mem[41] : 
                     (N94)? mem[48] : 
                     (N96)? mem[55] : 
                     (N98)? mem[62] : 
                     (N100)? mem[69] : 
                     (N102)? mem[76] : 
                     (N104)? mem[83] : 
                     (N106)? mem[90] : 
                     (N108)? mem[97] : 
                     (N110)? mem[104] : 
                     (N112)? mem[111] : 
                     (N114)? mem[118] : 
                     (N116)? mem[125] : 
                     (N118)? mem[132] : 
                     (N120)? mem[139] : 
                     (N122)? mem[146] : 
                     (N124)? mem[153] : 
                     (N126)? mem[160] : 
                     (N128)? mem[167] : 
                     (N130)? mem[174] : 
                     (N132)? mem[181] : 
                     (N134)? mem[188] : 
                     (N136)? mem[195] : 
                     (N138)? mem[202] : 
                     (N140)? mem[209] : 
                     (N142)? mem[216] : 
                     (N144)? mem[223] : 
                     (N83)? mem[230] : 
                     (N85)? mem[237] : 
                     (N87)? mem[244] : 
                     (N89)? mem[251] : 
                     (N91)? mem[258] : 
                     (N93)? mem[265] : 
                     (N95)? mem[272] : 
                     (N97)? mem[279] : 
                     (N99)? mem[286] : 
                     (N101)? mem[293] : 
                     (N103)? mem[300] : 
                     (N105)? mem[307] : 
                     (N107)? mem[314] : 
                     (N109)? mem[321] : 
                     (N111)? mem[328] : 
                     (N113)? mem[335] : 
                     (N115)? mem[342] : 
                     (N117)? mem[349] : 
                     (N119)? mem[356] : 
                     (N121)? mem[363] : 
                     (N123)? mem[370] : 
                     (N125)? mem[377] : 
                     (N127)? mem[384] : 
                     (N129)? mem[391] : 
                     (N131)? mem[398] : 
                     (N133)? mem[405] : 
                     (N135)? mem[412] : 
                     (N137)? mem[419] : 
                     (N139)? mem[426] : 
                     (N141)? mem[433] : 
                     (N143)? mem[440] : 
                     (N145)? mem[447] : 1'b0;
  assign data_o[5] = (N82)? mem[5] : 
                     (N84)? mem[12] : 
                     (N86)? mem[19] : 
                     (N88)? mem[26] : 
                     (N90)? mem[33] : 
                     (N92)? mem[40] : 
                     (N94)? mem[47] : 
                     (N96)? mem[54] : 
                     (N98)? mem[61] : 
                     (N100)? mem[68] : 
                     (N102)? mem[75] : 
                     (N104)? mem[82] : 
                     (N106)? mem[89] : 
                     (N108)? mem[96] : 
                     (N110)? mem[103] : 
                     (N112)? mem[110] : 
                     (N114)? mem[117] : 
                     (N116)? mem[124] : 
                     (N118)? mem[131] : 
                     (N120)? mem[138] : 
                     (N122)? mem[145] : 
                     (N124)? mem[152] : 
                     (N126)? mem[159] : 
                     (N128)? mem[166] : 
                     (N130)? mem[173] : 
                     (N132)? mem[180] : 
                     (N134)? mem[187] : 
                     (N136)? mem[194] : 
                     (N138)? mem[201] : 
                     (N140)? mem[208] : 
                     (N142)? mem[215] : 
                     (N144)? mem[222] : 
                     (N83)? mem[229] : 
                     (N85)? mem[236] : 
                     (N87)? mem[243] : 
                     (N89)? mem[250] : 
                     (N91)? mem[257] : 
                     (N93)? mem[264] : 
                     (N95)? mem[271] : 
                     (N97)? mem[278] : 
                     (N99)? mem[285] : 
                     (N101)? mem[292] : 
                     (N103)? mem[299] : 
                     (N105)? mem[306] : 
                     (N107)? mem[313] : 
                     (N109)? mem[320] : 
                     (N111)? mem[327] : 
                     (N113)? mem[334] : 
                     (N115)? mem[341] : 
                     (N117)? mem[348] : 
                     (N119)? mem[355] : 
                     (N121)? mem[362] : 
                     (N123)? mem[369] : 
                     (N125)? mem[376] : 
                     (N127)? mem[383] : 
                     (N129)? mem[390] : 
                     (N131)? mem[397] : 
                     (N133)? mem[404] : 
                     (N135)? mem[411] : 
                     (N137)? mem[418] : 
                     (N139)? mem[425] : 
                     (N141)? mem[432] : 
                     (N143)? mem[439] : 
                     (N145)? mem[446] : 1'b0;
  assign data_o[4] = (N82)? mem[4] : 
                     (N84)? mem[11] : 
                     (N86)? mem[18] : 
                     (N88)? mem[25] : 
                     (N90)? mem[32] : 
                     (N92)? mem[39] : 
                     (N94)? mem[46] : 
                     (N96)? mem[53] : 
                     (N98)? mem[60] : 
                     (N100)? mem[67] : 
                     (N102)? mem[74] : 
                     (N104)? mem[81] : 
                     (N106)? mem[88] : 
                     (N108)? mem[95] : 
                     (N110)? mem[102] : 
                     (N112)? mem[109] : 
                     (N114)? mem[116] : 
                     (N116)? mem[123] : 
                     (N118)? mem[130] : 
                     (N120)? mem[137] : 
                     (N122)? mem[144] : 
                     (N124)? mem[151] : 
                     (N126)? mem[158] : 
                     (N128)? mem[165] : 
                     (N130)? mem[172] : 
                     (N132)? mem[179] : 
                     (N134)? mem[186] : 
                     (N136)? mem[193] : 
                     (N138)? mem[200] : 
                     (N140)? mem[207] : 
                     (N142)? mem[214] : 
                     (N144)? mem[221] : 
                     (N83)? mem[228] : 
                     (N85)? mem[235] : 
                     (N87)? mem[242] : 
                     (N89)? mem[249] : 
                     (N91)? mem[256] : 
                     (N93)? mem[263] : 
                     (N95)? mem[270] : 
                     (N97)? mem[277] : 
                     (N99)? mem[284] : 
                     (N101)? mem[291] : 
                     (N103)? mem[298] : 
                     (N105)? mem[305] : 
                     (N107)? mem[312] : 
                     (N109)? mem[319] : 
                     (N111)? mem[326] : 
                     (N113)? mem[333] : 
                     (N115)? mem[340] : 
                     (N117)? mem[347] : 
                     (N119)? mem[354] : 
                     (N121)? mem[361] : 
                     (N123)? mem[368] : 
                     (N125)? mem[375] : 
                     (N127)? mem[382] : 
                     (N129)? mem[389] : 
                     (N131)? mem[396] : 
                     (N133)? mem[403] : 
                     (N135)? mem[410] : 
                     (N137)? mem[417] : 
                     (N139)? mem[424] : 
                     (N141)? mem[431] : 
                     (N143)? mem[438] : 
                     (N145)? mem[445] : 1'b0;
  assign data_o[3] = (N82)? mem[3] : 
                     (N84)? mem[10] : 
                     (N86)? mem[17] : 
                     (N88)? mem[24] : 
                     (N90)? mem[31] : 
                     (N92)? mem[38] : 
                     (N94)? mem[45] : 
                     (N96)? mem[52] : 
                     (N98)? mem[59] : 
                     (N100)? mem[66] : 
                     (N102)? mem[73] : 
                     (N104)? mem[80] : 
                     (N106)? mem[87] : 
                     (N108)? mem[94] : 
                     (N110)? mem[101] : 
                     (N112)? mem[108] : 
                     (N114)? mem[115] : 
                     (N116)? mem[122] : 
                     (N118)? mem[129] : 
                     (N120)? mem[136] : 
                     (N122)? mem[143] : 
                     (N124)? mem[150] : 
                     (N126)? mem[157] : 
                     (N128)? mem[164] : 
                     (N130)? mem[171] : 
                     (N132)? mem[178] : 
                     (N134)? mem[185] : 
                     (N136)? mem[192] : 
                     (N138)? mem[199] : 
                     (N140)? mem[206] : 
                     (N142)? mem[213] : 
                     (N144)? mem[220] : 
                     (N83)? mem[227] : 
                     (N85)? mem[234] : 
                     (N87)? mem[241] : 
                     (N89)? mem[248] : 
                     (N91)? mem[255] : 
                     (N93)? mem[262] : 
                     (N95)? mem[269] : 
                     (N97)? mem[276] : 
                     (N99)? mem[283] : 
                     (N101)? mem[290] : 
                     (N103)? mem[297] : 
                     (N105)? mem[304] : 
                     (N107)? mem[311] : 
                     (N109)? mem[318] : 
                     (N111)? mem[325] : 
                     (N113)? mem[332] : 
                     (N115)? mem[339] : 
                     (N117)? mem[346] : 
                     (N119)? mem[353] : 
                     (N121)? mem[360] : 
                     (N123)? mem[367] : 
                     (N125)? mem[374] : 
                     (N127)? mem[381] : 
                     (N129)? mem[388] : 
                     (N131)? mem[395] : 
                     (N133)? mem[402] : 
                     (N135)? mem[409] : 
                     (N137)? mem[416] : 
                     (N139)? mem[423] : 
                     (N141)? mem[430] : 
                     (N143)? mem[437] : 
                     (N145)? mem[444] : 1'b0;
  assign data_o[2] = (N82)? mem[2] : 
                     (N84)? mem[9] : 
                     (N86)? mem[16] : 
                     (N88)? mem[23] : 
                     (N90)? mem[30] : 
                     (N92)? mem[37] : 
                     (N94)? mem[44] : 
                     (N96)? mem[51] : 
                     (N98)? mem[58] : 
                     (N100)? mem[65] : 
                     (N102)? mem[72] : 
                     (N104)? mem[79] : 
                     (N106)? mem[86] : 
                     (N108)? mem[93] : 
                     (N110)? mem[100] : 
                     (N112)? mem[107] : 
                     (N114)? mem[114] : 
                     (N116)? mem[121] : 
                     (N118)? mem[128] : 
                     (N120)? mem[135] : 
                     (N122)? mem[142] : 
                     (N124)? mem[149] : 
                     (N126)? mem[156] : 
                     (N128)? mem[163] : 
                     (N130)? mem[170] : 
                     (N132)? mem[177] : 
                     (N134)? mem[184] : 
                     (N136)? mem[191] : 
                     (N138)? mem[198] : 
                     (N140)? mem[205] : 
                     (N142)? mem[212] : 
                     (N144)? mem[219] : 
                     (N83)? mem[226] : 
                     (N85)? mem[233] : 
                     (N87)? mem[240] : 
                     (N89)? mem[247] : 
                     (N91)? mem[254] : 
                     (N93)? mem[261] : 
                     (N95)? mem[268] : 
                     (N97)? mem[275] : 
                     (N99)? mem[282] : 
                     (N101)? mem[289] : 
                     (N103)? mem[296] : 
                     (N105)? mem[303] : 
                     (N107)? mem[310] : 
                     (N109)? mem[317] : 
                     (N111)? mem[324] : 
                     (N113)? mem[331] : 
                     (N115)? mem[338] : 
                     (N117)? mem[345] : 
                     (N119)? mem[352] : 
                     (N121)? mem[359] : 
                     (N123)? mem[366] : 
                     (N125)? mem[373] : 
                     (N127)? mem[380] : 
                     (N129)? mem[387] : 
                     (N131)? mem[394] : 
                     (N133)? mem[401] : 
                     (N135)? mem[408] : 
                     (N137)? mem[415] : 
                     (N139)? mem[422] : 
                     (N141)? mem[429] : 
                     (N143)? mem[436] : 
                     (N145)? mem[443] : 1'b0;
  assign data_o[1] = (N82)? mem[1] : 
                     (N84)? mem[8] : 
                     (N86)? mem[15] : 
                     (N88)? mem[22] : 
                     (N90)? mem[29] : 
                     (N92)? mem[36] : 
                     (N94)? mem[43] : 
                     (N96)? mem[50] : 
                     (N98)? mem[57] : 
                     (N100)? mem[64] : 
                     (N102)? mem[71] : 
                     (N104)? mem[78] : 
                     (N106)? mem[85] : 
                     (N108)? mem[92] : 
                     (N110)? mem[99] : 
                     (N112)? mem[106] : 
                     (N114)? mem[113] : 
                     (N116)? mem[120] : 
                     (N118)? mem[127] : 
                     (N120)? mem[134] : 
                     (N122)? mem[141] : 
                     (N124)? mem[148] : 
                     (N126)? mem[155] : 
                     (N128)? mem[162] : 
                     (N130)? mem[169] : 
                     (N132)? mem[176] : 
                     (N134)? mem[183] : 
                     (N136)? mem[190] : 
                     (N138)? mem[197] : 
                     (N140)? mem[204] : 
                     (N142)? mem[211] : 
                     (N144)? mem[218] : 
                     (N83)? mem[225] : 
                     (N85)? mem[232] : 
                     (N87)? mem[239] : 
                     (N89)? mem[246] : 
                     (N91)? mem[253] : 
                     (N93)? mem[260] : 
                     (N95)? mem[267] : 
                     (N97)? mem[274] : 
                     (N99)? mem[281] : 
                     (N101)? mem[288] : 
                     (N103)? mem[295] : 
                     (N105)? mem[302] : 
                     (N107)? mem[309] : 
                     (N109)? mem[316] : 
                     (N111)? mem[323] : 
                     (N113)? mem[330] : 
                     (N115)? mem[337] : 
                     (N117)? mem[344] : 
                     (N119)? mem[351] : 
                     (N121)? mem[358] : 
                     (N123)? mem[365] : 
                     (N125)? mem[372] : 
                     (N127)? mem[379] : 
                     (N129)? mem[386] : 
                     (N131)? mem[393] : 
                     (N133)? mem[400] : 
                     (N135)? mem[407] : 
                     (N137)? mem[414] : 
                     (N139)? mem[421] : 
                     (N141)? mem[428] : 
                     (N143)? mem[435] : 
                     (N145)? mem[442] : 1'b0;
  assign data_o[0] = (N82)? mem[0] : 
                     (N84)? mem[7] : 
                     (N86)? mem[14] : 
                     (N88)? mem[21] : 
                     (N90)? mem[28] : 
                     (N92)? mem[35] : 
                     (N94)? mem[42] : 
                     (N96)? mem[49] : 
                     (N98)? mem[56] : 
                     (N100)? mem[63] : 
                     (N102)? mem[70] : 
                     (N104)? mem[77] : 
                     (N106)? mem[84] : 
                     (N108)? mem[91] : 
                     (N110)? mem[98] : 
                     (N112)? mem[105] : 
                     (N114)? mem[112] : 
                     (N116)? mem[119] : 
                     (N118)? mem[126] : 
                     (N120)? mem[133] : 
                     (N122)? mem[140] : 
                     (N124)? mem[147] : 
                     (N126)? mem[154] : 
                     (N128)? mem[161] : 
                     (N130)? mem[168] : 
                     (N132)? mem[175] : 
                     (N134)? mem[182] : 
                     (N136)? mem[189] : 
                     (N138)? mem[196] : 
                     (N140)? mem[203] : 
                     (N142)? mem[210] : 
                     (N144)? mem[217] : 
                     (N83)? mem[224] : 
                     (N85)? mem[231] : 
                     (N87)? mem[238] : 
                     (N89)? mem[245] : 
                     (N91)? mem[252] : 
                     (N93)? mem[259] : 
                     (N95)? mem[266] : 
                     (N97)? mem[273] : 
                     (N99)? mem[280] : 
                     (N101)? mem[287] : 
                     (N103)? mem[294] : 
                     (N105)? mem[301] : 
                     (N107)? mem[308] : 
                     (N109)? mem[315] : 
                     (N111)? mem[322] : 
                     (N113)? mem[329] : 
                     (N115)? mem[336] : 
                     (N117)? mem[343] : 
                     (N119)? mem[350] : 
                     (N121)? mem[357] : 
                     (N123)? mem[364] : 
                     (N125)? mem[371] : 
                     (N127)? mem[378] : 
                     (N129)? mem[385] : 
                     (N131)? mem[392] : 
                     (N133)? mem[399] : 
                     (N135)? mem[406] : 
                     (N137)? mem[413] : 
                     (N139)? mem[420] : 
                     (N141)? mem[427] : 
                     (N143)? mem[434] : 
                     (N145)? mem[441] : 1'b0;

  always @(posedge clk_i) begin
    if(N1114) begin
      mem_447_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1113) begin
      mem_446_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1112) begin
      mem_445_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1111) begin
      mem_444_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1110) begin
      mem_443_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1109) begin
      mem_442_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1108) begin
      mem_441_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1107) begin
      mem_440_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1106) begin
      mem_439_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1105) begin
      mem_438_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1104) begin
      mem_437_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1103) begin
      mem_436_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1102) begin
      mem_435_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1101) begin
      mem_434_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1100) begin
      mem_433_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1099) begin
      mem_432_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1098) begin
      mem_431_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1097) begin
      mem_430_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1096) begin
      mem_429_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1095) begin
      mem_428_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1094) begin
      mem_427_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1093) begin
      mem_426_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1092) begin
      mem_425_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1091) begin
      mem_424_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1090) begin
      mem_423_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1089) begin
      mem_422_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1088) begin
      mem_421_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1087) begin
      mem_420_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1086) begin
      mem_419_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1085) begin
      mem_418_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1084) begin
      mem_417_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1083) begin
      mem_416_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1082) begin
      mem_415_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1081) begin
      mem_414_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1080) begin
      mem_413_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1079) begin
      mem_412_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1078) begin
      mem_411_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1077) begin
      mem_410_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1076) begin
      mem_409_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1075) begin
      mem_408_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1074) begin
      mem_407_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1073) begin
      mem_406_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1072) begin
      mem_405_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1071) begin
      mem_404_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1070) begin
      mem_403_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1069) begin
      mem_402_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1068) begin
      mem_401_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1067) begin
      mem_400_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1066) begin
      mem_399_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1065) begin
      mem_398_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1064) begin
      mem_397_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1063) begin
      mem_396_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1062) begin
      mem_395_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1061) begin
      mem_394_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1060) begin
      mem_393_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1059) begin
      mem_392_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1058) begin
      mem_391_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1057) begin
      mem_390_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1056) begin
      mem_389_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1055) begin
      mem_388_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1054) begin
      mem_387_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1053) begin
      mem_386_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1052) begin
      mem_385_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1051) begin
      mem_384_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1050) begin
      mem_383_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1049) begin
      mem_382_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1048) begin
      mem_381_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1047) begin
      mem_380_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1046) begin
      mem_379_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1045) begin
      mem_378_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1044) begin
      mem_377_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1043) begin
      mem_376_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1042) begin
      mem_375_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1041) begin
      mem_374_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1040) begin
      mem_373_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1039) begin
      mem_372_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1038) begin
      mem_371_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1037) begin
      mem_370_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1036) begin
      mem_369_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1035) begin
      mem_368_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1034) begin
      mem_367_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1033) begin
      mem_366_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1032) begin
      mem_365_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1031) begin
      mem_364_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1030) begin
      mem_363_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1029) begin
      mem_362_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1028) begin
      mem_361_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1027) begin
      mem_360_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1026) begin
      mem_359_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1025) begin
      mem_358_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1024) begin
      mem_357_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1023) begin
      mem_356_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1022) begin
      mem_355_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1021) begin
      mem_354_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1020) begin
      mem_353_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1019) begin
      mem_352_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1018) begin
      mem_351_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1017) begin
      mem_350_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1016) begin
      mem_349_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1015) begin
      mem_348_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1014) begin
      mem_347_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1013) begin
      mem_346_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1012) begin
      mem_345_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1011) begin
      mem_344_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1010) begin
      mem_343_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1009) begin
      mem_342_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1008) begin
      mem_341_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1007) begin
      mem_340_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N1006) begin
      mem_339_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N1005) begin
      mem_338_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N1004) begin
      mem_337_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N1003) begin
      mem_336_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N1002) begin
      mem_335_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N1001) begin
      mem_334_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N1000) begin
      mem_333_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N999) begin
      mem_332_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N998) begin
      mem_331_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N997) begin
      mem_330_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N996) begin
      mem_329_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N995) begin
      mem_328_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N994) begin
      mem_327_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N993) begin
      mem_326_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N992) begin
      mem_325_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N991) begin
      mem_324_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N990) begin
      mem_323_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N989) begin
      mem_322_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N988) begin
      mem_321_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N987) begin
      mem_320_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N986) begin
      mem_319_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N985) begin
      mem_318_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N984) begin
      mem_317_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N983) begin
      mem_316_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N982) begin
      mem_315_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N981) begin
      mem_314_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N980) begin
      mem_313_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N979) begin
      mem_312_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N978) begin
      mem_311_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N977) begin
      mem_310_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N976) begin
      mem_309_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N975) begin
      mem_308_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N974) begin
      mem_307_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N973) begin
      mem_306_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N972) begin
      mem_305_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N971) begin
      mem_304_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N970) begin
      mem_303_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N969) begin
      mem_302_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N968) begin
      mem_301_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N967) begin
      mem_300_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N966) begin
      mem_299_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N965) begin
      mem_298_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N964) begin
      mem_297_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N963) begin
      mem_296_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N962) begin
      mem_295_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N961) begin
      mem_294_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N960) begin
      mem_293_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N959) begin
      mem_292_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N958) begin
      mem_291_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N957) begin
      mem_290_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N956) begin
      mem_289_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N955) begin
      mem_288_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N954) begin
      mem_287_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N953) begin
      mem_286_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N952) begin
      mem_285_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N951) begin
      mem_284_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N950) begin
      mem_283_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N949) begin
      mem_282_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N948) begin
      mem_281_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N947) begin
      mem_280_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N946) begin
      mem_279_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N945) begin
      mem_278_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N944) begin
      mem_277_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N943) begin
      mem_276_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N942) begin
      mem_275_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N941) begin
      mem_274_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N940) begin
      mem_273_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N939) begin
      mem_272_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N938) begin
      mem_271_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N937) begin
      mem_270_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N936) begin
      mem_269_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N935) begin
      mem_268_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N934) begin
      mem_267_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N933) begin
      mem_266_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N932) begin
      mem_265_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N931) begin
      mem_264_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N930) begin
      mem_263_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N929) begin
      mem_262_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N928) begin
      mem_261_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N927) begin
      mem_260_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N926) begin
      mem_259_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N925) begin
      mem_258_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N924) begin
      mem_257_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N923) begin
      mem_256_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N922) begin
      mem_255_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N921) begin
      mem_254_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N920) begin
      mem_253_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N919) begin
      mem_252_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N918) begin
      mem_251_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N917) begin
      mem_250_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N916) begin
      mem_249_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N915) begin
      mem_248_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N914) begin
      mem_247_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N913) begin
      mem_246_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N912) begin
      mem_245_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N911) begin
      mem_244_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N910) begin
      mem_243_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N909) begin
      mem_242_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N908) begin
      mem_241_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N907) begin
      mem_240_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N906) begin
      mem_239_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N905) begin
      mem_238_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N904) begin
      mem_237_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N903) begin
      mem_236_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N902) begin
      mem_235_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N901) begin
      mem_234_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N900) begin
      mem_233_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N899) begin
      mem_232_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N898) begin
      mem_231_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N897) begin
      mem_230_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N896) begin
      mem_229_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N895) begin
      mem_228_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N894) begin
      mem_227_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N893) begin
      mem_226_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N892) begin
      mem_225_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N891) begin
      mem_224_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N890) begin
      mem_223_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N889) begin
      mem_222_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N888) begin
      mem_221_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N887) begin
      mem_220_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N886) begin
      mem_219_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N885) begin
      mem_218_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N884) begin
      mem_217_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N883) begin
      mem_216_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N882) begin
      mem_215_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N881) begin
      mem_214_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N880) begin
      mem_213_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N879) begin
      mem_212_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N878) begin
      mem_211_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N877) begin
      mem_210_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N876) begin
      mem_209_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N875) begin
      mem_208_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N874) begin
      mem_207_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N873) begin
      mem_206_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N872) begin
      mem_205_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N871) begin
      mem_204_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N870) begin
      mem_203_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N869) begin
      mem_202_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N868) begin
      mem_201_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N867) begin
      mem_200_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N866) begin
      mem_199_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N865) begin
      mem_198_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N864) begin
      mem_197_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N863) begin
      mem_196_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N862) begin
      mem_195_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N861) begin
      mem_194_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N860) begin
      mem_193_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N859) begin
      mem_192_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N858) begin
      mem_191_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N857) begin
      mem_190_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N856) begin
      mem_189_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N855) begin
      mem_188_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N854) begin
      mem_187_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N853) begin
      mem_186_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N852) begin
      mem_185_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N851) begin
      mem_184_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N850) begin
      mem_183_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N849) begin
      mem_182_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N848) begin
      mem_181_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N847) begin
      mem_180_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N846) begin
      mem_179_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N845) begin
      mem_178_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N844) begin
      mem_177_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N843) begin
      mem_176_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N842) begin
      mem_175_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N841) begin
      mem_174_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N840) begin
      mem_173_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N839) begin
      mem_172_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N838) begin
      mem_171_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N837) begin
      mem_170_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N836) begin
      mem_169_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N835) begin
      mem_168_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N834) begin
      mem_167_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N833) begin
      mem_166_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N832) begin
      mem_165_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N831) begin
      mem_164_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N830) begin
      mem_163_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N829) begin
      mem_162_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N828) begin
      mem_161_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N827) begin
      mem_160_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N826) begin
      mem_159_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N825) begin
      mem_158_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N824) begin
      mem_157_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N823) begin
      mem_156_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N822) begin
      mem_155_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N821) begin
      mem_154_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N820) begin
      mem_153_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N819) begin
      mem_152_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N818) begin
      mem_151_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N817) begin
      mem_150_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N816) begin
      mem_149_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N815) begin
      mem_148_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N814) begin
      mem_147_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N813) begin
      mem_146_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N812) begin
      mem_145_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N811) begin
      mem_144_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N810) begin
      mem_143_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N809) begin
      mem_142_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N808) begin
      mem_141_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N807) begin
      mem_140_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N806) begin
      mem_139_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N805) begin
      mem_138_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N804) begin
      mem_137_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N803) begin
      mem_136_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N802) begin
      mem_135_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N801) begin
      mem_134_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N800) begin
      mem_133_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N799) begin
      mem_132_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N798) begin
      mem_131_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N797) begin
      mem_130_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N796) begin
      mem_129_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N795) begin
      mem_128_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N794) begin
      mem_127_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N793) begin
      mem_126_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N792) begin
      mem_125_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N791) begin
      mem_124_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N790) begin
      mem_123_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N789) begin
      mem_122_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N788) begin
      mem_121_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N787) begin
      mem_120_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N786) begin
      mem_119_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N785) begin
      mem_118_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N784) begin
      mem_117_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N783) begin
      mem_116_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N782) begin
      mem_115_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N781) begin
      mem_114_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N780) begin
      mem_113_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N779) begin
      mem_112_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N778) begin
      mem_111_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N777) begin
      mem_110_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N776) begin
      mem_109_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N775) begin
      mem_108_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N774) begin
      mem_107_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N773) begin
      mem_106_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N772) begin
      mem_105_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N771) begin
      mem_104_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N770) begin
      mem_103_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N769) begin
      mem_102_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N768) begin
      mem_101_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N767) begin
      mem_100_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N766) begin
      mem_99_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N765) begin
      mem_98_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N764) begin
      mem_97_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N763) begin
      mem_96_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N762) begin
      mem_95_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N761) begin
      mem_94_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N760) begin
      mem_93_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N759) begin
      mem_92_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N758) begin
      mem_91_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N757) begin
      mem_90_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N756) begin
      mem_89_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N755) begin
      mem_88_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N754) begin
      mem_87_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N753) begin
      mem_86_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N752) begin
      mem_85_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N751) begin
      mem_84_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N750) begin
      mem_83_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N749) begin
      mem_82_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N748) begin
      mem_81_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N747) begin
      mem_80_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N746) begin
      mem_79_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N745) begin
      mem_78_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N744) begin
      mem_77_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N743) begin
      mem_76_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N742) begin
      mem_75_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N741) begin
      mem_74_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N740) begin
      mem_73_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N739) begin
      mem_72_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N738) begin
      mem_71_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N737) begin
      mem_70_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N736) begin
      mem_69_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N735) begin
      mem_68_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N734) begin
      mem_67_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N733) begin
      mem_66_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N732) begin
      mem_65_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N731) begin
      mem_64_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N730) begin
      mem_63_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N729) begin
      mem_62_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N728) begin
      mem_61_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N727) begin
      mem_60_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N726) begin
      mem_59_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N725) begin
      mem_58_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N724) begin
      mem_57_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N723) begin
      mem_56_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N722) begin
      mem_55_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N721) begin
      mem_54_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N720) begin
      mem_53_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N719) begin
      mem_52_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N718) begin
      mem_51_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N717) begin
      mem_50_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N716) begin
      mem_49_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N715) begin
      mem_48_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N714) begin
      mem_47_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N713) begin
      mem_46_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N712) begin
      mem_45_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N711) begin
      mem_44_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N710) begin
      mem_43_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N709) begin
      mem_42_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N708) begin
      mem_41_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N707) begin
      mem_40_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N706) begin
      mem_39_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N705) begin
      mem_38_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N704) begin
      mem_37_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N703) begin
      mem_36_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N702) begin
      mem_35_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N701) begin
      mem_34_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N700) begin
      mem_33_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N699) begin
      mem_32_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N698) begin
      mem_31_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N697) begin
      mem_30_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N696) begin
      mem_29_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N695) begin
      mem_28_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N694) begin
      mem_27_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N693) begin
      mem_26_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N692) begin
      mem_25_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N691) begin
      mem_24_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N690) begin
      mem_23_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N689) begin
      mem_22_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N688) begin
      mem_21_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N687) begin
      mem_20_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N686) begin
      mem_19_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N685) begin
      mem_18_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N684) begin
      mem_17_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N683) begin
      mem_16_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N682) begin
      mem_15_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N681) begin
      mem_14_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N680) begin
      mem_13_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N679) begin
      mem_12_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N678) begin
      mem_11_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N677) begin
      mem_10_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N676) begin
      mem_9_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N675) begin
      mem_8_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N674) begin
      mem_7_sv2v_reg <= data_i[0];
    end 
  end


  always @(posedge clk_i) begin
    if(N673) begin
      mem_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(N672) begin
      mem_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(N671) begin
      mem_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(N670) begin
      mem_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(N669) begin
      mem_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(N668) begin
      mem_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(N667) begin
      mem_0_sv2v_reg <= data_i[0];
    end 
  end

  assign N1115 = ~addr_i[5];
  assign N1116 = addr_i[3] & addr_i[4];
  assign N1117 = N0 & addr_i[4];
  assign N0 = ~addr_i[3];
  assign N1118 = addr_i[3] & N1;
  assign N1 = ~addr_i[4];
  assign N1119 = N2 & N3;
  assign N2 = ~addr_i[3];
  assign N3 = ~addr_i[4];
  assign N1120 = addr_i[5] & N1116;
  assign N1121 = addr_i[5] & N1117;
  assign N1122 = addr_i[5] & N1118;
  assign N1123 = addr_i[5] & N1119;
  assign N1124 = N1115 & N1116;
  assign N1125 = N1115 & N1117;
  assign N1126 = N1115 & N1118;
  assign N1127 = N1115 & N1119;
  assign N1128 = ~addr_i[2];
  assign N1129 = addr_i[0] & addr_i[1];
  assign N1130 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N1131 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N1132 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N1133 = addr_i[2] & N1129;
  assign N1134 = addr_i[2] & N1130;
  assign N1135 = addr_i[2] & N1131;
  assign N1136 = addr_i[2] & N1132;
  assign N1137 = N1128 & N1129;
  assign N1138 = N1128 & N1130;
  assign N1139 = N1128 & N1131;
  assign N1140 = N1128 & N1132;
  assign N602 = N1120 & N1133;
  assign N601 = N1120 & N1134;
  assign N600 = N1120 & N1135;
  assign N599 = N1120 & N1136;
  assign N598 = N1120 & N1137;
  assign N597 = N1120 & N1138;
  assign N596 = N1120 & N1139;
  assign N595 = N1120 & N1140;
  assign N594 = N1121 & N1133;
  assign N593 = N1121 & N1134;
  assign N592 = N1121 & N1135;
  assign N591 = N1121 & N1136;
  assign N590 = N1121 & N1137;
  assign N589 = N1121 & N1138;
  assign N588 = N1121 & N1139;
  assign N587 = N1121 & N1140;
  assign N586 = N1122 & N1133;
  assign N585 = N1122 & N1134;
  assign N584 = N1122 & N1135;
  assign N583 = N1122 & N1136;
  assign N582 = N1122 & N1137;
  assign N581 = N1122 & N1138;
  assign N580 = N1122 & N1139;
  assign N579 = N1122 & N1140;
  assign N578 = N1123 & N1133;
  assign N577 = N1123 & N1134;
  assign N576 = N1123 & N1135;
  assign N575 = N1123 & N1136;
  assign N574 = N1123 & N1137;
  assign N573 = N1123 & N1138;
  assign N572 = N1123 & N1139;
  assign N571 = N1123 & N1140;
  assign N570 = N1124 & N1133;
  assign N569 = N1124 & N1134;
  assign N568 = N1124 & N1135;
  assign N567 = N1124 & N1136;
  assign N566 = N1124 & N1137;
  assign N565 = N1124 & N1138;
  assign N564 = N1124 & N1139;
  assign N563 = N1124 & N1140;
  assign N562 = N1125 & N1133;
  assign N561 = N1125 & N1134;
  assign N560 = N1125 & N1135;
  assign N559 = N1125 & N1136;
  assign N558 = N1125 & N1137;
  assign N557 = N1125 & N1138;
  assign N556 = N1125 & N1139;
  assign N555 = N1125 & N1140;
  assign N554 = N1126 & N1133;
  assign N553 = N1126 & N1134;
  assign N552 = N1126 & N1135;
  assign N551 = N1126 & N1136;
  assign N550 = N1126 & N1137;
  assign N549 = N1126 & N1138;
  assign N548 = N1126 & N1139;
  assign N547 = N1126 & N1140;
  assign N546 = N1127 & N1133;
  assign N545 = N1127 & N1134;
  assign N544 = N1127 & N1135;
  assign N543 = N1127 & N1136;
  assign N542 = N1127 & N1137;
  assign N541 = N1127 & N1138;
  assign N540 = N1127 & N1139;
  assign N539 = N1127 & N1140;
  assign { N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149 } = (N8)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_mask_i[0];
  assign { N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214 } = (N9)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N213)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = w_mask_i[1];
  assign { N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279 } = (N10)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N278)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = w_mask_i[2];
  assign { N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344 } = (N11)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N343)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N11 = w_mask_i[3];
  assign { N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409 } = (N12)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N408)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = w_mask_i[4];
  assign { N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474 } = (N13)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N473)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = w_mask_i[5];
  assign { N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603 } = (N14)? { N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N538)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = w_mask_i[6];
  assign { N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667 } = (N15)? { N666, N537, N472, N407, N342, N277, N212, N665, N536, N471, N406, N341, N276, N211, N664, N535, N470, N405, N340, N275, N210, N663, N534, N469, N404, N339, N274, N209, N662, N533, N468, N403, N338, N273, N208, N661, N532, N467, N402, N337, N272, N207, N660, N531, N466, N401, N336, N271, N206, N659, N530, N465, N400, N335, N270, N205, N658, N529, N464, N399, N334, N269, N204, N657, N528, N463, N398, N333, N268, N203, N656, N527, N462, N397, N332, N267, N202, N655, N526, N461, N396, N331, N266, N201, N654, N525, N460, N395, N330, N265, N200, N653, N524, N459, N394, N329, N264, N199, N652, N523, N458, N393, N328, N263, N198, N651, N522, N457, N392, N327, N262, N197, N650, N521, N456, N391, N326, N261, N196, N649, N520, N455, N390, N325, N260, N195, N648, N519, N454, N389, N324, N259, N194, N647, N518, N453, N388, N323, N258, N193, N646, N517, N452, N387, N322, N257, N192, N645, N516, N451, N386, N321, N256, N191, N644, N515, N450, N385, N320, N255, N190, N643, N514, N449, N384, N319, N254, N189, N642, N513, N448, N383, N318, N253, N188, N641, N512, N447, N382, N317, N252, N187, N640, N511, N446, N381, N316, N251, N186, N639, N510, N445, N380, N315, N250, N185, N638, N509, N444, N379, N314, N249, N184, N637, N508, N443, N378, N313, N248, N183, N636, N507, N442, N377, N312, N247, N182, N635, N506, N441, N376, N311, N246, N181, N634, N505, N440, N375, N310, N245, N180, N633, N504, N439, N374, N309, N244, N179, N632, N503, N438, N373, N308, N243, N178, N631, N502, N437, N372, N307, N242, N177, N630, N501, N436, N371, N306, N241, N176, N629, N500, N435, N370, N305, N240, N175, N628, N499, N434, N369, N304, N239, N174, N627, N498, N433, N368, N303, N238, N173, N626, N497, N432, N367, N302, N237, N172, N625, N496, N431, N366, N301, N236, N171, N624, N495, N430, N365, N300, N235, N170, N623, N494, N429, N364, N299, N234, N169, N622, N493, N428, N363, N298, N233, N168, N621, N492, N427, N362, N297, N232, N167, N620, N491, N426, N361, N296, N231, N166, N619, N490, N425, N360, N295, N230, N165, N618, N489, N424, N359, N294, N229, N164, N617, N488, N423, N358, N293, N228, N163, N616, N487, N422, N357, N292, N227, N162, N615, N486, N421, N356, N291, N226, N161, N614, N485, N420, N355, N290, N225, N160, N613, N484, N419, N354, N289, N224, N159, N612, N483, N418, N353, N288, N223, N158, N611, N482, N417, N352, N287, N222, N157, N610, N481, N416, N351, N286, N221, N156, N609, N480, N415, N350, N285, N220, N155, N608, N479, N414, N349, N284, N219, N154, N607, N478, N413, N348, N283, N218, N153, N606, N477, N412, N347, N282, N217, N152, N605, N476, N411, N346, N281, N216, N151, N604, N475, N410, N345, N280, N215, N150, N603, N474, N409, N344, N279, N214, N149 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (N147)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N15 = N146;
  assign N16 = ~addr_r[0];
  assign N17 = ~addr_r[1];
  assign N18 = N16 & N17;
  assign N19 = N16 & addr_r[1];
  assign N20 = addr_r[0] & N17;
  assign N21 = addr_r[0] & addr_r[1];
  assign N22 = ~addr_r[2];
  assign N23 = N18 & N22;
  assign N24 = N18 & addr_r[2];
  assign N25 = N20 & N22;
  assign N26 = N20 & addr_r[2];
  assign N27 = N19 & N22;
  assign N28 = N19 & addr_r[2];
  assign N29 = N21 & N22;
  assign N30 = N21 & addr_r[2];
  assign N31 = ~addr_r[3];
  assign N32 = N23 & N31;
  assign N33 = N23 & addr_r[3];
  assign N34 = N25 & N31;
  assign N35 = N25 & addr_r[3];
  assign N36 = N27 & N31;
  assign N37 = N27 & addr_r[3];
  assign N38 = N29 & N31;
  assign N39 = N29 & addr_r[3];
  assign N40 = N24 & N31;
  assign N41 = N24 & addr_r[3];
  assign N42 = N26 & N31;
  assign N43 = N26 & addr_r[3];
  assign N44 = N28 & N31;
  assign N45 = N28 & addr_r[3];
  assign N46 = N30 & N31;
  assign N47 = N30 & addr_r[3];
  assign N48 = ~addr_r[4];
  assign N49 = N32 & N48;
  assign N50 = N32 & addr_r[4];
  assign N51 = N34 & N48;
  assign N52 = N34 & addr_r[4];
  assign N53 = N36 & N48;
  assign N54 = N36 & addr_r[4];
  assign N55 = N38 & N48;
  assign N56 = N38 & addr_r[4];
  assign N57 = N40 & N48;
  assign N58 = N40 & addr_r[4];
  assign N59 = N42 & N48;
  assign N60 = N42 & addr_r[4];
  assign N61 = N44 & N48;
  assign N62 = N44 & addr_r[4];
  assign N63 = N46 & N48;
  assign N64 = N46 & addr_r[4];
  assign N65 = N33 & N48;
  assign N66 = N33 & addr_r[4];
  assign N67 = N35 & N48;
  assign N68 = N35 & addr_r[4];
  assign N69 = N37 & N48;
  assign N70 = N37 & addr_r[4];
  assign N71 = N39 & N48;
  assign N72 = N39 & addr_r[4];
  assign N73 = N41 & N48;
  assign N74 = N41 & addr_r[4];
  assign N75 = N43 & N48;
  assign N76 = N43 & addr_r[4];
  assign N77 = N45 & N48;
  assign N78 = N45 & addr_r[4];
  assign N79 = N47 & N48;
  assign N80 = N47 & addr_r[4];
  assign N81 = ~addr_r[5];
  assign N82 = N49 & N81;
  assign N83 = N49 & addr_r[5];
  assign N84 = N51 & N81;
  assign N85 = N51 & addr_r[5];
  assign N86 = N53 & N81;
  assign N87 = N53 & addr_r[5];
  assign N88 = N55 & N81;
  assign N89 = N55 & addr_r[5];
  assign N90 = N57 & N81;
  assign N91 = N57 & addr_r[5];
  assign N92 = N59 & N81;
  assign N93 = N59 & addr_r[5];
  assign N94 = N61 & N81;
  assign N95 = N61 & addr_r[5];
  assign N96 = N63 & N81;
  assign N97 = N63 & addr_r[5];
  assign N98 = N65 & N81;
  assign N99 = N65 & addr_r[5];
  assign N100 = N67 & N81;
  assign N101 = N67 & addr_r[5];
  assign N102 = N69 & N81;
  assign N103 = N69 & addr_r[5];
  assign N104 = N71 & N81;
  assign N105 = N71 & addr_r[5];
  assign N106 = N73 & N81;
  assign N107 = N73 & addr_r[5];
  assign N108 = N75 & N81;
  assign N109 = N75 & addr_r[5];
  assign N110 = N77 & N81;
  assign N111 = N77 & addr_r[5];
  assign N112 = N79 & N81;
  assign N113 = N79 & addr_r[5];
  assign N114 = N50 & N81;
  assign N115 = N50 & addr_r[5];
  assign N116 = N52 & N81;
  assign N117 = N52 & addr_r[5];
  assign N118 = N54 & N81;
  assign N119 = N54 & addr_r[5];
  assign N120 = N56 & N81;
  assign N121 = N56 & addr_r[5];
  assign N122 = N58 & N81;
  assign N123 = N58 & addr_r[5];
  assign N124 = N60 & N81;
  assign N125 = N60 & addr_r[5];
  assign N126 = N62 & N81;
  assign N127 = N62 & addr_r[5];
  assign N128 = N64 & N81;
  assign N129 = N64 & addr_r[5];
  assign N130 = N66 & N81;
  assign N131 = N66 & addr_r[5];
  assign N132 = N68 & N81;
  assign N133 = N68 & addr_r[5];
  assign N134 = N70 & N81;
  assign N135 = N70 & addr_r[5];
  assign N136 = N72 & N81;
  assign N137 = N72 & addr_r[5];
  assign N138 = N74 & N81;
  assign N139 = N74 & addr_r[5];
  assign N140 = N76 & N81;
  assign N141 = N76 & addr_r[5];
  assign N142 = N78 & N81;
  assign N143 = N78 & addr_r[5];
  assign N144 = N80 & N81;
  assign N145 = N80 & addr_r[5];
  assign N146 = v_i & w_i;
  assign N147 = ~N146;
  assign N148 = ~w_mask_i[0];
  assign N213 = ~w_mask_i[1];
  assign N278 = ~w_mask_i[2];
  assign N343 = ~w_mask_i[3];
  assign N408 = ~w_mask_i[4];
  assign N473 = ~w_mask_i[5];
  assign N538 = ~w_mask_i[6];

endmodule