module bsg_dff_width_p295
(
  clk_i,
  data_i,
  data_o
);

  input [294:0] data_i;
  output [294:0] data_o;
  input clk_i;
  wire [294:0] data_o;
  reg data_o_294_sv2v_reg,data_o_293_sv2v_reg,data_o_292_sv2v_reg,data_o_291_sv2v_reg,
  data_o_290_sv2v_reg,data_o_289_sv2v_reg,data_o_288_sv2v_reg,data_o_287_sv2v_reg,
  data_o_286_sv2v_reg,data_o_285_sv2v_reg,data_o_284_sv2v_reg,data_o_283_sv2v_reg,
  data_o_282_sv2v_reg,data_o_281_sv2v_reg,data_o_280_sv2v_reg,data_o_279_sv2v_reg,
  data_o_278_sv2v_reg,data_o_277_sv2v_reg,data_o_276_sv2v_reg,data_o_275_sv2v_reg,
  data_o_274_sv2v_reg,data_o_273_sv2v_reg,data_o_272_sv2v_reg,data_o_271_sv2v_reg,
  data_o_270_sv2v_reg,data_o_269_sv2v_reg,data_o_268_sv2v_reg,data_o_267_sv2v_reg,
  data_o_266_sv2v_reg,data_o_265_sv2v_reg,data_o_264_sv2v_reg,data_o_263_sv2v_reg,
  data_o_262_sv2v_reg,data_o_261_sv2v_reg,data_o_260_sv2v_reg,data_o_259_sv2v_reg,
  data_o_258_sv2v_reg,data_o_257_sv2v_reg,data_o_256_sv2v_reg,data_o_255_sv2v_reg,
  data_o_254_sv2v_reg,data_o_253_sv2v_reg,data_o_252_sv2v_reg,data_o_251_sv2v_reg,
  data_o_250_sv2v_reg,data_o_249_sv2v_reg,data_o_248_sv2v_reg,data_o_247_sv2v_reg,
  data_o_246_sv2v_reg,data_o_245_sv2v_reg,data_o_244_sv2v_reg,data_o_243_sv2v_reg,
  data_o_242_sv2v_reg,data_o_241_sv2v_reg,data_o_240_sv2v_reg,data_o_239_sv2v_reg,
  data_o_238_sv2v_reg,data_o_237_sv2v_reg,data_o_236_sv2v_reg,data_o_235_sv2v_reg,
  data_o_234_sv2v_reg,data_o_233_sv2v_reg,data_o_232_sv2v_reg,data_o_231_sv2v_reg,
  data_o_230_sv2v_reg,data_o_229_sv2v_reg,data_o_228_sv2v_reg,data_o_227_sv2v_reg,
  data_o_226_sv2v_reg,data_o_225_sv2v_reg,data_o_224_sv2v_reg,data_o_223_sv2v_reg,
  data_o_222_sv2v_reg,data_o_221_sv2v_reg,data_o_220_sv2v_reg,data_o_219_sv2v_reg,
  data_o_218_sv2v_reg,data_o_217_sv2v_reg,data_o_216_sv2v_reg,data_o_215_sv2v_reg,
  data_o_214_sv2v_reg,data_o_213_sv2v_reg,data_o_212_sv2v_reg,data_o_211_sv2v_reg,
  data_o_210_sv2v_reg,data_o_209_sv2v_reg,data_o_208_sv2v_reg,data_o_207_sv2v_reg,
  data_o_206_sv2v_reg,data_o_205_sv2v_reg,data_o_204_sv2v_reg,data_o_203_sv2v_reg,
  data_o_202_sv2v_reg,data_o_201_sv2v_reg,data_o_200_sv2v_reg,data_o_199_sv2v_reg,
  data_o_198_sv2v_reg,data_o_197_sv2v_reg,data_o_196_sv2v_reg,data_o_195_sv2v_reg,
  data_o_194_sv2v_reg,data_o_193_sv2v_reg,data_o_192_sv2v_reg,data_o_191_sv2v_reg,
  data_o_190_sv2v_reg,data_o_189_sv2v_reg,data_o_188_sv2v_reg,data_o_187_sv2v_reg,
  data_o_186_sv2v_reg,data_o_185_sv2v_reg,data_o_184_sv2v_reg,data_o_183_sv2v_reg,
  data_o_182_sv2v_reg,data_o_181_sv2v_reg,data_o_180_sv2v_reg,data_o_179_sv2v_reg,
  data_o_178_sv2v_reg,data_o_177_sv2v_reg,data_o_176_sv2v_reg,data_o_175_sv2v_reg,
  data_o_174_sv2v_reg,data_o_173_sv2v_reg,data_o_172_sv2v_reg,data_o_171_sv2v_reg,
  data_o_170_sv2v_reg,data_o_169_sv2v_reg,data_o_168_sv2v_reg,data_o_167_sv2v_reg,
  data_o_166_sv2v_reg,data_o_165_sv2v_reg,data_o_164_sv2v_reg,data_o_163_sv2v_reg,
  data_o_162_sv2v_reg,data_o_161_sv2v_reg,data_o_160_sv2v_reg,data_o_159_sv2v_reg,
  data_o_158_sv2v_reg,data_o_157_sv2v_reg,data_o_156_sv2v_reg,data_o_155_sv2v_reg,
  data_o_154_sv2v_reg,data_o_153_sv2v_reg,data_o_152_sv2v_reg,data_o_151_sv2v_reg,
  data_o_150_sv2v_reg,data_o_149_sv2v_reg,data_o_148_sv2v_reg,data_o_147_sv2v_reg,
  data_o_146_sv2v_reg,data_o_145_sv2v_reg,data_o_144_sv2v_reg,data_o_143_sv2v_reg,
  data_o_142_sv2v_reg,data_o_141_sv2v_reg,data_o_140_sv2v_reg,data_o_139_sv2v_reg,
  data_o_138_sv2v_reg,data_o_137_sv2v_reg,data_o_136_sv2v_reg,data_o_135_sv2v_reg,
  data_o_134_sv2v_reg,data_o_133_sv2v_reg,data_o_132_sv2v_reg,data_o_131_sv2v_reg,
  data_o_130_sv2v_reg,data_o_129_sv2v_reg,data_o_128_sv2v_reg,data_o_127_sv2v_reg,
  data_o_126_sv2v_reg,data_o_125_sv2v_reg,data_o_124_sv2v_reg,data_o_123_sv2v_reg,
  data_o_122_sv2v_reg,data_o_121_sv2v_reg,data_o_120_sv2v_reg,data_o_119_sv2v_reg,
  data_o_118_sv2v_reg,data_o_117_sv2v_reg,data_o_116_sv2v_reg,data_o_115_sv2v_reg,
  data_o_114_sv2v_reg,data_o_113_sv2v_reg,data_o_112_sv2v_reg,data_o_111_sv2v_reg,
  data_o_110_sv2v_reg,data_o_109_sv2v_reg,data_o_108_sv2v_reg,data_o_107_sv2v_reg,
  data_o_106_sv2v_reg,data_o_105_sv2v_reg,data_o_104_sv2v_reg,data_o_103_sv2v_reg,
  data_o_102_sv2v_reg,data_o_101_sv2v_reg,data_o_100_sv2v_reg,data_o_99_sv2v_reg,
  data_o_98_sv2v_reg,data_o_97_sv2v_reg,data_o_96_sv2v_reg,data_o_95_sv2v_reg,
  data_o_94_sv2v_reg,data_o_93_sv2v_reg,data_o_92_sv2v_reg,data_o_91_sv2v_reg,
  data_o_90_sv2v_reg,data_o_89_sv2v_reg,data_o_88_sv2v_reg,data_o_87_sv2v_reg,
  data_o_86_sv2v_reg,data_o_85_sv2v_reg,data_o_84_sv2v_reg,data_o_83_sv2v_reg,
  data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,data_o_79_sv2v_reg,data_o_78_sv2v_reg,
  data_o_77_sv2v_reg,data_o_76_sv2v_reg,data_o_75_sv2v_reg,data_o_74_sv2v_reg,
  data_o_73_sv2v_reg,data_o_72_sv2v_reg,data_o_71_sv2v_reg,data_o_70_sv2v_reg,
  data_o_69_sv2v_reg,data_o_68_sv2v_reg,data_o_67_sv2v_reg,data_o_66_sv2v_reg,
  data_o_65_sv2v_reg,data_o_64_sv2v_reg,data_o_63_sv2v_reg,data_o_62_sv2v_reg,
  data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,data_o_58_sv2v_reg,data_o_57_sv2v_reg,
  data_o_56_sv2v_reg,data_o_55_sv2v_reg,data_o_54_sv2v_reg,data_o_53_sv2v_reg,
  data_o_52_sv2v_reg,data_o_51_sv2v_reg,data_o_50_sv2v_reg,data_o_49_sv2v_reg,
  data_o_48_sv2v_reg,data_o_47_sv2v_reg,data_o_46_sv2v_reg,data_o_45_sv2v_reg,
  data_o_44_sv2v_reg,data_o_43_sv2v_reg,data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,
  data_o_39_sv2v_reg,data_o_38_sv2v_reg,data_o_37_sv2v_reg,data_o_36_sv2v_reg,
  data_o_35_sv2v_reg,data_o_34_sv2v_reg,data_o_33_sv2v_reg,data_o_32_sv2v_reg,
  data_o_31_sv2v_reg,data_o_30_sv2v_reg,data_o_29_sv2v_reg,data_o_28_sv2v_reg,
  data_o_27_sv2v_reg,data_o_26_sv2v_reg,data_o_25_sv2v_reg,data_o_24_sv2v_reg,
  data_o_23_sv2v_reg,data_o_22_sv2v_reg,data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,
  data_o_18_sv2v_reg,data_o_17_sv2v_reg,data_o_16_sv2v_reg,data_o_15_sv2v_reg,
  data_o_14_sv2v_reg,data_o_13_sv2v_reg,data_o_12_sv2v_reg,data_o_11_sv2v_reg,
  data_o_10_sv2v_reg,data_o_9_sv2v_reg,data_o_8_sv2v_reg,data_o_7_sv2v_reg,
  data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,data_o_3_sv2v_reg,data_o_2_sv2v_reg,
  data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[294] = data_o_294_sv2v_reg;
  assign data_o[293] = data_o_293_sv2v_reg;
  assign data_o[292] = data_o_292_sv2v_reg;
  assign data_o[291] = data_o_291_sv2v_reg;
  assign data_o[290] = data_o_290_sv2v_reg;
  assign data_o[289] = data_o_289_sv2v_reg;
  assign data_o[288] = data_o_288_sv2v_reg;
  assign data_o[287] = data_o_287_sv2v_reg;
  assign data_o[286] = data_o_286_sv2v_reg;
  assign data_o[285] = data_o_285_sv2v_reg;
  assign data_o[284] = data_o_284_sv2v_reg;
  assign data_o[283] = data_o_283_sv2v_reg;
  assign data_o[282] = data_o_282_sv2v_reg;
  assign data_o[281] = data_o_281_sv2v_reg;
  assign data_o[280] = data_o_280_sv2v_reg;
  assign data_o[279] = data_o_279_sv2v_reg;
  assign data_o[278] = data_o_278_sv2v_reg;
  assign data_o[277] = data_o_277_sv2v_reg;
  assign data_o[276] = data_o_276_sv2v_reg;
  assign data_o[275] = data_o_275_sv2v_reg;
  assign data_o[274] = data_o_274_sv2v_reg;
  assign data_o[273] = data_o_273_sv2v_reg;
  assign data_o[272] = data_o_272_sv2v_reg;
  assign data_o[271] = data_o_271_sv2v_reg;
  assign data_o[270] = data_o_270_sv2v_reg;
  assign data_o[269] = data_o_269_sv2v_reg;
  assign data_o[268] = data_o_268_sv2v_reg;
  assign data_o[267] = data_o_267_sv2v_reg;
  assign data_o[266] = data_o_266_sv2v_reg;
  assign data_o[265] = data_o_265_sv2v_reg;
  assign data_o[264] = data_o_264_sv2v_reg;
  assign data_o[263] = data_o_263_sv2v_reg;
  assign data_o[262] = data_o_262_sv2v_reg;
  assign data_o[261] = data_o_261_sv2v_reg;
  assign data_o[260] = data_o_260_sv2v_reg;
  assign data_o[259] = data_o_259_sv2v_reg;
  assign data_o[258] = data_o_258_sv2v_reg;
  assign data_o[257] = data_o_257_sv2v_reg;
  assign data_o[256] = data_o_256_sv2v_reg;
  assign data_o[255] = data_o_255_sv2v_reg;
  assign data_o[254] = data_o_254_sv2v_reg;
  assign data_o[253] = data_o_253_sv2v_reg;
  assign data_o[252] = data_o_252_sv2v_reg;
  assign data_o[251] = data_o_251_sv2v_reg;
  assign data_o[250] = data_o_250_sv2v_reg;
  assign data_o[249] = data_o_249_sv2v_reg;
  assign data_o[248] = data_o_248_sv2v_reg;
  assign data_o[247] = data_o_247_sv2v_reg;
  assign data_o[246] = data_o_246_sv2v_reg;
  assign data_o[245] = data_o_245_sv2v_reg;
  assign data_o[244] = data_o_244_sv2v_reg;
  assign data_o[243] = data_o_243_sv2v_reg;
  assign data_o[242] = data_o_242_sv2v_reg;
  assign data_o[241] = data_o_241_sv2v_reg;
  assign data_o[240] = data_o_240_sv2v_reg;
  assign data_o[239] = data_o_239_sv2v_reg;
  assign data_o[238] = data_o_238_sv2v_reg;
  assign data_o[237] = data_o_237_sv2v_reg;
  assign data_o[236] = data_o_236_sv2v_reg;
  assign data_o[235] = data_o_235_sv2v_reg;
  assign data_o[234] = data_o_234_sv2v_reg;
  assign data_o[233] = data_o_233_sv2v_reg;
  assign data_o[232] = data_o_232_sv2v_reg;
  assign data_o[231] = data_o_231_sv2v_reg;
  assign data_o[230] = data_o_230_sv2v_reg;
  assign data_o[229] = data_o_229_sv2v_reg;
  assign data_o[228] = data_o_228_sv2v_reg;
  assign data_o[227] = data_o_227_sv2v_reg;
  assign data_o[226] = data_o_226_sv2v_reg;
  assign data_o[225] = data_o_225_sv2v_reg;
  assign data_o[224] = data_o_224_sv2v_reg;
  assign data_o[223] = data_o_223_sv2v_reg;
  assign data_o[222] = data_o_222_sv2v_reg;
  assign data_o[221] = data_o_221_sv2v_reg;
  assign data_o[220] = data_o_220_sv2v_reg;
  assign data_o[219] = data_o_219_sv2v_reg;
  assign data_o[218] = data_o_218_sv2v_reg;
  assign data_o[217] = data_o_217_sv2v_reg;
  assign data_o[216] = data_o_216_sv2v_reg;
  assign data_o[215] = data_o_215_sv2v_reg;
  assign data_o[214] = data_o_214_sv2v_reg;
  assign data_o[213] = data_o_213_sv2v_reg;
  assign data_o[212] = data_o_212_sv2v_reg;
  assign data_o[211] = data_o_211_sv2v_reg;
  assign data_o[210] = data_o_210_sv2v_reg;
  assign data_o[209] = data_o_209_sv2v_reg;
  assign data_o[208] = data_o_208_sv2v_reg;
  assign data_o[207] = data_o_207_sv2v_reg;
  assign data_o[206] = data_o_206_sv2v_reg;
  assign data_o[205] = data_o_205_sv2v_reg;
  assign data_o[204] = data_o_204_sv2v_reg;
  assign data_o[203] = data_o_203_sv2v_reg;
  assign data_o[202] = data_o_202_sv2v_reg;
  assign data_o[201] = data_o_201_sv2v_reg;
  assign data_o[200] = data_o_200_sv2v_reg;
  assign data_o[199] = data_o_199_sv2v_reg;
  assign data_o[198] = data_o_198_sv2v_reg;
  assign data_o[197] = data_o_197_sv2v_reg;
  assign data_o[196] = data_o_196_sv2v_reg;
  assign data_o[195] = data_o_195_sv2v_reg;
  assign data_o[194] = data_o_194_sv2v_reg;
  assign data_o[193] = data_o_193_sv2v_reg;
  assign data_o[192] = data_o_192_sv2v_reg;
  assign data_o[191] = data_o_191_sv2v_reg;
  assign data_o[190] = data_o_190_sv2v_reg;
  assign data_o[189] = data_o_189_sv2v_reg;
  assign data_o[188] = data_o_188_sv2v_reg;
  assign data_o[187] = data_o_187_sv2v_reg;
  assign data_o[186] = data_o_186_sv2v_reg;
  assign data_o[185] = data_o_185_sv2v_reg;
  assign data_o[184] = data_o_184_sv2v_reg;
  assign data_o[183] = data_o_183_sv2v_reg;
  assign data_o[182] = data_o_182_sv2v_reg;
  assign data_o[181] = data_o_181_sv2v_reg;
  assign data_o[180] = data_o_180_sv2v_reg;
  assign data_o[179] = data_o_179_sv2v_reg;
  assign data_o[178] = data_o_178_sv2v_reg;
  assign data_o[177] = data_o_177_sv2v_reg;
  assign data_o[176] = data_o_176_sv2v_reg;
  assign data_o[175] = data_o_175_sv2v_reg;
  assign data_o[174] = data_o_174_sv2v_reg;
  assign data_o[173] = data_o_173_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_294_sv2v_reg <= data_i[294];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_293_sv2v_reg <= data_i[293];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_292_sv2v_reg <= data_i[292];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_291_sv2v_reg <= data_i[291];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_290_sv2v_reg <= data_i[290];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_289_sv2v_reg <= data_i[289];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_288_sv2v_reg <= data_i[288];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_287_sv2v_reg <= data_i[287];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_286_sv2v_reg <= data_i[286];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_285_sv2v_reg <= data_i[285];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_284_sv2v_reg <= data_i[284];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_283_sv2v_reg <= data_i[283];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_282_sv2v_reg <= data_i[282];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_281_sv2v_reg <= data_i[281];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_280_sv2v_reg <= data_i[280];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_279_sv2v_reg <= data_i[279];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_278_sv2v_reg <= data_i[278];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_277_sv2v_reg <= data_i[277];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_276_sv2v_reg <= data_i[276];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_275_sv2v_reg <= data_i[275];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_274_sv2v_reg <= data_i[274];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_273_sv2v_reg <= data_i[273];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_272_sv2v_reg <= data_i[272];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_271_sv2v_reg <= data_i[271];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_270_sv2v_reg <= data_i[270];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_269_sv2v_reg <= data_i[269];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_268_sv2v_reg <= data_i[268];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_267_sv2v_reg <= data_i[267];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_266_sv2v_reg <= data_i[266];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_265_sv2v_reg <= data_i[265];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_264_sv2v_reg <= data_i[264];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_263_sv2v_reg <= data_i[263];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_262_sv2v_reg <= data_i[262];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_261_sv2v_reg <= data_i[261];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_260_sv2v_reg <= data_i[260];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_259_sv2v_reg <= data_i[259];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_258_sv2v_reg <= data_i[258];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_257_sv2v_reg <= data_i[257];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_256_sv2v_reg <= data_i[256];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_255_sv2v_reg <= data_i[255];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_254_sv2v_reg <= data_i[254];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_253_sv2v_reg <= data_i[253];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_252_sv2v_reg <= data_i[252];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_251_sv2v_reg <= data_i[251];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_250_sv2v_reg <= data_i[250];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_249_sv2v_reg <= data_i[249];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_248_sv2v_reg <= data_i[248];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_247_sv2v_reg <= data_i[247];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_246_sv2v_reg <= data_i[246];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_245_sv2v_reg <= data_i[245];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_244_sv2v_reg <= data_i[244];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_243_sv2v_reg <= data_i[243];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_242_sv2v_reg <= data_i[242];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_241_sv2v_reg <= data_i[241];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_240_sv2v_reg <= data_i[240];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_239_sv2v_reg <= data_i[239];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_238_sv2v_reg <= data_i[238];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_237_sv2v_reg <= data_i[237];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_236_sv2v_reg <= data_i[236];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_235_sv2v_reg <= data_i[235];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_234_sv2v_reg <= data_i[234];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_233_sv2v_reg <= data_i[233];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_232_sv2v_reg <= data_i[232];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_231_sv2v_reg <= data_i[231];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_230_sv2v_reg <= data_i[230];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_229_sv2v_reg <= data_i[229];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_228_sv2v_reg <= data_i[228];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_227_sv2v_reg <= data_i[227];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_226_sv2v_reg <= data_i[226];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_225_sv2v_reg <= data_i[225];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_224_sv2v_reg <= data_i[224];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_223_sv2v_reg <= data_i[223];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_222_sv2v_reg <= data_i[222];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_221_sv2v_reg <= data_i[221];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_220_sv2v_reg <= data_i[220];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_219_sv2v_reg <= data_i[219];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_218_sv2v_reg <= data_i[218];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_217_sv2v_reg <= data_i[217];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_216_sv2v_reg <= data_i[216];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_215_sv2v_reg <= data_i[215];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_214_sv2v_reg <= data_i[214];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_213_sv2v_reg <= data_i[213];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_212_sv2v_reg <= data_i[212];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_211_sv2v_reg <= data_i[211];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_210_sv2v_reg <= data_i[210];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_209_sv2v_reg <= data_i[209];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_208_sv2v_reg <= data_i[208];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_207_sv2v_reg <= data_i[207];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_206_sv2v_reg <= data_i[206];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_205_sv2v_reg <= data_i[205];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_204_sv2v_reg <= data_i[204];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_203_sv2v_reg <= data_i[203];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_202_sv2v_reg <= data_i[202];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_201_sv2v_reg <= data_i[201];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_200_sv2v_reg <= data_i[200];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_199_sv2v_reg <= data_i[199];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_198_sv2v_reg <= data_i[198];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_197_sv2v_reg <= data_i[197];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_196_sv2v_reg <= data_i[196];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_195_sv2v_reg <= data_i[195];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_194_sv2v_reg <= data_i[194];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_193_sv2v_reg <= data_i[193];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_192_sv2v_reg <= data_i[192];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_191_sv2v_reg <= data_i[191];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_190_sv2v_reg <= data_i[190];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_189_sv2v_reg <= data_i[189];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_188_sv2v_reg <= data_i[188];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_187_sv2v_reg <= data_i[187];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_186_sv2v_reg <= data_i[186];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_185_sv2v_reg <= data_i[185];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_184_sv2v_reg <= data_i[184];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_183_sv2v_reg <= data_i[183];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_182_sv2v_reg <= data_i[182];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_181_sv2v_reg <= data_i[181];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_180_sv2v_reg <= data_i[180];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_179_sv2v_reg <= data_i[179];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_178_sv2v_reg <= data_i[178];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_177_sv2v_reg <= data_i[177];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_176_sv2v_reg <= data_i[176];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_175_sv2v_reg <= data_i[175];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_174_sv2v_reg <= data_i[174];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_173_sv2v_reg <= data_i[173];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_172_sv2v_reg <= data_i[172];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_171_sv2v_reg <= data_i[171];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_170_sv2v_reg <= data_i[170];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_169_sv2v_reg <= data_i[169];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_168_sv2v_reg <= data_i[168];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_167_sv2v_reg <= data_i[167];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_166_sv2v_reg <= data_i[166];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_165_sv2v_reg <= data_i[165];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_164_sv2v_reg <= data_i[164];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_163_sv2v_reg <= data_i[163];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_162_sv2v_reg <= data_i[162];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_161_sv2v_reg <= data_i[161];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_160_sv2v_reg <= data_i[160];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_159_sv2v_reg <= data_i[159];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_158_sv2v_reg <= data_i[158];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_157_sv2v_reg <= data_i[157];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_156_sv2v_reg <= data_i[156];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_155_sv2v_reg <= data_i[155];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_154_sv2v_reg <= data_i[154];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_153_sv2v_reg <= data_i[153];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_152_sv2v_reg <= data_i[152];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_151_sv2v_reg <= data_i[151];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_150_sv2v_reg <= data_i[150];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_149_sv2v_reg <= data_i[149];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_148_sv2v_reg <= data_i[148];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_147_sv2v_reg <= data_i[147];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_146_sv2v_reg <= data_i[146];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_145_sv2v_reg <= data_i[145];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_144_sv2v_reg <= data_i[144];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_143_sv2v_reg <= data_i[143];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_142_sv2v_reg <= data_i[142];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_141_sv2v_reg <= data_i[141];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_140_sv2v_reg <= data_i[140];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_139_sv2v_reg <= data_i[139];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_138_sv2v_reg <= data_i[138];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_137_sv2v_reg <= data_i[137];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_136_sv2v_reg <= data_i[136];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_135_sv2v_reg <= data_i[135];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_134_sv2v_reg <= data_i[134];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_133_sv2v_reg <= data_i[133];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_132_sv2v_reg <= data_i[132];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_131_sv2v_reg <= data_i[131];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_130_sv2v_reg <= data_i[130];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_129_sv2v_reg <= data_i[129];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_128_sv2v_reg <= data_i[128];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_127_sv2v_reg <= data_i[127];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_126_sv2v_reg <= data_i[126];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_125_sv2v_reg <= data_i[125];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_124_sv2v_reg <= data_i[124];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_123_sv2v_reg <= data_i[123];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_122_sv2v_reg <= data_i[122];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_121_sv2v_reg <= data_i[121];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_120_sv2v_reg <= data_i[120];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_119_sv2v_reg <= data_i[119];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_118_sv2v_reg <= data_i[118];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_117_sv2v_reg <= data_i[117];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_116_sv2v_reg <= data_i[116];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_115_sv2v_reg <= data_i[115];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_114_sv2v_reg <= data_i[114];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_113_sv2v_reg <= data_i[113];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_112_sv2v_reg <= data_i[112];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_111_sv2v_reg <= data_i[111];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_110_sv2v_reg <= data_i[110];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_109_sv2v_reg <= data_i[109];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_108_sv2v_reg <= data_i[108];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_107_sv2v_reg <= data_i[107];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_106_sv2v_reg <= data_i[106];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_105_sv2v_reg <= data_i[105];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_104_sv2v_reg <= data_i[104];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_103_sv2v_reg <= data_i[103];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_102_sv2v_reg <= data_i[102];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_101_sv2v_reg <= data_i[101];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_100_sv2v_reg <= data_i[100];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_99_sv2v_reg <= data_i[99];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_98_sv2v_reg <= data_i[98];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_97_sv2v_reg <= data_i[97];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_96_sv2v_reg <= data_i[96];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_95_sv2v_reg <= data_i[95];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_94_sv2v_reg <= data_i[94];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_93_sv2v_reg <= data_i[93];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_92_sv2v_reg <= data_i[92];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_91_sv2v_reg <= data_i[91];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_90_sv2v_reg <= data_i[90];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_89_sv2v_reg <= data_i[89];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_88_sv2v_reg <= data_i[88];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_87_sv2v_reg <= data_i[87];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_86_sv2v_reg <= data_i[86];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_85_sv2v_reg <= data_i[85];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_84_sv2v_reg <= data_i[84];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_83_sv2v_reg <= data_i[83];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_82_sv2v_reg <= data_i[82];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_81_sv2v_reg <= data_i[81];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_80_sv2v_reg <= data_i[80];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_79_sv2v_reg <= data_i[79];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_78_sv2v_reg <= data_i[78];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_77_sv2v_reg <= data_i[77];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_76_sv2v_reg <= data_i[76];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_75_sv2v_reg <= data_i[75];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_74_sv2v_reg <= data_i[74];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_73_sv2v_reg <= data_i[73];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_72_sv2v_reg <= data_i[72];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_71_sv2v_reg <= data_i[71];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_70_sv2v_reg <= data_i[70];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_69_sv2v_reg <= data_i[69];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_68_sv2v_reg <= data_i[68];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_67_sv2v_reg <= data_i[67];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_66_sv2v_reg <= data_i[66];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_65_sv2v_reg <= data_i[65];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_64_sv2v_reg <= data_i[64];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_63_sv2v_reg <= data_i[63];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_62_sv2v_reg <= data_i[62];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_61_sv2v_reg <= data_i[61];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_60_sv2v_reg <= data_i[60];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_59_sv2v_reg <= data_i[59];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_58_sv2v_reg <= data_i[58];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_57_sv2v_reg <= data_i[57];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_56_sv2v_reg <= data_i[56];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_55_sv2v_reg <= data_i[55];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_54_sv2v_reg <= data_i[54];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_53_sv2v_reg <= data_i[53];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_52_sv2v_reg <= data_i[52];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_51_sv2v_reg <= data_i[51];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_50_sv2v_reg <= data_i[50];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_49_sv2v_reg <= data_i[49];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_48_sv2v_reg <= data_i[48];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_47_sv2v_reg <= data_i[47];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_46_sv2v_reg <= data_i[46];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_45_sv2v_reg <= data_i[45];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_44_sv2v_reg <= data_i[44];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_43_sv2v_reg <= data_i[43];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_42_sv2v_reg <= data_i[42];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_41_sv2v_reg <= data_i[41];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_40_sv2v_reg <= data_i[40];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_39_sv2v_reg <= data_i[39];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_38_sv2v_reg <= data_i[38];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_37_sv2v_reg <= data_i[37];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_36_sv2v_reg <= data_i[36];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_35_sv2v_reg <= data_i[35];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_34_sv2v_reg <= data_i[34];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_33_sv2v_reg <= data_i[33];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_32_sv2v_reg <= data_i[32];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_31_sv2v_reg <= data_i[31];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_30_sv2v_reg <= data_i[30];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_29_sv2v_reg <= data_i[29];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_28_sv2v_reg <= data_i[28];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_27_sv2v_reg <= data_i[27];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_26_sv2v_reg <= data_i[26];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_25_sv2v_reg <= data_i[25];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_24_sv2v_reg <= data_i[24];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_23_sv2v_reg <= data_i[23];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_22_sv2v_reg <= data_i[22];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_21_sv2v_reg <= data_i[21];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_20_sv2v_reg <= data_i[20];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_19_sv2v_reg <= data_i[19];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_18_sv2v_reg <= data_i[18];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_17_sv2v_reg <= data_i[17];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_16_sv2v_reg <= data_i[16];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_15_sv2v_reg <= data_i[15];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_14_sv2v_reg <= data_i[14];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_13_sv2v_reg <= data_i[13];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_12_sv2v_reg <= data_i[12];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_11_sv2v_reg <= data_i[11];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_10_sv2v_reg <= data_i[10];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_9_sv2v_reg <= data_i[9];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_8_sv2v_reg <= data_i[8];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_7_sv2v_reg <= data_i[7];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_6_sv2v_reg <= data_i[6];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_5_sv2v_reg <= data_i[5];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_4_sv2v_reg <= data_i[4];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_3_sv2v_reg <= data_i[3];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_2_sv2v_reg <= data_i[2];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_1_sv2v_reg <= data_i[1];
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      data_o_0_sv2v_reg <= data_i[0];
    end 
  end


endmodule