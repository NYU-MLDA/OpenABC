module bsg_mesh_stitch_width_p64_x_max_p2_y_max_p1
(
  outs_i,
  ins_o,
  hor_i,
  hor_o,
  ver_i,
  ver_o
);

  input [511:0] outs_i;
  output [511:0] ins_o;
  input [127:0] hor_i;
  output [127:0] hor_o;
  input [255:0] ver_i;
  output [255:0] ver_o;
  wire [511:0] ins_o;
  wire [127:0] hor_o;
  wire [255:0] ver_o;
  assign ins_o[511] = ver_i[255];
  assign ins_o[510] = ver_i[254];
  assign ins_o[509] = ver_i[253];
  assign ins_o[508] = ver_i[252];
  assign ins_o[507] = ver_i[251];
  assign ins_o[506] = ver_i[250];
  assign ins_o[505] = ver_i[249];
  assign ins_o[504] = ver_i[248];
  assign ins_o[503] = ver_i[247];
  assign ins_o[502] = ver_i[246];
  assign ins_o[501] = ver_i[245];
  assign ins_o[500] = ver_i[244];
  assign ins_o[499] = ver_i[243];
  assign ins_o[498] = ver_i[242];
  assign ins_o[497] = ver_i[241];
  assign ins_o[496] = ver_i[240];
  assign ins_o[495] = ver_i[239];
  assign ins_o[494] = ver_i[238];
  assign ins_o[493] = ver_i[237];
  assign ins_o[492] = ver_i[236];
  assign ins_o[491] = ver_i[235];
  assign ins_o[490] = ver_i[234];
  assign ins_o[489] = ver_i[233];
  assign ins_o[488] = ver_i[232];
  assign ins_o[487] = ver_i[231];
  assign ins_o[486] = ver_i[230];
  assign ins_o[485] = ver_i[229];
  assign ins_o[484] = ver_i[228];
  assign ins_o[483] = ver_i[227];
  assign ins_o[482] = ver_i[226];
  assign ins_o[481] = ver_i[225];
  assign ins_o[480] = ver_i[224];
  assign ins_o[479] = ver_i[223];
  assign ins_o[478] = ver_i[222];
  assign ins_o[477] = ver_i[221];
  assign ins_o[476] = ver_i[220];
  assign ins_o[475] = ver_i[219];
  assign ins_o[474] = ver_i[218];
  assign ins_o[473] = ver_i[217];
  assign ins_o[472] = ver_i[216];
  assign ins_o[471] = ver_i[215];
  assign ins_o[470] = ver_i[214];
  assign ins_o[469] = ver_i[213];
  assign ins_o[468] = ver_i[212];
  assign ins_o[467] = ver_i[211];
  assign ins_o[466] = ver_i[210];
  assign ins_o[465] = ver_i[209];
  assign ins_o[464] = ver_i[208];
  assign ins_o[463] = ver_i[207];
  assign ins_o[462] = ver_i[206];
  assign ins_o[461] = ver_i[205];
  assign ins_o[460] = ver_i[204];
  assign ins_o[459] = ver_i[203];
  assign ins_o[458] = ver_i[202];
  assign ins_o[457] = ver_i[201];
  assign ins_o[456] = ver_i[200];
  assign ins_o[455] = ver_i[199];
  assign ins_o[454] = ver_i[198];
  assign ins_o[453] = ver_i[197];
  assign ins_o[452] = ver_i[196];
  assign ins_o[451] = ver_i[195];
  assign ins_o[450] = ver_i[194];
  assign ins_o[449] = ver_i[193];
  assign ins_o[448] = ver_i[192];
  assign ins_o[447] = ver_i[127];
  assign ins_o[446] = ver_i[126];
  assign ins_o[445] = ver_i[125];
  assign ins_o[444] = ver_i[124];
  assign ins_o[443] = ver_i[123];
  assign ins_o[442] = ver_i[122];
  assign ins_o[441] = ver_i[121];
  assign ins_o[440] = ver_i[120];
  assign ins_o[439] = ver_i[119];
  assign ins_o[438] = ver_i[118];
  assign ins_o[437] = ver_i[117];
  assign ins_o[436] = ver_i[116];
  assign ins_o[435] = ver_i[115];
  assign ins_o[434] = ver_i[114];
  assign ins_o[433] = ver_i[113];
  assign ins_o[432] = ver_i[112];
  assign ins_o[431] = ver_i[111];
  assign ins_o[430] = ver_i[110];
  assign ins_o[429] = ver_i[109];
  assign ins_o[428] = ver_i[108];
  assign ins_o[427] = ver_i[107];
  assign ins_o[426] = ver_i[106];
  assign ins_o[425] = ver_i[105];
  assign ins_o[424] = ver_i[104];
  assign ins_o[423] = ver_i[103];
  assign ins_o[422] = ver_i[102];
  assign ins_o[421] = ver_i[101];
  assign ins_o[420] = ver_i[100];
  assign ins_o[419] = ver_i[99];
  assign ins_o[418] = ver_i[98];
  assign ins_o[417] = ver_i[97];
  assign ins_o[416] = ver_i[96];
  assign ins_o[415] = ver_i[95];
  assign ins_o[414] = ver_i[94];
  assign ins_o[413] = ver_i[93];
  assign ins_o[412] = ver_i[92];
  assign ins_o[411] = ver_i[91];
  assign ins_o[410] = ver_i[90];
  assign ins_o[409] = ver_i[89];
  assign ins_o[408] = ver_i[88];
  assign ins_o[407] = ver_i[87];
  assign ins_o[406] = ver_i[86];
  assign ins_o[405] = ver_i[85];
  assign ins_o[404] = ver_i[84];
  assign ins_o[403] = ver_i[83];
  assign ins_o[402] = ver_i[82];
  assign ins_o[401] = ver_i[81];
  assign ins_o[400] = ver_i[80];
  assign ins_o[399] = ver_i[79];
  assign ins_o[398] = ver_i[78];
  assign ins_o[397] = ver_i[77];
  assign ins_o[396] = ver_i[76];
  assign ins_o[395] = ver_i[75];
  assign ins_o[394] = ver_i[74];
  assign ins_o[393] = ver_i[73];
  assign ins_o[392] = ver_i[72];
  assign ins_o[391] = ver_i[71];
  assign ins_o[390] = ver_i[70];
  assign ins_o[389] = ver_i[69];
  assign ins_o[388] = ver_i[68];
  assign ins_o[387] = ver_i[67];
  assign ins_o[386] = ver_i[66];
  assign ins_o[385] = ver_i[65];
  assign ins_o[384] = ver_i[64];
  assign ins_o[383] = hor_i[127];
  assign ins_o[382] = hor_i[126];
  assign ins_o[381] = hor_i[125];
  assign ins_o[380] = hor_i[124];
  assign ins_o[379] = hor_i[123];
  assign ins_o[378] = hor_i[122];
  assign ins_o[377] = hor_i[121];
  assign ins_o[376] = hor_i[120];
  assign ins_o[375] = hor_i[119];
  assign ins_o[374] = hor_i[118];
  assign ins_o[373] = hor_i[117];
  assign ins_o[372] = hor_i[116];
  assign ins_o[371] = hor_i[115];
  assign ins_o[370] = hor_i[114];
  assign ins_o[369] = hor_i[113];
  assign ins_o[368] = hor_i[112];
  assign ins_o[367] = hor_i[111];
  assign ins_o[366] = hor_i[110];
  assign ins_o[365] = hor_i[109];
  assign ins_o[364] = hor_i[108];
  assign ins_o[363] = hor_i[107];
  assign ins_o[362] = hor_i[106];
  assign ins_o[361] = hor_i[105];
  assign ins_o[360] = hor_i[104];
  assign ins_o[359] = hor_i[103];
  assign ins_o[358] = hor_i[102];
  assign ins_o[357] = hor_i[101];
  assign ins_o[356] = hor_i[100];
  assign ins_o[355] = hor_i[99];
  assign ins_o[354] = hor_i[98];
  assign ins_o[353] = hor_i[97];
  assign ins_o[352] = hor_i[96];
  assign ins_o[351] = hor_i[95];
  assign ins_o[350] = hor_i[94];
  assign ins_o[349] = hor_i[93];
  assign ins_o[348] = hor_i[92];
  assign ins_o[347] = hor_i[91];
  assign ins_o[346] = hor_i[90];
  assign ins_o[345] = hor_i[89];
  assign ins_o[344] = hor_i[88];
  assign ins_o[343] = hor_i[87];
  assign ins_o[342] = hor_i[86];
  assign ins_o[341] = hor_i[85];
  assign ins_o[340] = hor_i[84];
  assign ins_o[339] = hor_i[83];
  assign ins_o[338] = hor_i[82];
  assign ins_o[337] = hor_i[81];
  assign ins_o[336] = hor_i[80];
  assign ins_o[335] = hor_i[79];
  assign ins_o[334] = hor_i[78];
  assign ins_o[333] = hor_i[77];
  assign ins_o[332] = hor_i[76];
  assign ins_o[331] = hor_i[75];
  assign ins_o[330] = hor_i[74];
  assign ins_o[329] = hor_i[73];
  assign ins_o[328] = hor_i[72];
  assign ins_o[327] = hor_i[71];
  assign ins_o[326] = hor_i[70];
  assign ins_o[325] = hor_i[69];
  assign ins_o[324] = hor_i[68];
  assign ins_o[323] = hor_i[67];
  assign ins_o[322] = hor_i[66];
  assign ins_o[321] = hor_i[65];
  assign ins_o[320] = hor_i[64];
  assign ins_o[319] = outs_i[127];
  assign ins_o[318] = outs_i[126];
  assign ins_o[317] = outs_i[125];
  assign ins_o[316] = outs_i[124];
  assign ins_o[315] = outs_i[123];
  assign ins_o[314] = outs_i[122];
  assign ins_o[313] = outs_i[121];
  assign ins_o[312] = outs_i[120];
  assign ins_o[311] = outs_i[119];
  assign ins_o[310] = outs_i[118];
  assign ins_o[309] = outs_i[117];
  assign ins_o[308] = outs_i[116];
  assign ins_o[307] = outs_i[115];
  assign ins_o[306] = outs_i[114];
  assign ins_o[305] = outs_i[113];
  assign ins_o[304] = outs_i[112];
  assign ins_o[303] = outs_i[111];
  assign ins_o[302] = outs_i[110];
  assign ins_o[301] = outs_i[109];
  assign ins_o[300] = outs_i[108];
  assign ins_o[299] = outs_i[107];
  assign ins_o[298] = outs_i[106];
  assign ins_o[297] = outs_i[105];
  assign ins_o[296] = outs_i[104];
  assign ins_o[295] = outs_i[103];
  assign ins_o[294] = outs_i[102];
  assign ins_o[293] = outs_i[101];
  assign ins_o[292] = outs_i[100];
  assign ins_o[291] = outs_i[99];
  assign ins_o[290] = outs_i[98];
  assign ins_o[289] = outs_i[97];
  assign ins_o[288] = outs_i[96];
  assign ins_o[287] = outs_i[95];
  assign ins_o[286] = outs_i[94];
  assign ins_o[285] = outs_i[93];
  assign ins_o[284] = outs_i[92];
  assign ins_o[283] = outs_i[91];
  assign ins_o[282] = outs_i[90];
  assign ins_o[281] = outs_i[89];
  assign ins_o[280] = outs_i[88];
  assign ins_o[279] = outs_i[87];
  assign ins_o[278] = outs_i[86];
  assign ins_o[277] = outs_i[85];
  assign ins_o[276] = outs_i[84];
  assign ins_o[275] = outs_i[83];
  assign ins_o[274] = outs_i[82];
  assign ins_o[273] = outs_i[81];
  assign ins_o[272] = outs_i[80];
  assign ins_o[271] = outs_i[79];
  assign ins_o[270] = outs_i[78];
  assign ins_o[269] = outs_i[77];
  assign ins_o[268] = outs_i[76];
  assign ins_o[267] = outs_i[75];
  assign ins_o[266] = outs_i[74];
  assign ins_o[265] = outs_i[73];
  assign ins_o[264] = outs_i[72];
  assign ins_o[263] = outs_i[71];
  assign ins_o[262] = outs_i[70];
  assign ins_o[261] = outs_i[69];
  assign ins_o[260] = outs_i[68];
  assign ins_o[259] = outs_i[67];
  assign ins_o[258] = outs_i[66];
  assign ins_o[257] = outs_i[65];
  assign ins_o[256] = outs_i[64];
  assign ins_o[255] = ver_i[191];
  assign ins_o[254] = ver_i[190];
  assign ins_o[253] = ver_i[189];
  assign ins_o[252] = ver_i[188];
  assign ins_o[251] = ver_i[187];
  assign ins_o[250] = ver_i[186];
  assign ins_o[249] = ver_i[185];
  assign ins_o[248] = ver_i[184];
  assign ins_o[247] = ver_i[183];
  assign ins_o[246] = ver_i[182];
  assign ins_o[245] = ver_i[181];
  assign ins_o[244] = ver_i[180];
  assign ins_o[243] = ver_i[179];
  assign ins_o[242] = ver_i[178];
  assign ins_o[241] = ver_i[177];
  assign ins_o[240] = ver_i[176];
  assign ins_o[239] = ver_i[175];
  assign ins_o[238] = ver_i[174];
  assign ins_o[237] = ver_i[173];
  assign ins_o[236] = ver_i[172];
  assign ins_o[235] = ver_i[171];
  assign ins_o[234] = ver_i[170];
  assign ins_o[233] = ver_i[169];
  assign ins_o[232] = ver_i[168];
  assign ins_o[231] = ver_i[167];
  assign ins_o[230] = ver_i[166];
  assign ins_o[229] = ver_i[165];
  assign ins_o[228] = ver_i[164];
  assign ins_o[227] = ver_i[163];
  assign ins_o[226] = ver_i[162];
  assign ins_o[225] = ver_i[161];
  assign ins_o[224] = ver_i[160];
  assign ins_o[223] = ver_i[159];
  assign ins_o[222] = ver_i[158];
  assign ins_o[221] = ver_i[157];
  assign ins_o[220] = ver_i[156];
  assign ins_o[219] = ver_i[155];
  assign ins_o[218] = ver_i[154];
  assign ins_o[217] = ver_i[153];
  assign ins_o[216] = ver_i[152];
  assign ins_o[215] = ver_i[151];
  assign ins_o[214] = ver_i[150];
  assign ins_o[213] = ver_i[149];
  assign ins_o[212] = ver_i[148];
  assign ins_o[211] = ver_i[147];
  assign ins_o[210] = ver_i[146];
  assign ins_o[209] = ver_i[145];
  assign ins_o[208] = ver_i[144];
  assign ins_o[207] = ver_i[143];
  assign ins_o[206] = ver_i[142];
  assign ins_o[205] = ver_i[141];
  assign ins_o[204] = ver_i[140];
  assign ins_o[203] = ver_i[139];
  assign ins_o[202] = ver_i[138];
  assign ins_o[201] = ver_i[137];
  assign ins_o[200] = ver_i[136];
  assign ins_o[199] = ver_i[135];
  assign ins_o[198] = ver_i[134];
  assign ins_o[197] = ver_i[133];
  assign ins_o[196] = ver_i[132];
  assign ins_o[195] = ver_i[131];
  assign ins_o[194] = ver_i[130];
  assign ins_o[193] = ver_i[129];
  assign ins_o[192] = ver_i[128];
  assign ins_o[191] = ver_i[63];
  assign ins_o[190] = ver_i[62];
  assign ins_o[189] = ver_i[61];
  assign ins_o[188] = ver_i[60];
  assign ins_o[187] = ver_i[59];
  assign ins_o[186] = ver_i[58];
  assign ins_o[185] = ver_i[57];
  assign ins_o[184] = ver_i[56];
  assign ins_o[183] = ver_i[55];
  assign ins_o[182] = ver_i[54];
  assign ins_o[181] = ver_i[53];
  assign ins_o[180] = ver_i[52];
  assign ins_o[179] = ver_i[51];
  assign ins_o[178] = ver_i[50];
  assign ins_o[177] = ver_i[49];
  assign ins_o[176] = ver_i[48];
  assign ins_o[175] = ver_i[47];
  assign ins_o[174] = ver_i[46];
  assign ins_o[173] = ver_i[45];
  assign ins_o[172] = ver_i[44];
  assign ins_o[171] = ver_i[43];
  assign ins_o[170] = ver_i[42];
  assign ins_o[169] = ver_i[41];
  assign ins_o[168] = ver_i[40];
  assign ins_o[167] = ver_i[39];
  assign ins_o[166] = ver_i[38];
  assign ins_o[165] = ver_i[37];
  assign ins_o[164] = ver_i[36];
  assign ins_o[163] = ver_i[35];
  assign ins_o[162] = ver_i[34];
  assign ins_o[161] = ver_i[33];
  assign ins_o[160] = ver_i[32];
  assign ins_o[159] = ver_i[31];
  assign ins_o[158] = ver_i[30];
  assign ins_o[157] = ver_i[29];
  assign ins_o[156] = ver_i[28];
  assign ins_o[155] = ver_i[27];
  assign ins_o[154] = ver_i[26];
  assign ins_o[153] = ver_i[25];
  assign ins_o[152] = ver_i[24];
  assign ins_o[151] = ver_i[23];
  assign ins_o[150] = ver_i[22];
  assign ins_o[149] = ver_i[21];
  assign ins_o[148] = ver_i[20];
  assign ins_o[147] = ver_i[19];
  assign ins_o[146] = ver_i[18];
  assign ins_o[145] = ver_i[17];
  assign ins_o[144] = ver_i[16];
  assign ins_o[143] = ver_i[15];
  assign ins_o[142] = ver_i[14];
  assign ins_o[141] = ver_i[13];
  assign ins_o[140] = ver_i[12];
  assign ins_o[139] = ver_i[11];
  assign ins_o[138] = ver_i[10];
  assign ins_o[137] = ver_i[9];
  assign ins_o[136] = ver_i[8];
  assign ins_o[135] = ver_i[7];
  assign ins_o[134] = ver_i[6];
  assign ins_o[133] = ver_i[5];
  assign ins_o[132] = ver_i[4];
  assign ins_o[131] = ver_i[3];
  assign ins_o[130] = ver_i[2];
  assign ins_o[129] = ver_i[1];
  assign ins_o[128] = ver_i[0];
  assign ins_o[127] = outs_i[319];
  assign ins_o[126] = outs_i[318];
  assign ins_o[125] = outs_i[317];
  assign ins_o[124] = outs_i[316];
  assign ins_o[123] = outs_i[315];
  assign ins_o[122] = outs_i[314];
  assign ins_o[121] = outs_i[313];
  assign ins_o[120] = outs_i[312];
  assign ins_o[119] = outs_i[311];
  assign ins_o[118] = outs_i[310];
  assign ins_o[117] = outs_i[309];
  assign ins_o[116] = outs_i[308];
  assign ins_o[115] = outs_i[307];
  assign ins_o[114] = outs_i[306];
  assign ins_o[113] = outs_i[305];
  assign ins_o[112] = outs_i[304];
  assign ins_o[111] = outs_i[303];
  assign ins_o[110] = outs_i[302];
  assign ins_o[109] = outs_i[301];
  assign ins_o[108] = outs_i[300];
  assign ins_o[107] = outs_i[299];
  assign ins_o[106] = outs_i[298];
  assign ins_o[105] = outs_i[297];
  assign ins_o[104] = outs_i[296];
  assign ins_o[103] = outs_i[295];
  assign ins_o[102] = outs_i[294];
  assign ins_o[101] = outs_i[293];
  assign ins_o[100] = outs_i[292];
  assign ins_o[99] = outs_i[291];
  assign ins_o[98] = outs_i[290];
  assign ins_o[97] = outs_i[289];
  assign ins_o[96] = outs_i[288];
  assign ins_o[95] = outs_i[287];
  assign ins_o[94] = outs_i[286];
  assign ins_o[93] = outs_i[285];
  assign ins_o[92] = outs_i[284];
  assign ins_o[91] = outs_i[283];
  assign ins_o[90] = outs_i[282];
  assign ins_o[89] = outs_i[281];
  assign ins_o[88] = outs_i[280];
  assign ins_o[87] = outs_i[279];
  assign ins_o[86] = outs_i[278];
  assign ins_o[85] = outs_i[277];
  assign ins_o[84] = outs_i[276];
  assign ins_o[83] = outs_i[275];
  assign ins_o[82] = outs_i[274];
  assign ins_o[81] = outs_i[273];
  assign ins_o[80] = outs_i[272];
  assign ins_o[79] = outs_i[271];
  assign ins_o[78] = outs_i[270];
  assign ins_o[77] = outs_i[269];
  assign ins_o[76] = outs_i[268];
  assign ins_o[75] = outs_i[267];
  assign ins_o[74] = outs_i[266];
  assign ins_o[73] = outs_i[265];
  assign ins_o[72] = outs_i[264];
  assign ins_o[71] = outs_i[263];
  assign ins_o[70] = outs_i[262];
  assign ins_o[69] = outs_i[261];
  assign ins_o[68] = outs_i[260];
  assign ins_o[67] = outs_i[259];
  assign ins_o[66] = outs_i[258];
  assign ins_o[65] = outs_i[257];
  assign ins_o[64] = outs_i[256];
  assign ins_o[63] = hor_i[63];
  assign ins_o[62] = hor_i[62];
  assign ins_o[61] = hor_i[61];
  assign ins_o[60] = hor_i[60];
  assign ins_o[59] = hor_i[59];
  assign ins_o[58] = hor_i[58];
  assign ins_o[57] = hor_i[57];
  assign ins_o[56] = hor_i[56];
  assign ins_o[55] = hor_i[55];
  assign ins_o[54] = hor_i[54];
  assign ins_o[53] = hor_i[53];
  assign ins_o[52] = hor_i[52];
  assign ins_o[51] = hor_i[51];
  assign ins_o[50] = hor_i[50];
  assign ins_o[49] = hor_i[49];
  assign ins_o[48] = hor_i[48];
  assign ins_o[47] = hor_i[47];
  assign ins_o[46] = hor_i[46];
  assign ins_o[45] = hor_i[45];
  assign ins_o[44] = hor_i[44];
  assign ins_o[43] = hor_i[43];
  assign ins_o[42] = hor_i[42];
  assign ins_o[41] = hor_i[41];
  assign ins_o[40] = hor_i[40];
  assign ins_o[39] = hor_i[39];
  assign ins_o[38] = hor_i[38];
  assign ins_o[37] = hor_i[37];
  assign ins_o[36] = hor_i[36];
  assign ins_o[35] = hor_i[35];
  assign ins_o[34] = hor_i[34];
  assign ins_o[33] = hor_i[33];
  assign ins_o[32] = hor_i[32];
  assign ins_o[31] = hor_i[31];
  assign ins_o[30] = hor_i[30];
  assign ins_o[29] = hor_i[29];
  assign ins_o[28] = hor_i[28];
  assign ins_o[27] = hor_i[27];
  assign ins_o[26] = hor_i[26];
  assign ins_o[25] = hor_i[25];
  assign ins_o[24] = hor_i[24];
  assign ins_o[23] = hor_i[23];
  assign ins_o[22] = hor_i[22];
  assign ins_o[21] = hor_i[21];
  assign ins_o[20] = hor_i[20];
  assign ins_o[19] = hor_i[19];
  assign ins_o[18] = hor_i[18];
  assign ins_o[17] = hor_i[17];
  assign ins_o[16] = hor_i[16];
  assign ins_o[15] = hor_i[15];
  assign ins_o[14] = hor_i[14];
  assign ins_o[13] = hor_i[13];
  assign ins_o[12] = hor_i[12];
  assign ins_o[11] = hor_i[11];
  assign ins_o[10] = hor_i[10];
  assign ins_o[9] = hor_i[9];
  assign ins_o[8] = hor_i[8];
  assign ins_o[7] = hor_i[7];
  assign ins_o[6] = hor_i[6];
  assign ins_o[5] = hor_i[5];
  assign ins_o[4] = hor_i[4];
  assign ins_o[3] = hor_i[3];
  assign ins_o[2] = hor_i[2];
  assign ins_o[1] = hor_i[1];
  assign ins_o[0] = hor_i[0];
  assign hor_o[127] = outs_i[383];
  assign hor_o[126] = outs_i[382];
  assign hor_o[125] = outs_i[381];
  assign hor_o[124] = outs_i[380];
  assign hor_o[123] = outs_i[379];
  assign hor_o[122] = outs_i[378];
  assign hor_o[121] = outs_i[377];
  assign hor_o[120] = outs_i[376];
  assign hor_o[119] = outs_i[375];
  assign hor_o[118] = outs_i[374];
  assign hor_o[117] = outs_i[373];
  assign hor_o[116] = outs_i[372];
  assign hor_o[115] = outs_i[371];
  assign hor_o[114] = outs_i[370];
  assign hor_o[113] = outs_i[369];
  assign hor_o[112] = outs_i[368];
  assign hor_o[111] = outs_i[367];
  assign hor_o[110] = outs_i[366];
  assign hor_o[109] = outs_i[365];
  assign hor_o[108] = outs_i[364];
  assign hor_o[107] = outs_i[363];
  assign hor_o[106] = outs_i[362];
  assign hor_o[105] = outs_i[361];
  assign hor_o[104] = outs_i[360];
  assign hor_o[103] = outs_i[359];
  assign hor_o[102] = outs_i[358];
  assign hor_o[101] = outs_i[357];
  assign hor_o[100] = outs_i[356];
  assign hor_o[99] = outs_i[355];
  assign hor_o[98] = outs_i[354];
  assign hor_o[97] = outs_i[353];
  assign hor_o[96] = outs_i[352];
  assign hor_o[95] = outs_i[351];
  assign hor_o[94] = outs_i[350];
  assign hor_o[93] = outs_i[349];
  assign hor_o[92] = outs_i[348];
  assign hor_o[91] = outs_i[347];
  assign hor_o[90] = outs_i[346];
  assign hor_o[89] = outs_i[345];
  assign hor_o[88] = outs_i[344];
  assign hor_o[87] = outs_i[343];
  assign hor_o[86] = outs_i[342];
  assign hor_o[85] = outs_i[341];
  assign hor_o[84] = outs_i[340];
  assign hor_o[83] = outs_i[339];
  assign hor_o[82] = outs_i[338];
  assign hor_o[81] = outs_i[337];
  assign hor_o[80] = outs_i[336];
  assign hor_o[79] = outs_i[335];
  assign hor_o[78] = outs_i[334];
  assign hor_o[77] = outs_i[333];
  assign hor_o[76] = outs_i[332];
  assign hor_o[75] = outs_i[331];
  assign hor_o[74] = outs_i[330];
  assign hor_o[73] = outs_i[329];
  assign hor_o[72] = outs_i[328];
  assign hor_o[71] = outs_i[327];
  assign hor_o[70] = outs_i[326];
  assign hor_o[69] = outs_i[325];
  assign hor_o[68] = outs_i[324];
  assign hor_o[67] = outs_i[323];
  assign hor_o[66] = outs_i[322];
  assign hor_o[65] = outs_i[321];
  assign hor_o[64] = outs_i[320];
  assign hor_o[63] = outs_i[63];
  assign hor_o[62] = outs_i[62];
  assign hor_o[61] = outs_i[61];
  assign hor_o[60] = outs_i[60];
  assign hor_o[59] = outs_i[59];
  assign hor_o[58] = outs_i[58];
  assign hor_o[57] = outs_i[57];
  assign hor_o[56] = outs_i[56];
  assign hor_o[55] = outs_i[55];
  assign hor_o[54] = outs_i[54];
  assign hor_o[53] = outs_i[53];
  assign hor_o[52] = outs_i[52];
  assign hor_o[51] = outs_i[51];
  assign hor_o[50] = outs_i[50];
  assign hor_o[49] = outs_i[49];
  assign hor_o[48] = outs_i[48];
  assign hor_o[47] = outs_i[47];
  assign hor_o[46] = outs_i[46];
  assign hor_o[45] = outs_i[45];
  assign hor_o[44] = outs_i[44];
  assign hor_o[43] = outs_i[43];
  assign hor_o[42] = outs_i[42];
  assign hor_o[41] = outs_i[41];
  assign hor_o[40] = outs_i[40];
  assign hor_o[39] = outs_i[39];
  assign hor_o[38] = outs_i[38];
  assign hor_o[37] = outs_i[37];
  assign hor_o[36] = outs_i[36];
  assign hor_o[35] = outs_i[35];
  assign hor_o[34] = outs_i[34];
  assign hor_o[33] = outs_i[33];
  assign hor_o[32] = outs_i[32];
  assign hor_o[31] = outs_i[31];
  assign hor_o[30] = outs_i[30];
  assign hor_o[29] = outs_i[29];
  assign hor_o[28] = outs_i[28];
  assign hor_o[27] = outs_i[27];
  assign hor_o[26] = outs_i[26];
  assign hor_o[25] = outs_i[25];
  assign hor_o[24] = outs_i[24];
  assign hor_o[23] = outs_i[23];
  assign hor_o[22] = outs_i[22];
  assign hor_o[21] = outs_i[21];
  assign hor_o[20] = outs_i[20];
  assign hor_o[19] = outs_i[19];
  assign hor_o[18] = outs_i[18];
  assign hor_o[17] = outs_i[17];
  assign hor_o[16] = outs_i[16];
  assign hor_o[15] = outs_i[15];
  assign hor_o[14] = outs_i[14];
  assign hor_o[13] = outs_i[13];
  assign hor_o[12] = outs_i[12];
  assign hor_o[11] = outs_i[11];
  assign hor_o[10] = outs_i[10];
  assign hor_o[9] = outs_i[9];
  assign hor_o[8] = outs_i[8];
  assign hor_o[7] = outs_i[7];
  assign hor_o[6] = outs_i[6];
  assign hor_o[5] = outs_i[5];
  assign hor_o[4] = outs_i[4];
  assign hor_o[3] = outs_i[3];
  assign hor_o[2] = outs_i[2];
  assign hor_o[1] = outs_i[1];
  assign hor_o[0] = outs_i[0];
  assign ver_o[255] = outs_i[511];
  assign ver_o[254] = outs_i[510];
  assign ver_o[253] = outs_i[509];
  assign ver_o[252] = outs_i[508];
  assign ver_o[251] = outs_i[507];
  assign ver_o[250] = outs_i[506];
  assign ver_o[249] = outs_i[505];
  assign ver_o[248] = outs_i[504];
  assign ver_o[247] = outs_i[503];
  assign ver_o[246] = outs_i[502];
  assign ver_o[245] = outs_i[501];
  assign ver_o[244] = outs_i[500];
  assign ver_o[243] = outs_i[499];
  assign ver_o[242] = outs_i[498];
  assign ver_o[241] = outs_i[497];
  assign ver_o[240] = outs_i[496];
  assign ver_o[239] = outs_i[495];
  assign ver_o[238] = outs_i[494];
  assign ver_o[237] = outs_i[493];
  assign ver_o[236] = outs_i[492];
  assign ver_o[235] = outs_i[491];
  assign ver_o[234] = outs_i[490];
  assign ver_o[233] = outs_i[489];
  assign ver_o[232] = outs_i[488];
  assign ver_o[231] = outs_i[487];
  assign ver_o[230] = outs_i[486];
  assign ver_o[229] = outs_i[485];
  assign ver_o[228] = outs_i[484];
  assign ver_o[227] = outs_i[483];
  assign ver_o[226] = outs_i[482];
  assign ver_o[225] = outs_i[481];
  assign ver_o[224] = outs_i[480];
  assign ver_o[223] = outs_i[479];
  assign ver_o[222] = outs_i[478];
  assign ver_o[221] = outs_i[477];
  assign ver_o[220] = outs_i[476];
  assign ver_o[219] = outs_i[475];
  assign ver_o[218] = outs_i[474];
  assign ver_o[217] = outs_i[473];
  assign ver_o[216] = outs_i[472];
  assign ver_o[215] = outs_i[471];
  assign ver_o[214] = outs_i[470];
  assign ver_o[213] = outs_i[469];
  assign ver_o[212] = outs_i[468];
  assign ver_o[211] = outs_i[467];
  assign ver_o[210] = outs_i[466];
  assign ver_o[209] = outs_i[465];
  assign ver_o[208] = outs_i[464];
  assign ver_o[207] = outs_i[463];
  assign ver_o[206] = outs_i[462];
  assign ver_o[205] = outs_i[461];
  assign ver_o[204] = outs_i[460];
  assign ver_o[203] = outs_i[459];
  assign ver_o[202] = outs_i[458];
  assign ver_o[201] = outs_i[457];
  assign ver_o[200] = outs_i[456];
  assign ver_o[199] = outs_i[455];
  assign ver_o[198] = outs_i[454];
  assign ver_o[197] = outs_i[453];
  assign ver_o[196] = outs_i[452];
  assign ver_o[195] = outs_i[451];
  assign ver_o[194] = outs_i[450];
  assign ver_o[193] = outs_i[449];
  assign ver_o[192] = outs_i[448];
  assign ver_o[191] = outs_i[255];
  assign ver_o[190] = outs_i[254];
  assign ver_o[189] = outs_i[253];
  assign ver_o[188] = outs_i[252];
  assign ver_o[187] = outs_i[251];
  assign ver_o[186] = outs_i[250];
  assign ver_o[185] = outs_i[249];
  assign ver_o[184] = outs_i[248];
  assign ver_o[183] = outs_i[247];
  assign ver_o[182] = outs_i[246];
  assign ver_o[181] = outs_i[245];
  assign ver_o[180] = outs_i[244];
  assign ver_o[179] = outs_i[243];
  assign ver_o[178] = outs_i[242];
  assign ver_o[177] = outs_i[241];
  assign ver_o[176] = outs_i[240];
  assign ver_o[175] = outs_i[239];
  assign ver_o[174] = outs_i[238];
  assign ver_o[173] = outs_i[237];
  assign ver_o[172] = outs_i[236];
  assign ver_o[171] = outs_i[235];
  assign ver_o[170] = outs_i[234];
  assign ver_o[169] = outs_i[233];
  assign ver_o[168] = outs_i[232];
  assign ver_o[167] = outs_i[231];
  assign ver_o[166] = outs_i[230];
  assign ver_o[165] = outs_i[229];
  assign ver_o[164] = outs_i[228];
  assign ver_o[163] = outs_i[227];
  assign ver_o[162] = outs_i[226];
  assign ver_o[161] = outs_i[225];
  assign ver_o[160] = outs_i[224];
  assign ver_o[159] = outs_i[223];
  assign ver_o[158] = outs_i[222];
  assign ver_o[157] = outs_i[221];
  assign ver_o[156] = outs_i[220];
  assign ver_o[155] = outs_i[219];
  assign ver_o[154] = outs_i[218];
  assign ver_o[153] = outs_i[217];
  assign ver_o[152] = outs_i[216];
  assign ver_o[151] = outs_i[215];
  assign ver_o[150] = outs_i[214];
  assign ver_o[149] = outs_i[213];
  assign ver_o[148] = outs_i[212];
  assign ver_o[147] = outs_i[211];
  assign ver_o[146] = outs_i[210];
  assign ver_o[145] = outs_i[209];
  assign ver_o[144] = outs_i[208];
  assign ver_o[143] = outs_i[207];
  assign ver_o[142] = outs_i[206];
  assign ver_o[141] = outs_i[205];
  assign ver_o[140] = outs_i[204];
  assign ver_o[139] = outs_i[203];
  assign ver_o[138] = outs_i[202];
  assign ver_o[137] = outs_i[201];
  assign ver_o[136] = outs_i[200];
  assign ver_o[135] = outs_i[199];
  assign ver_o[134] = outs_i[198];
  assign ver_o[133] = outs_i[197];
  assign ver_o[132] = outs_i[196];
  assign ver_o[131] = outs_i[195];
  assign ver_o[130] = outs_i[194];
  assign ver_o[129] = outs_i[193];
  assign ver_o[128] = outs_i[192];
  assign ver_o[127] = outs_i[447];
  assign ver_o[126] = outs_i[446];
  assign ver_o[125] = outs_i[445];
  assign ver_o[124] = outs_i[444];
  assign ver_o[123] = outs_i[443];
  assign ver_o[122] = outs_i[442];
  assign ver_o[121] = outs_i[441];
  assign ver_o[120] = outs_i[440];
  assign ver_o[119] = outs_i[439];
  assign ver_o[118] = outs_i[438];
  assign ver_o[117] = outs_i[437];
  assign ver_o[116] = outs_i[436];
  assign ver_o[115] = outs_i[435];
  assign ver_o[114] = outs_i[434];
  assign ver_o[113] = outs_i[433];
  assign ver_o[112] = outs_i[432];
  assign ver_o[111] = outs_i[431];
  assign ver_o[110] = outs_i[430];
  assign ver_o[109] = outs_i[429];
  assign ver_o[108] = outs_i[428];
  assign ver_o[107] = outs_i[427];
  assign ver_o[106] = outs_i[426];
  assign ver_o[105] = outs_i[425];
  assign ver_o[104] = outs_i[424];
  assign ver_o[103] = outs_i[423];
  assign ver_o[102] = outs_i[422];
  assign ver_o[101] = outs_i[421];
  assign ver_o[100] = outs_i[420];
  assign ver_o[99] = outs_i[419];
  assign ver_o[98] = outs_i[418];
  assign ver_o[97] = outs_i[417];
  assign ver_o[96] = outs_i[416];
  assign ver_o[95] = outs_i[415];
  assign ver_o[94] = outs_i[414];
  assign ver_o[93] = outs_i[413];
  assign ver_o[92] = outs_i[412];
  assign ver_o[91] = outs_i[411];
  assign ver_o[90] = outs_i[410];
  assign ver_o[89] = outs_i[409];
  assign ver_o[88] = outs_i[408];
  assign ver_o[87] = outs_i[407];
  assign ver_o[86] = outs_i[406];
  assign ver_o[85] = outs_i[405];
  assign ver_o[84] = outs_i[404];
  assign ver_o[83] = outs_i[403];
  assign ver_o[82] = outs_i[402];
  assign ver_o[81] = outs_i[401];
  assign ver_o[80] = outs_i[400];
  assign ver_o[79] = outs_i[399];
  assign ver_o[78] = outs_i[398];
  assign ver_o[77] = outs_i[397];
  assign ver_o[76] = outs_i[396];
  assign ver_o[75] = outs_i[395];
  assign ver_o[74] = outs_i[394];
  assign ver_o[73] = outs_i[393];
  assign ver_o[72] = outs_i[392];
  assign ver_o[71] = outs_i[391];
  assign ver_o[70] = outs_i[390];
  assign ver_o[69] = outs_i[389];
  assign ver_o[68] = outs_i[388];
  assign ver_o[67] = outs_i[387];
  assign ver_o[66] = outs_i[386];
  assign ver_o[65] = outs_i[385];
  assign ver_o[64] = outs_i[384];
  assign ver_o[63] = outs_i[191];
  assign ver_o[62] = outs_i[190];
  assign ver_o[61] = outs_i[189];
  assign ver_o[60] = outs_i[188];
  assign ver_o[59] = outs_i[187];
  assign ver_o[58] = outs_i[186];
  assign ver_o[57] = outs_i[185];
  assign ver_o[56] = outs_i[184];
  assign ver_o[55] = outs_i[183];
  assign ver_o[54] = outs_i[182];
  assign ver_o[53] = outs_i[181];
  assign ver_o[52] = outs_i[180];
  assign ver_o[51] = outs_i[179];
  assign ver_o[50] = outs_i[178];
  assign ver_o[49] = outs_i[177];
  assign ver_o[48] = outs_i[176];
  assign ver_o[47] = outs_i[175];
  assign ver_o[46] = outs_i[174];
  assign ver_o[45] = outs_i[173];
  assign ver_o[44] = outs_i[172];
  assign ver_o[43] = outs_i[171];
  assign ver_o[42] = outs_i[170];
  assign ver_o[41] = outs_i[169];
  assign ver_o[40] = outs_i[168];
  assign ver_o[39] = outs_i[167];
  assign ver_o[38] = outs_i[166];
  assign ver_o[37] = outs_i[165];
  assign ver_o[36] = outs_i[164];
  assign ver_o[35] = outs_i[163];
  assign ver_o[34] = outs_i[162];
  assign ver_o[33] = outs_i[161];
  assign ver_o[32] = outs_i[160];
  assign ver_o[31] = outs_i[159];
  assign ver_o[30] = outs_i[158];
  assign ver_o[29] = outs_i[157];
  assign ver_o[28] = outs_i[156];
  assign ver_o[27] = outs_i[155];
  assign ver_o[26] = outs_i[154];
  assign ver_o[25] = outs_i[153];
  assign ver_o[24] = outs_i[152];
  assign ver_o[23] = outs_i[151];
  assign ver_o[22] = outs_i[150];
  assign ver_o[21] = outs_i[149];
  assign ver_o[20] = outs_i[148];
  assign ver_o[19] = outs_i[147];
  assign ver_o[18] = outs_i[146];
  assign ver_o[17] = outs_i[145];
  assign ver_o[16] = outs_i[144];
  assign ver_o[15] = outs_i[143];
  assign ver_o[14] = outs_i[142];
  assign ver_o[13] = outs_i[141];
  assign ver_o[12] = outs_i[140];
  assign ver_o[11] = outs_i[139];
  assign ver_o[10] = outs_i[138];
  assign ver_o[9] = outs_i[137];
  assign ver_o[8] = outs_i[136];
  assign ver_o[7] = outs_i[135];
  assign ver_o[6] = outs_i[134];
  assign ver_o[5] = outs_i[133];
  assign ver_o[4] = outs_i[132];
  assign ver_o[3] = outs_i[131];
  assign ver_o[2] = outs_i[130];
  assign ver_o[1] = outs_i[129];
  assign ver_o[0] = outs_i[128];

endmodule