module ptw_s00000001
(
  clk_i,
  rst_ni,
  flush_i,
  ptw_active_o,
  walking_instr_o,
  ptw_error_o,
  enable_translation_i,
  en_ld_st_translation_i,
  lsu_is_store_i,
  req_port_i,
  req_port_o,
  itlb_update_o,
  dtlb_update_o,
  update_vaddr_o,
  asid_i,
  itlb_access_i,
  itlb_hit_i,
  itlb_vaddr_i,
  dtlb_access_i,
  dtlb_hit_i,
  dtlb_vaddr_i,
  satp_ppn_i,
  mxr_i,
  itlb_miss_o,
  dtlb_miss_o
);

  input [65:0] req_port_i;
  output [133:0] req_port_o;
  output [94:0] itlb_update_o;
  output [94:0] dtlb_update_o;
  output [38:0] update_vaddr_o;
  input [0:0] asid_i;
  input [63:0] itlb_vaddr_i;
  input [63:0] dtlb_vaddr_i;
  input [43:0] satp_ppn_i;
  input clk_i;
  input rst_ni;
  input flush_i;
  input enable_translation_i;
  input en_ld_st_translation_i;
  input lsu_is_store_i;
  input itlb_access_i;
  input itlb_hit_i;
  input dtlb_access_i;
  input dtlb_hit_i;
  input mxr_i;
  output ptw_active_o;
  output walking_instr_o;
  output ptw_error_o;
  output itlb_miss_o;
  output dtlb_miss_o;
  wire [94:0] dtlb_update_o;
  wire ptw_active_o,ptw_error_o,itlb_miss_o,dtlb_miss_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,tag_valid_n,
  global_mapping_n,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,
  N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,
  N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,
  N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N320,N321,N323,N325,N327,N329,N330,
  N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,
  N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,
  N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390;
  wire [1:0] ptw_lvl_n;
  wire [55:0] ptw_pptr_n;
  wire [2:0] state_d;
  reg data_rvalid_q,walking_instr_o,global_mapping_q,pte_g_;
  reg [2:0] state_q;
  reg [1:0] ptw_lvl_q;
  reg [133:0] req_port_o;
  reg [94:0] itlb_update_o;
  reg [38:0] update_vaddr_o;
  assign req_port_o[2] = 1'b1;
  assign req_port_o[3] = 1'b1;
  assign req_port_o[4] = 1'b1;
  assign req_port_o[5] = 1'b1;
  assign req_port_o[6] = 1'b1;
  assign req_port_o[7] = 1'b1;
  assign req_port_o[8] = 1'b1;
  assign req_port_o[9] = 1'b1;
  assign req_port_o[10] = 1'b1;
  assign req_port_o[11] = 1'b1;
  assign req_port_o[12] = 1'b0;
  assign req_port_o[14] = 1'b0;
  assign req_port_o[15] = 1'b0;
  assign req_port_o[16] = 1'b0;
  assign req_port_o[17] = 1'b0;
  assign req_port_o[18] = 1'b0;
  assign req_port_o[19] = 1'b0;
  assign req_port_o[20] = 1'b0;
  assign req_port_o[21] = 1'b0;
  assign req_port_o[22] = 1'b0;
  assign req_port_o[23] = 1'b0;
  assign req_port_o[24] = 1'b0;
  assign req_port_o[25] = 1'b0;
  assign req_port_o[26] = 1'b0;
  assign req_port_o[27] = 1'b0;
  assign req_port_o[28] = 1'b0;
  assign req_port_o[29] = 1'b0;
  assign req_port_o[30] = 1'b0;
  assign req_port_o[31] = 1'b0;
  assign req_port_o[32] = 1'b0;
  assign req_port_o[33] = 1'b0;
  assign req_port_o[34] = 1'b0;
  assign req_port_o[35] = 1'b0;
  assign req_port_o[36] = 1'b0;
  assign req_port_o[37] = 1'b0;
  assign req_port_o[38] = 1'b0;
  assign req_port_o[39] = 1'b0;
  assign req_port_o[40] = 1'b0;
  assign req_port_o[41] = 1'b0;
  assign req_port_o[42] = 1'b0;
  assign req_port_o[43] = 1'b0;
  assign req_port_o[44] = 1'b0;
  assign req_port_o[45] = 1'b0;
  assign req_port_o[46] = 1'b0;
  assign req_port_o[47] = 1'b0;
  assign req_port_o[48] = 1'b0;
  assign req_port_o[49] = 1'b0;
  assign req_port_o[50] = 1'b0;
  assign req_port_o[51] = 1'b0;
  assign req_port_o[52] = 1'b0;
  assign req_port_o[53] = 1'b0;
  assign req_port_o[54] = 1'b0;
  assign req_port_o[55] = 1'b0;
  assign req_port_o[56] = 1'b0;
  assign req_port_o[57] = 1'b0;
  assign req_port_o[58] = 1'b0;
  assign req_port_o[59] = 1'b0;
  assign req_port_o[60] = 1'b0;
  assign req_port_o[61] = 1'b0;
  assign req_port_o[62] = 1'b0;
  assign req_port_o[63] = 1'b0;
  assign req_port_o[64] = 1'b0;
  assign req_port_o[65] = 1'b0;
  assign req_port_o[66] = 1'b0;
  assign req_port_o[67] = 1'b0;
  assign req_port_o[68] = 1'b0;
  assign req_port_o[69] = 1'b0;
  assign req_port_o[70] = 1'b0;
  assign req_port_o[71] = 1'b0;
  assign req_port_o[72] = 1'b0;
  assign req_port_o[73] = 1'b0;
  assign req_port_o[74] = 1'b0;
  assign req_port_o[75] = 1'b0;
  assign req_port_o[76] = 1'b0;
  assign req_port_o[77] = 1'b0;
  assign req_port_o[1] = 1'b0;
  assign dtlb_update_o[64] = itlb_update_o[64];
  assign dtlb_update_o[63] = itlb_update_o[63];
  assign dtlb_update_o[62] = itlb_update_o[62];
  assign dtlb_update_o[61] = itlb_update_o[61];
  assign dtlb_update_o[60] = itlb_update_o[60];
  assign dtlb_update_o[59] = itlb_update_o[59];
  assign dtlb_update_o[58] = itlb_update_o[58];
  assign dtlb_update_o[57] = itlb_update_o[57];
  assign dtlb_update_o[56] = itlb_update_o[56];
  assign dtlb_update_o[55] = itlb_update_o[55];
  assign dtlb_update_o[54] = itlb_update_o[54];
  assign dtlb_update_o[53] = itlb_update_o[53];
  assign dtlb_update_o[52] = itlb_update_o[52];
  assign dtlb_update_o[51] = itlb_update_o[51];
  assign dtlb_update_o[50] = itlb_update_o[50];
  assign dtlb_update_o[49] = itlb_update_o[49];
  assign dtlb_update_o[48] = itlb_update_o[48];
  assign dtlb_update_o[47] = itlb_update_o[47];
  assign dtlb_update_o[46] = itlb_update_o[46];
  assign dtlb_update_o[45] = itlb_update_o[45];
  assign dtlb_update_o[44] = itlb_update_o[44];
  assign dtlb_update_o[43] = itlb_update_o[43];
  assign dtlb_update_o[42] = itlb_update_o[42];
  assign dtlb_update_o[41] = itlb_update_o[41];
  assign dtlb_update_o[40] = itlb_update_o[40];
  assign dtlb_update_o[39] = itlb_update_o[39];
  assign dtlb_update_o[38] = itlb_update_o[38];
  assign dtlb_update_o[37] = itlb_update_o[37];
  assign dtlb_update_o[36] = itlb_update_o[36];
  assign dtlb_update_o[35] = itlb_update_o[35];
  assign dtlb_update_o[34] = itlb_update_o[34];
  assign dtlb_update_o[33] = itlb_update_o[33];
  assign dtlb_update_o[32] = itlb_update_o[32];
  assign dtlb_update_o[31] = itlb_update_o[31];
  assign dtlb_update_o[30] = itlb_update_o[30];
  assign dtlb_update_o[29] = itlb_update_o[29];
  assign dtlb_update_o[28] = itlb_update_o[28];
  assign dtlb_update_o[27] = itlb_update_o[27];
  assign dtlb_update_o[26] = itlb_update_o[26];
  assign dtlb_update_o[25] = itlb_update_o[25];
  assign dtlb_update_o[24] = itlb_update_o[24];
  assign dtlb_update_o[23] = itlb_update_o[23];
  assign dtlb_update_o[22] = itlb_update_o[22];
  assign dtlb_update_o[21] = itlb_update_o[21];
  assign dtlb_update_o[20] = itlb_update_o[20];
  assign dtlb_update_o[19] = itlb_update_o[19];
  assign dtlb_update_o[18] = itlb_update_o[18];
  assign dtlb_update_o[17] = itlb_update_o[17];
  assign dtlb_update_o[16] = itlb_update_o[16];
  assign dtlb_update_o[15] = itlb_update_o[15];
  assign dtlb_update_o[14] = itlb_update_o[14];
  assign dtlb_update_o[13] = itlb_update_o[13];
  assign dtlb_update_o[12] = itlb_update_o[12];
  assign dtlb_update_o[11] = itlb_update_o[11];
  assign dtlb_update_o[10] = itlb_update_o[10];
  assign dtlb_update_o[9] = itlb_update_o[9];
  assign dtlb_update_o[8] = itlb_update_o[8];
  assign dtlb_update_o[7] = itlb_update_o[7];
  assign dtlb_update_o[6] = itlb_update_o[6];
  assign dtlb_update_o[4] = itlb_update_o[4];
  assign dtlb_update_o[3] = itlb_update_o[3];
  assign dtlb_update_o[2] = itlb_update_o[2];
  assign dtlb_update_o[1] = itlb_update_o[1];
  assign dtlb_update_o[0] = itlb_update_o[0];
  assign dtlb_update_o[91] = update_vaddr_o[38];
  assign itlb_update_o[91] = update_vaddr_o[38];
  assign dtlb_update_o[90] = update_vaddr_o[37];
  assign itlb_update_o[90] = update_vaddr_o[37];
  assign dtlb_update_o[89] = update_vaddr_o[36];
  assign itlb_update_o[89] = update_vaddr_o[36];
  assign dtlb_update_o[88] = update_vaddr_o[35];
  assign itlb_update_o[88] = update_vaddr_o[35];
  assign dtlb_update_o[87] = update_vaddr_o[34];
  assign itlb_update_o[87] = update_vaddr_o[34];
  assign dtlb_update_o[86] = update_vaddr_o[33];
  assign itlb_update_o[86] = update_vaddr_o[33];
  assign dtlb_update_o[85] = update_vaddr_o[32];
  assign itlb_update_o[85] = update_vaddr_o[32];
  assign dtlb_update_o[84] = update_vaddr_o[31];
  assign itlb_update_o[84] = update_vaddr_o[31];
  assign dtlb_update_o[83] = update_vaddr_o[30];
  assign itlb_update_o[83] = update_vaddr_o[30];
  assign dtlb_update_o[82] = update_vaddr_o[29];
  assign itlb_update_o[82] = update_vaddr_o[29];
  assign dtlb_update_o[81] = update_vaddr_o[28];
  assign itlb_update_o[81] = update_vaddr_o[28];
  assign dtlb_update_o[80] = update_vaddr_o[27];
  assign itlb_update_o[80] = update_vaddr_o[27];
  assign dtlb_update_o[79] = update_vaddr_o[26];
  assign itlb_update_o[79] = update_vaddr_o[26];
  assign dtlb_update_o[78] = update_vaddr_o[25];
  assign itlb_update_o[78] = update_vaddr_o[25];
  assign dtlb_update_o[77] = update_vaddr_o[24];
  assign itlb_update_o[77] = update_vaddr_o[24];
  assign dtlb_update_o[76] = update_vaddr_o[23];
  assign itlb_update_o[76] = update_vaddr_o[23];
  assign dtlb_update_o[75] = update_vaddr_o[22];
  assign itlb_update_o[75] = update_vaddr_o[22];
  assign dtlb_update_o[74] = update_vaddr_o[21];
  assign itlb_update_o[74] = update_vaddr_o[21];
  assign dtlb_update_o[73] = update_vaddr_o[20];
  assign itlb_update_o[73] = update_vaddr_o[20];
  assign dtlb_update_o[72] = update_vaddr_o[19];
  assign itlb_update_o[72] = update_vaddr_o[19];
  assign dtlb_update_o[71] = update_vaddr_o[18];
  assign itlb_update_o[71] = update_vaddr_o[18];
  assign dtlb_update_o[70] = update_vaddr_o[17];
  assign itlb_update_o[70] = update_vaddr_o[17];
  assign dtlb_update_o[69] = update_vaddr_o[16];
  assign itlb_update_o[69] = update_vaddr_o[16];
  assign dtlb_update_o[68] = update_vaddr_o[15];
  assign itlb_update_o[68] = update_vaddr_o[15];
  assign dtlb_update_o[67] = update_vaddr_o[14];
  assign itlb_update_o[67] = update_vaddr_o[14];
  assign dtlb_update_o[66] = update_vaddr_o[13];
  assign itlb_update_o[66] = update_vaddr_o[13];
  assign dtlb_update_o[65] = update_vaddr_o[12];
  assign itlb_update_o[65] = update_vaddr_o[12];
  assign N27 = N26 & N329;
  assign N28 = N27 & N333;
  assign N29 = state_q[2] | state_q[1];
  assign N30 = N29 | N333;
  assign N32 = state_q[2] | N329;
  assign N33 = N32 | state_q[0];
  assign N35 = N26 | state_q[1];
  assign N36 = N35 | state_q[0];
  assign N38 = state_q[2] | N329;
  assign N39 = N38 | N333;
  assign N41 = state_q[2] & state_q[0];
  assign N42 = state_q[2] & state_q[1];

  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      data_rvalid_q <= 1'b0;
    end else if(1'b1) begin
      data_rvalid_q <= req_port_i[64];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      state_q[2] <= 1'b0;
    end else if(N261) begin
      state_q[2] <= state_d[2];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      state_q[1] <= 1'b0;
    end else if(N261) begin
      state_q[1] <= state_d[1];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      state_q[0] <= 1'b0;
    end else if(N261) begin
      state_q[0] <= state_d[0];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      walking_instr_o <= 1'b0;
    end else if(N266) begin
      walking_instr_o <= N88;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      ptw_lvl_q[1] <= 1'b0;
    end else if(N279) begin
      ptw_lvl_q[1] <= ptw_lvl_n[1];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      ptw_lvl_q[0] <= 1'b0;
    end else if(N287) begin
      ptw_lvl_q[0] <= ptw_lvl_n[0];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[0] <= 1'b0;
    end else if(1'b1) begin
      req_port_o[0] <= tag_valid_n;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[64] <= 1'b0;
    end else if(N294) begin
      itlb_update_o[64] <= asid_i[0];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[38] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[38] <= N56;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[37] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[37] <= N55;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[36] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[36] <= N54;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[35] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[35] <= N53;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[34] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[34] <= N52;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[33] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[33] <= N51;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[32] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[32] <= N50;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[31] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[31] <= N49;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[30] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[30] <= N48;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[29] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[29] <= N86;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[28] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[28] <= N85;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[27] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[27] <= N84;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[26] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[26] <= N83;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[25] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[25] <= N82;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[24] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[24] <= N81;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[23] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[23] <= N80;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[22] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[22] <= N79;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[21] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[21] <= N78;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[20] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[20] <= N77;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[19] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[19] <= N76;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[18] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[18] <= N75;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[17] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[17] <= N74;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[16] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[16] <= N73;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[15] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[15] <= N72;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[14] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[14] <= N71;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[13] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[13] <= N70;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[12] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[12] <= N69;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[11] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[11] <= N68;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[10] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[10] <= N67;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[9] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[9] <= N66;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[8] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[8] <= N65;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[7] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[7] <= N64;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[6] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[6] <= N63;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[5] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[5] <= N62;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[4] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[4] <= N61;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[3] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[3] <= N60;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[2] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[2] <= N59;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[1] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[1] <= N58;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      update_vaddr_o[0] <= 1'b0;
    end else if(N294) begin
      update_vaddr_o[0] <= N57;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[121] <= 1'b0;
    end else if(N301) begin
      req_port_o[121] <= ptw_pptr_n[55];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[120] <= 1'b0;
    end else if(N301) begin
      req_port_o[120] <= ptw_pptr_n[54];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[119] <= 1'b0;
    end else if(N301) begin
      req_port_o[119] <= ptw_pptr_n[53];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[118] <= 1'b0;
    end else if(N301) begin
      req_port_o[118] <= ptw_pptr_n[52];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[117] <= 1'b0;
    end else if(N301) begin
      req_port_o[117] <= ptw_pptr_n[51];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[116] <= 1'b0;
    end else if(N301) begin
      req_port_o[116] <= ptw_pptr_n[50];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[115] <= 1'b0;
    end else if(N301) begin
      req_port_o[115] <= ptw_pptr_n[49];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[114] <= 1'b0;
    end else if(N310) begin
      req_port_o[114] <= ptw_pptr_n[48];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[113] <= 1'b0;
    end else if(N310) begin
      req_port_o[113] <= ptw_pptr_n[47];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[112] <= 1'b0;
    end else if(N310) begin
      req_port_o[112] <= ptw_pptr_n[46];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[111] <= 1'b0;
    end else if(N310) begin
      req_port_o[111] <= ptw_pptr_n[45];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[110] <= 1'b0;
    end else if(N310) begin
      req_port_o[110] <= ptw_pptr_n[44];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[109] <= 1'b0;
    end else if(N310) begin
      req_port_o[109] <= ptw_pptr_n[43];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[108] <= 1'b0;
    end else if(N310) begin
      req_port_o[108] <= ptw_pptr_n[42];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[107] <= 1'b0;
    end else if(N310) begin
      req_port_o[107] <= ptw_pptr_n[41];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[106] <= 1'b0;
    end else if(N310) begin
      req_port_o[106] <= ptw_pptr_n[40];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[105] <= 1'b0;
    end else if(N310) begin
      req_port_o[105] <= ptw_pptr_n[39];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[104] <= 1'b0;
    end else if(N310) begin
      req_port_o[104] <= ptw_pptr_n[38];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[103] <= 1'b0;
    end else if(N310) begin
      req_port_o[103] <= ptw_pptr_n[37];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[102] <= 1'b0;
    end else if(N310) begin
      req_port_o[102] <= ptw_pptr_n[36];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[101] <= 1'b0;
    end else if(N310) begin
      req_port_o[101] <= ptw_pptr_n[35];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[100] <= 1'b0;
    end else if(N310) begin
      req_port_o[100] <= ptw_pptr_n[34];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[99] <= 1'b0;
    end else if(N310) begin
      req_port_o[99] <= ptw_pptr_n[33];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[98] <= 1'b0;
    end else if(N310) begin
      req_port_o[98] <= ptw_pptr_n[32];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[97] <= 1'b0;
    end else if(N310) begin
      req_port_o[97] <= ptw_pptr_n[31];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[96] <= 1'b0;
    end else if(N310) begin
      req_port_o[96] <= ptw_pptr_n[30];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[95] <= 1'b0;
    end else if(N310) begin
      req_port_o[95] <= ptw_pptr_n[29];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[94] <= 1'b0;
    end else if(N310) begin
      req_port_o[94] <= ptw_pptr_n[28];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[93] <= 1'b0;
    end else if(N310) begin
      req_port_o[93] <= ptw_pptr_n[27];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[92] <= 1'b0;
    end else if(N310) begin
      req_port_o[92] <= ptw_pptr_n[26];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[91] <= 1'b0;
    end else if(N310) begin
      req_port_o[91] <= ptw_pptr_n[25];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[90] <= 1'b0;
    end else if(N310) begin
      req_port_o[90] <= ptw_pptr_n[24];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[89] <= 1'b0;
    end else if(N310) begin
      req_port_o[89] <= ptw_pptr_n[23];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[88] <= 1'b0;
    end else if(N310) begin
      req_port_o[88] <= ptw_pptr_n[22];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[87] <= 1'b0;
    end else if(N310) begin
      req_port_o[87] <= ptw_pptr_n[21];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[86] <= 1'b0;
    end else if(N310) begin
      req_port_o[86] <= ptw_pptr_n[20];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[85] <= 1'b0;
    end else if(N310) begin
      req_port_o[85] <= ptw_pptr_n[19];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[84] <= 1'b0;
    end else if(N310) begin
      req_port_o[84] <= ptw_pptr_n[18];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[83] <= 1'b0;
    end else if(N310) begin
      req_port_o[83] <= ptw_pptr_n[17];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[82] <= 1'b0;
    end else if(N310) begin
      req_port_o[82] <= ptw_pptr_n[16];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[81] <= 1'b0;
    end else if(N310) begin
      req_port_o[81] <= ptw_pptr_n[15];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[80] <= 1'b0;
    end else if(N310) begin
      req_port_o[80] <= ptw_pptr_n[14];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[79] <= 1'b0;
    end else if(N310) begin
      req_port_o[79] <= ptw_pptr_n[13];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[78] <= 1'b0;
    end else if(N310) begin
      req_port_o[78] <= ptw_pptr_n[12];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[133] <= 1'b0;
    end else if(N310) begin
      req_port_o[133] <= ptw_pptr_n[11];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[132] <= 1'b0;
    end else if(N310) begin
      req_port_o[132] <= ptw_pptr_n[10];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[131] <= 1'b0;
    end else if(N310) begin
      req_port_o[131] <= ptw_pptr_n[9];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[130] <= 1'b0;
    end else if(N310) begin
      req_port_o[130] <= ptw_pptr_n[8];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[129] <= 1'b0;
    end else if(N310) begin
      req_port_o[129] <= ptw_pptr_n[7];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[128] <= 1'b0;
    end else if(N310) begin
      req_port_o[128] <= ptw_pptr_n[6];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[127] <= 1'b0;
    end else if(N310) begin
      req_port_o[127] <= ptw_pptr_n[5];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[126] <= 1'b0;
    end else if(N310) begin
      req_port_o[126] <= ptw_pptr_n[4];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[125] <= 1'b0;
    end else if(N310) begin
      req_port_o[125] <= ptw_pptr_n[3];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[124] <= 1'b0;
    end else if(N310) begin
      req_port_o[124] <= ptw_pptr_n[2];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[123] <= 1'b0;
    end else if(N310) begin
      req_port_o[123] <= ptw_pptr_n[1];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      req_port_o[122] <= 1'b0;
    end else if(N310) begin
      req_port_o[122] <= ptw_pptr_n[0];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      global_mapping_q <= 1'b0;
    end else if(N317) begin
      global_mapping_q <= global_mapping_n;
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[63] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[63] <= req_port_i[63];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[62] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[62] <= req_port_i[62];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[61] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[61] <= req_port_i[61];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[60] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[60] <= req_port_i[60];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[59] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[59] <= req_port_i[59];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[58] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[58] <= req_port_i[58];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[57] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[57] <= req_port_i[57];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[56] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[56] <= req_port_i[56];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[55] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[55] <= req_port_i[55];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[54] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[54] <= req_port_i[54];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[53] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[53] <= req_port_i[53];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[52] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[52] <= req_port_i[52];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[51] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[51] <= req_port_i[51];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[50] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[50] <= req_port_i[50];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[49] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[49] <= req_port_i[49];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[48] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[48] <= req_port_i[48];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[47] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[47] <= req_port_i[47];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[46] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[46] <= req_port_i[46];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[45] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[45] <= req_port_i[45];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[44] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[44] <= req_port_i[44];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[43] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[43] <= req_port_i[43];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[42] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[42] <= req_port_i[42];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[41] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[41] <= req_port_i[41];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[40] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[40] <= req_port_i[40];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[39] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[39] <= req_port_i[39];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[38] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[38] <= req_port_i[38];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[37] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[37] <= req_port_i[37];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[36] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[36] <= req_port_i[36];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[35] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[35] <= req_port_i[35];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[34] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[34] <= req_port_i[34];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[33] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[33] <= req_port_i[33];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[32] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[32] <= req_port_i[32];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[31] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[31] <= req_port_i[31];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[30] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[30] <= req_port_i[30];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[29] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[29] <= req_port_i[29];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[28] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[28] <= req_port_i[28];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[27] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[27] <= req_port_i[27];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[26] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[26] <= req_port_i[26];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[25] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[25] <= req_port_i[25];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[24] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[24] <= req_port_i[24];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[23] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[23] <= req_port_i[23];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[22] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[22] <= req_port_i[22];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[21] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[21] <= req_port_i[21];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[20] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[20] <= req_port_i[20];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[19] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[19] <= req_port_i[19];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[18] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[18] <= req_port_i[18];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[17] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[17] <= req_port_i[17];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[16] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[16] <= req_port_i[16];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[15] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[15] <= req_port_i[15];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[14] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[14] <= req_port_i[14];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[13] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[13] <= req_port_i[13];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[12] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[12] <= req_port_i[12];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[11] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[11] <= req_port_i[11];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[10] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[10] <= req_port_i[10];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[9] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[9] <= req_port_i[9];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[8] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[8] <= req_port_i[8];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[7] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[7] <= req_port_i[7];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[6] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[6] <= req_port_i[6];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      pte_g_ <= 1'b0;
    end else if(1'b1) begin
      pte_g_ <= req_port_i[5];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[4] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[4] <= req_port_i[4];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[3] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[3] <= req_port_i[3];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[2] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[2] <= req_port_i[2];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[1] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[1] <= req_port_i[1];
    end 
  end


  always @(posedge clk_i or posedge N249) begin
    if(N249) begin
      itlb_update_o[0] <= 1'b0;
    end else if(1'b1) begin
      itlb_update_o[0] <= req_port_i[0];
    end 
  end

  assign N318 = state_q[1] | state_q[2];
  assign ptw_active_o = state_q[0] | N318;
  assign N320 = ~ptw_lvl_q[0];
  assign N321 = N320 | ptw_lvl_q[1];
  assign itlb_update_o[93] = ~N321;
  assign N323 = ptw_lvl_q[0] | ptw_lvl_q[1];
  assign itlb_update_o[92] = ~N323;
  assign N325 = N320 | ptw_lvl_q[1];
  assign dtlb_update_o[93] = ~N325;
  assign N327 = ptw_lvl_q[0] | ptw_lvl_q[1];
  assign dtlb_update_o[92] = ~N327;
  assign N329 = ~state_q[1];
  assign N330 = N329 | state_q[2];
  assign N331 = state_q[0] | N330;
  assign N332 = ~N331;
  assign N333 = ~state_q[0];
  assign N334 = state_q[1] | state_q[2];
  assign N335 = N333 | N334;
  assign N336 = ~N335;
  assign N337 = ~ptw_lvl_q[1];
  assign N338 = ptw_lvl_q[0] | N337;
  assign N339 = ~N338;
  assign N340 = N320 | ptw_lvl_q[1];
  assign N341 = ~N340;
  assign N342 = ptw_lvl_q[0] | ptw_lvl_q[1];
  assign N343 = ~N342;
  assign N344 = N320 | ptw_lvl_q[1];
  assign N345 = ~N344;
  assign N346 = itlb_update_o[17] | itlb_update_o[18];
  assign N347 = itlb_update_o[16] | N346;
  assign N348 = itlb_update_o[15] | N347;
  assign N349 = itlb_update_o[14] | N348;
  assign N350 = itlb_update_o[13] | N349;
  assign N351 = itlb_update_o[12] | N350;
  assign N352 = itlb_update_o[11] | N351;
  assign N353 = itlb_update_o[10] | N352;
  assign N354 = ptw_lvl_q[0] | ptw_lvl_q[1];
  assign N355 = ~N354;
  assign N356 = itlb_update_o[26] | itlb_update_o[27];
  assign N357 = itlb_update_o[25] | N356;
  assign N358 = itlb_update_o[24] | N357;
  assign N359 = itlb_update_o[23] | N358;
  assign N360 = itlb_update_o[22] | N359;
  assign N361 = itlb_update_o[21] | N360;
  assign N362 = itlb_update_o[20] | N361;
  assign N363 = itlb_update_o[19] | N362;
  assign N364 = itlb_update_o[18] | N363;
  assign N365 = itlb_update_o[17] | N364;
  assign N366 = itlb_update_o[16] | N365;
  assign N367 = itlb_update_o[15] | N366;
  assign N368 = itlb_update_o[14] | N367;
  assign N369 = itlb_update_o[13] | N368;
  assign N370 = itlb_update_o[12] | N369;
  assign N371 = itlb_update_o[11] | N370;
  assign N372 = itlb_update_o[10] | N371;
  assign { N56, N55, N54, N53, N52, N51, N50, N49, N48 } = (N0)? itlb_vaddr_i[38:30] : 
                                                           (N1)? dtlb_vaddr_i[38:30] : 1'b0;
  assign N0 = N44;
  assign N1 = N45;
  assign { N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57 } = (N0)? itlb_vaddr_i[29:0] : 
                                                                                                                                                                    (N1)? dtlb_vaddr_i[29:0] : 1'b0;
  assign N88 = (N0)? 1'b1 : 
               (N87)? 1'b0 : 
               (N2)? 1'b0 : 1'b0;
  assign N2 = 1'b0;
  assign N89 = (N0)? 1'b0 : 
               (N1)? 1'b1 : 
               (N47)? 1'b0 : 1'b0;
  assign N99 = ~N98;
  assign N101 = ~N100;
  assign N104 = (N3)? 1'b0 : 
                (N103)? N100 : 1'b0;
  assign N3 = N102;
  assign N105 = (N3)? 1'b1 : 
                (N103)? N101 : 1'b0;
  assign N106 = (N4)? N99 : 
                (N5)? 1'b0 : 1'b0;
  assign N4 = walking_instr_o;
  assign N5 = N97;
  assign N107 = (N4)? N98 : 
                (N5)? N105 : 1'b0;
  assign N108 = (N4)? 1'b0 : 
                (N5)? N104 : 1'b0;
  assign N113 = (N6)? 1'b1 : 
                (N7)? 1'b1 : 
                (N112)? N107 : 1'b0;
  assign N6 = N109;
  assign N7 = N110;
  assign N114 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N112)? N108 : 1'b0;
  assign N115 = (N6)? 1'b0 : 
                (N7)? 1'b0 : 
                (N112)? N106 : 1'b0;
  assign { N117, N116 } = (N8)? { 1'b0, 1'b1 } : 
                          (N9)? ptw_lvl_q : 1'b0;
  assign N8 = N343;
  assign N9 = N342;
  assign { N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118 } = (N8)? { itlb_update_o[53:10], update_vaddr_o[29:21], 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                              (N9)? { req_port_o[121:78], req_port_o[133:122] } : 1'b0;
  assign { N175, N174 } = (N10)? { 1'b1, 1'b0 } : 
                          (N11)? { N117, N116 } : 1'b0;
  assign N10 = N341;
  assign N11 = N340;
  assign { N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176 } = (N10)? { itlb_update_o[53:10], update_vaddr_o[20:12], 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                              (N11)? { N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118 } : 1'b0;
  assign { N233, N232 } = (N12)? { 1'b1, 1'b0 } : 
                          (N13)? { N175, N174 } : 1'b0;
  assign N12 = N339;
  assign N13 = N338;
  assign N234 = (N14)? N114 : 
                (N96)? 1'b0 : 1'b0;
  assign N14 = N95;
  assign N235 = (N14)? N115 : 
                (N96)? 1'b0 : 1'b0;
  assign { N237, N236 } = (N14)? { N113, 1'b0 } : 
                          (N96)? { N339, N338 } : 1'b0;
  assign { N239, N238 } = (N15)? { 1'b1, 1'b0 } : 
                          (N94)? { N237, N236 } : 1'b0;
  assign N15 = N93;
  assign N240 = (N15)? 1'b0 : 
                (N94)? N234 : 1'b0;
  assign N241 = (N15)? 1'b0 : 
                (N94)? N235 : 1'b0;
  assign N242 = (N16)? N240 : 
                (N17)? 1'b0 : 1'b0;
  assign N16 = data_rvalid_q;
  assign N17 = N91;
  assign N243 = (N16)? N241 : 
                (N17)? 1'b0 : 1'b0;
  assign ptw_lvl_n = (N18)? { 1'b0, 1'b0 } : 
                     (N19)? { N233, N232 } : 1'b0;
  assign N18 = N28;
  assign N19 = N34;
  assign global_mapping_n = (N18)? 1'b0 : 
                            (N19)? 1'b1 : 1'b0;
  assign dtlb_miss_o = (N18)? N89 : 
                       (N20)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b0 : 1'b0;
  assign N20 = N31;
  assign N21 = N37;
  assign N22 = N40;
  assign N23 = N43;
  assign ptw_pptr_n = (N18)? { satp_ppn_i, N56, N55, N54, N53, N52, N51, N50, N49, N48, 1'b0, 1'b0, 1'b0 } : 
                      (N19)? { N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176 } : 1'b0;
  assign { N246, N245, N244 } = (N18)? { 1'b0, 1'b0, 1'b1 } : 
                                (N20)? { 1'b0, 1'b1, 1'b0 } : 
                                (N19)? { N239, 1'b0, N238 } : 
                                (N21)? { 1'b0, 1'b0, 1'b0 } : 
                                (N22)? { 1'b0, 1'b0, 1'b0 } : 
                                (N23)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign itlb_miss_o = (N18)? N88 : 
                       (N20)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b0 : 1'b0;
  assign req_port_o[13] = (N18)? 1'b0 : 
                          (N20)? 1'b1 : 
                          (N19)? 1'b0 : 
                          (N21)? 1'b0 : 
                          (N22)? 1'b0 : 
                          (N23)? 1'b0 : 1'b0;
  assign tag_valid_n = (N18)? 1'b0 : 
                       (N20)? req_port_i[65] : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b0 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b0 : 1'b0;
  assign itlb_update_o[94] = (N18)? 1'b0 : 
                             (N20)? 1'b0 : 
                             (N19)? N243 : 
                             (N21)? 1'b0 : 
                             (N22)? 1'b0 : 
                             (N23)? 1'b0 : 1'b0;
  assign dtlb_update_o[94] = (N18)? 1'b0 : 
                             (N20)? 1'b0 : 
                             (N19)? N242 : 
                             (N21)? 1'b0 : 
                             (N22)? 1'b0 : 
                             (N23)? 1'b0 : 1'b0;
  assign ptw_error_o = (N18)? 1'b0 : 
                       (N20)? 1'b0 : 
                       (N19)? 1'b0 : 
                       (N21)? 1'b1 : 
                       (N22)? 1'b0 : 
                       (N23)? 1'b0 : 1'b0;
  assign state_d = (N24)? { 1'b0, N248, N248 } : 
                   (N25)? { N246, N245, N244 } : 1'b0;
  assign N24 = flush_i;
  assign N25 = N247;
  assign itlb_update_o[5] = pte_g_ | global_mapping_q;
  assign dtlb_update_o[5] = pte_g_ | global_mapping_q;
  assign N26 = ~state_q[2];
  assign N31 = ~N30;
  assign N34 = ~N33;
  assign N37 = ~N36;
  assign N40 = ~N39;
  assign N43 = N41 | N42;
  assign N44 = N375 & N376;
  assign N375 = N373 & N374;
  assign N373 = enable_translation_i & itlb_access_i;
  assign N374 = ~itlb_hit_i;
  assign N376 = ~dtlb_access_i;
  assign N45 = N377 & N378;
  assign N377 = en_ld_st_translation_i & dtlb_access_i;
  assign N378 = ~dtlb_hit_i;
  assign N46 = N45 | N44;
  assign N47 = ~N46;
  assign N87 = ~N44;
  assign N90 = ~req_port_i[65];
  assign N91 = ~data_rvalid_q;
  assign N92 = ~pte_g_;
  assign N93 = N379 | N381;
  assign N379 = ~itlb_update_o[0];
  assign N381 = N380 & itlb_update_o[2];
  assign N380 = ~itlb_update_o[1];
  assign N94 = ~N93;
  assign N95 = itlb_update_o[1] | itlb_update_o[3];
  assign N96 = ~N95;
  assign N97 = ~walking_instr_o;
  assign N98 = N382 | N383;
  assign N382 = ~itlb_update_o[3];
  assign N383 = ~itlb_update_o[6];
  assign N100 = itlb_update_o[6] & N385;
  assign N385 = itlb_update_o[1] | N384;
  assign N384 = itlb_update_o[3] & mxr_i;
  assign N102 = lsu_is_store_i & N388;
  assign N388 = N386 | N387;
  assign N386 = ~itlb_update_o[2];
  assign N387 = ~itlb_update_o[7];
  assign N103 = ~N102;
  assign N109 = N355 & N372;
  assign N110 = N345 & N353;
  assign N111 = N110 | N109;
  assign N112 = ~N111;
  assign N247 = ~flush_i;
  assign N248 = N389 | N390;
  assign N389 = N332 & N91;
  assign N390 = N336 & req_port_i[65];
  assign N249 = ~rst_ni;
  assign N250 = N28 & N247;
  assign N251 = N47 & N250;
  assign N252 = N31 & N247;
  assign N253 = N90 & N252;
  assign N254 = N251 | N253;
  assign N255 = N34 & N247;
  assign N256 = N91 & N255;
  assign N257 = N254 | N256;
  assign N258 = N40 & N247;
  assign N259 = N91 & N258;
  assign N260 = N257 | N259;
  assign N261 = ~N260;
  assign N262 = N31 | N34;
  assign N263 = N262 | N37;
  assign N264 = N263 | N40;
  assign N265 = N264 | N43;
  assign N266 = ~N265;
  assign N267 = data_rvalid_q & N34;
  assign N268 = N93 & N267;
  assign N269 = N31 | N268;
  assign N270 = data_rvalid_q & N34;
  assign N271 = N94 & N270;
  assign N272 = N95 & N271;
  assign N273 = N269 | N272;
  assign N274 = N91 & N34;
  assign N275 = N273 | N274;
  assign N276 = N275 | N37;
  assign N277 = N276 | N40;
  assign N278 = N277 | N43;
  assign N279 = ~N278;
  assign N280 = N93 & N270;
  assign N281 = N31 | N280;
  assign N282 = N281 | N272;
  assign N283 = N282 | N274;
  assign N284 = N283 | N37;
  assign N285 = N284 | N40;
  assign N286 = N285 | N43;
  assign N287 = ~N286;
  assign N288 = N47 & N28;
  assign N289 = N288 | N31;
  assign N290 = N289 | N34;
  assign N291 = N290 | N37;
  assign N292 = N291 | N40;
  assign N293 = N292 | N43;
  assign N294 = ~N293;
  assign N295 = N289 | N280;
  assign N296 = N295 | N272;
  assign N297 = N296 | N274;
  assign N298 = N297 | N37;
  assign N299 = N298 | N40;
  assign N300 = N299 | N43;
  assign N301 = ~N300;
  assign N302 = N289 | N268;
  assign N303 = N94 & N267;
  assign N304 = N95 & N303;
  assign N305 = N302 | N304;
  assign N306 = N305 | N274;
  assign N307 = N306 | N37;
  assign N308 = N307 | N40;
  assign N309 = N308 | N43;
  assign N310 = ~N309;
  assign N311 = N92 & N267;
  assign N312 = N31 | N311;
  assign N313 = N312 | N274;
  assign N314 = N313 | N37;
  assign N315 = N314 | N40;
  assign N316 = N315 | N43;
  assign N317 = ~N316;

endmodule