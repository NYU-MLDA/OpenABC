module PMPChecker( // @[:freechips.rocketchip.system.TinyConfig.fir@103215.2]
  input         io_pmp_0_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_0_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_0_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_0_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_0_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_0_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_0_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_1_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_1_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_1_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_1_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_1_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_1_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_1_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_2_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_2_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_2_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_2_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_2_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_2_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_2_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_3_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_3_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_3_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_3_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_3_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_3_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_3_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_4_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_4_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_4_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_4_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_4_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_4_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_4_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_5_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_5_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_5_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_5_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_5_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_5_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_5_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_6_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_6_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_6_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_6_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_6_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_6_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_6_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_7_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [1:0]  io_pmp_7_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_7_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_7_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input         io_pmp_7_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [29:0] io_pmp_7_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_pmp_7_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  input  [31:0] io_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  output        io_r, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  output        io_w, // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
  output        io_x // @[:freechips.rocketchip.system.TinyConfig.fir@103218.4]
);
  wire  _T_10; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103251.4]
  wire [31:0] _T_11; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103252.4]
  wire [31:0] _T_12; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103253.4]
  wire [31:0] _T_13; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103254.4]
  wire [31:0] _T_14; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103255.4]
  wire [31:0] _T_15; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103256.4]
  wire [31:0] _T_16; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103257.4]
  wire [31:0] _T_17; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103258.4]
  wire  _T_18; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103259.4]
  wire  _T_19; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103260.4]
  wire [31:0] _T_24; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103265.4]
  wire [31:0] _T_25; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103266.4]
  wire [31:0] _T_26; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103267.4]
  wire [31:0] _T_27; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103268.4]
  wire  _T_28; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103269.4]
  wire  _T_29; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103270.4]
  wire  _T_34; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103275.4]
  wire  _T_35; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103276.4]
  wire  _T_36; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103277.4]
  wire  _T_37; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103278.4]
  wire  _T_38; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103279.4]
  wire  _T_91; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103334.4]
  wire  _T_93; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103337.4]
  wire  _T_95; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103340.4]
  wire  _T_97_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  wire  _T_97_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  wire  _T_97_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  wire  _T_98; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103344.4]
  wire [31:0] _T_103; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103349.4]
  wire [31:0] _T_104; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103350.4]
  wire [31:0] _T_105; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103351.4]
  wire  _T_106; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103352.4]
  wire  _T_107; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103353.4]
  wire [31:0] _T_112; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103358.4]
  wire [31:0] _T_113; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103359.4]
  wire [31:0] _T_114; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103360.4]
  wire [31:0] _T_115; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103361.4]
  wire  _T_116; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103362.4]
  wire  _T_117; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103363.4]
  wire  _T_123; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103369.4]
  wire  _T_124; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103370.4]
  wire  _T_125; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103371.4]
  wire  _T_126; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103372.4]
  wire  _T_179; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103427.4]
  wire  _T_181; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103430.4]
  wire  _T_183; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103433.4]
  wire  _T_185_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  wire  _T_185_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  wire  _T_185_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  wire  _T_186; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103437.4]
  wire [31:0] _T_191; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103442.4]
  wire [31:0] _T_192; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103443.4]
  wire [31:0] _T_193; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103444.4]
  wire  _T_194; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103445.4]
  wire  _T_195; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103446.4]
  wire [31:0] _T_200; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103451.4]
  wire [31:0] _T_201; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103452.4]
  wire [31:0] _T_202; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103453.4]
  wire [31:0] _T_203; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103454.4]
  wire  _T_204; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103455.4]
  wire  _T_205; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103456.4]
  wire  _T_211; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103462.4]
  wire  _T_212; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103463.4]
  wire  _T_213; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103464.4]
  wire  _T_214; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103465.4]
  wire  _T_267; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103520.4]
  wire  _T_269; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103523.4]
  wire  _T_271; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103526.4]
  wire  _T_273_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  wire  _T_273_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  wire  _T_273_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  wire  _T_274; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103530.4]
  wire [31:0] _T_279; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103535.4]
  wire [31:0] _T_280; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103536.4]
  wire [31:0] _T_281; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103537.4]
  wire  _T_282; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103538.4]
  wire  _T_283; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103539.4]
  wire [31:0] _T_288; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103544.4]
  wire [31:0] _T_289; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103545.4]
  wire [31:0] _T_290; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103546.4]
  wire [31:0] _T_291; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103547.4]
  wire  _T_292; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103548.4]
  wire  _T_293; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103549.4]
  wire  _T_299; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103555.4]
  wire  _T_300; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103556.4]
  wire  _T_301; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103557.4]
  wire  _T_302; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103558.4]
  wire  _T_355; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103613.4]
  wire  _T_357; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103616.4]
  wire  _T_359; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103619.4]
  wire  _T_361_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  wire  _T_361_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  wire  _T_361_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  wire  _T_362; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103623.4]
  wire [31:0] _T_367; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103628.4]
  wire [31:0] _T_368; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103629.4]
  wire [31:0] _T_369; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103630.4]
  wire  _T_370; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103631.4]
  wire  _T_371; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103632.4]
  wire [31:0] _T_376; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103637.4]
  wire [31:0] _T_377; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103638.4]
  wire [31:0] _T_378; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103639.4]
  wire [31:0] _T_379; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103640.4]
  wire  _T_380; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103641.4]
  wire  _T_381; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103642.4]
  wire  _T_387; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103648.4]
  wire  _T_388; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103649.4]
  wire  _T_389; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103650.4]
  wire  _T_390; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103651.4]
  wire  _T_443; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103706.4]
  wire  _T_445; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103709.4]
  wire  _T_447; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103712.4]
  wire  _T_449_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  wire  _T_449_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  wire  _T_449_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  wire  _T_450; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103716.4]
  wire [31:0] _T_455; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103721.4]
  wire [31:0] _T_456; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103722.4]
  wire [31:0] _T_457; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103723.4]
  wire  _T_458; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103724.4]
  wire  _T_459; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103725.4]
  wire [31:0] _T_464; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103730.4]
  wire [31:0] _T_465; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103731.4]
  wire [31:0] _T_466; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103732.4]
  wire [31:0] _T_467; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103733.4]
  wire  _T_468; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103734.4]
  wire  _T_469; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103735.4]
  wire  _T_475; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103741.4]
  wire  _T_476; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103742.4]
  wire  _T_477; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103743.4]
  wire  _T_478; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103744.4]
  wire  _T_531; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103799.4]
  wire  _T_533; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103802.4]
  wire  _T_535; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103805.4]
  wire  _T_537_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  wire  _T_537_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  wire  _T_537_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  wire  _T_538; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103809.4]
  wire [31:0] _T_543; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103814.4]
  wire [31:0] _T_544; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103815.4]
  wire [31:0] _T_545; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103816.4]
  wire  _T_546; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103817.4]
  wire  _T_547; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103818.4]
  wire [31:0] _T_552; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103823.4]
  wire [31:0] _T_553; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103824.4]
  wire [31:0] _T_554; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103825.4]
  wire [31:0] _T_555; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103826.4]
  wire  _T_556; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103827.4]
  wire  _T_557; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103828.4]
  wire  _T_563; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103834.4]
  wire  _T_564; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103835.4]
  wire  _T_565; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103836.4]
  wire  _T_566; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103837.4]
  wire  _T_619; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103892.4]
  wire  _T_621; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103895.4]
  wire  _T_623; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103898.4]
  wire  _T_625_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  wire  _T_625_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  wire  _T_625_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  wire  _T_626; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103902.4]
  wire [31:0] _T_631; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103907.4]
  wire [31:0] _T_632; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103908.4]
  wire [31:0] _T_633; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103909.4]
  wire  _T_634; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103910.4]
  wire  _T_635; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103911.4]
  wire  _T_652; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103928.4]
  wire  _T_653; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103929.4]
  wire  _T_654; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103930.4]
  wire  _T_707; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103985.4]
  wire  _T_709; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103988.4]
  wire  _T_711; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103991.4]
  assign _T_10 = io_pmp_7_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103251.4]
  assign _T_11 = {io_pmp_7_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103252.4]
  assign _T_12 = ~ _T_11; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103253.4]
  assign _T_13 = _T_12 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103254.4]
  assign _T_14 = ~ _T_13; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103255.4]
  assign _T_15 = io_addr ^ _T_14; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103256.4]
  assign _T_16 = ~ io_pmp_7_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103257.4]
  assign _T_17 = _T_15 & _T_16; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103258.4]
  assign _T_18 = _T_17 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103259.4]
  assign _T_19 = io_pmp_7_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103260.4]
  assign _T_24 = {io_pmp_6_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103265.4]
  assign _T_25 = ~ _T_24; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103266.4]
  assign _T_26 = _T_25 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103267.4]
  assign _T_27 = ~ _T_26; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103268.4]
  assign _T_28 = io_addr < _T_27; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103269.4]
  assign _T_29 = _T_28 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103270.4]
  assign _T_34 = io_addr < _T_14; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103275.4]
  assign _T_35 = _T_29 & _T_34; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103276.4]
  assign _T_36 = _T_19 & _T_35; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103277.4]
  assign _T_37 = _T_10 ? _T_18 : _T_36; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103278.4]
  assign _T_38 = io_pmp_7_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103279.4]
  assign _T_91 = io_pmp_7_cfg_r | _T_38; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103334.4]
  assign _T_93 = io_pmp_7_cfg_w | _T_38; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103337.4]
  assign _T_95 = io_pmp_7_cfg_x | _T_38; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103340.4]
  assign _T_97_cfg_x = _T_37 ? _T_95 : 1'h1; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  assign _T_97_cfg_w = _T_37 ? _T_93 : 1'h1; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  assign _T_97_cfg_r = _T_37 ? _T_91 : 1'h1; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103343.4]
  assign _T_98 = io_pmp_6_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103344.4]
  assign _T_103 = io_addr ^ _T_27; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103349.4]
  assign _T_104 = ~ io_pmp_6_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103350.4]
  assign _T_105 = _T_103 & _T_104; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103351.4]
  assign _T_106 = _T_105 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103352.4]
  assign _T_107 = io_pmp_6_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103353.4]
  assign _T_112 = {io_pmp_5_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103358.4]
  assign _T_113 = ~ _T_112; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103359.4]
  assign _T_114 = _T_113 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103360.4]
  assign _T_115 = ~ _T_114; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103361.4]
  assign _T_116 = io_addr < _T_115; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103362.4]
  assign _T_117 = _T_116 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103363.4]
  assign _T_123 = _T_117 & _T_28; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103369.4]
  assign _T_124 = _T_107 & _T_123; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103370.4]
  assign _T_125 = _T_98 ? _T_106 : _T_124; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103371.4]
  assign _T_126 = io_pmp_6_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103372.4]
  assign _T_179 = io_pmp_6_cfg_r | _T_126; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103427.4]
  assign _T_181 = io_pmp_6_cfg_w | _T_126; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103430.4]
  assign _T_183 = io_pmp_6_cfg_x | _T_126; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103433.4]
  assign _T_185_cfg_x = _T_125 ? _T_183 : _T_97_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  assign _T_185_cfg_w = _T_125 ? _T_181 : _T_97_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  assign _T_185_cfg_r = _T_125 ? _T_179 : _T_97_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103436.4]
  assign _T_186 = io_pmp_5_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103437.4]
  assign _T_191 = io_addr ^ _T_115; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103442.4]
  assign _T_192 = ~ io_pmp_5_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103443.4]
  assign _T_193 = _T_191 & _T_192; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103444.4]
  assign _T_194 = _T_193 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103445.4]
  assign _T_195 = io_pmp_5_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103446.4]
  assign _T_200 = {io_pmp_4_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103451.4]
  assign _T_201 = ~ _T_200; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103452.4]
  assign _T_202 = _T_201 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103453.4]
  assign _T_203 = ~ _T_202; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103454.4]
  assign _T_204 = io_addr < _T_203; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103455.4]
  assign _T_205 = _T_204 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103456.4]
  assign _T_211 = _T_205 & _T_116; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103462.4]
  assign _T_212 = _T_195 & _T_211; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103463.4]
  assign _T_213 = _T_186 ? _T_194 : _T_212; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103464.4]
  assign _T_214 = io_pmp_5_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103465.4]
  assign _T_267 = io_pmp_5_cfg_r | _T_214; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103520.4]
  assign _T_269 = io_pmp_5_cfg_w | _T_214; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103523.4]
  assign _T_271 = io_pmp_5_cfg_x | _T_214; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103526.4]
  assign _T_273_cfg_x = _T_213 ? _T_271 : _T_185_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  assign _T_273_cfg_w = _T_213 ? _T_269 : _T_185_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  assign _T_273_cfg_r = _T_213 ? _T_267 : _T_185_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103529.4]
  assign _T_274 = io_pmp_4_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103530.4]
  assign _T_279 = io_addr ^ _T_203; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103535.4]
  assign _T_280 = ~ io_pmp_4_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103536.4]
  assign _T_281 = _T_279 & _T_280; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103537.4]
  assign _T_282 = _T_281 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103538.4]
  assign _T_283 = io_pmp_4_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103539.4]
  assign _T_288 = {io_pmp_3_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103544.4]
  assign _T_289 = ~ _T_288; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103545.4]
  assign _T_290 = _T_289 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103546.4]
  assign _T_291 = ~ _T_290; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103547.4]
  assign _T_292 = io_addr < _T_291; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103548.4]
  assign _T_293 = _T_292 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103549.4]
  assign _T_299 = _T_293 & _T_204; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103555.4]
  assign _T_300 = _T_283 & _T_299; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103556.4]
  assign _T_301 = _T_274 ? _T_282 : _T_300; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103557.4]
  assign _T_302 = io_pmp_4_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103558.4]
  assign _T_355 = io_pmp_4_cfg_r | _T_302; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103613.4]
  assign _T_357 = io_pmp_4_cfg_w | _T_302; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103616.4]
  assign _T_359 = io_pmp_4_cfg_x | _T_302; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103619.4]
  assign _T_361_cfg_x = _T_301 ? _T_359 : _T_273_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  assign _T_361_cfg_w = _T_301 ? _T_357 : _T_273_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  assign _T_361_cfg_r = _T_301 ? _T_355 : _T_273_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103622.4]
  assign _T_362 = io_pmp_3_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103623.4]
  assign _T_367 = io_addr ^ _T_291; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103628.4]
  assign _T_368 = ~ io_pmp_3_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103629.4]
  assign _T_369 = _T_367 & _T_368; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103630.4]
  assign _T_370 = _T_369 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103631.4]
  assign _T_371 = io_pmp_3_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103632.4]
  assign _T_376 = {io_pmp_2_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103637.4]
  assign _T_377 = ~ _T_376; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103638.4]
  assign _T_378 = _T_377 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103639.4]
  assign _T_379 = ~ _T_378; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103640.4]
  assign _T_380 = io_addr < _T_379; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103641.4]
  assign _T_381 = _T_380 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103642.4]
  assign _T_387 = _T_381 & _T_292; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103648.4]
  assign _T_388 = _T_371 & _T_387; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103649.4]
  assign _T_389 = _T_362 ? _T_370 : _T_388; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103650.4]
  assign _T_390 = io_pmp_3_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103651.4]
  assign _T_443 = io_pmp_3_cfg_r | _T_390; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103706.4]
  assign _T_445 = io_pmp_3_cfg_w | _T_390; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103709.4]
  assign _T_447 = io_pmp_3_cfg_x | _T_390; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103712.4]
  assign _T_449_cfg_x = _T_389 ? _T_447 : _T_361_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  assign _T_449_cfg_w = _T_389 ? _T_445 : _T_361_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  assign _T_449_cfg_r = _T_389 ? _T_443 : _T_361_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103715.4]
  assign _T_450 = io_pmp_2_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103716.4]
  assign _T_455 = io_addr ^ _T_379; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103721.4]
  assign _T_456 = ~ io_pmp_2_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103722.4]
  assign _T_457 = _T_455 & _T_456; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103723.4]
  assign _T_458 = _T_457 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103724.4]
  assign _T_459 = io_pmp_2_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103725.4]
  assign _T_464 = {io_pmp_1_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103730.4]
  assign _T_465 = ~ _T_464; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103731.4]
  assign _T_466 = _T_465 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103732.4]
  assign _T_467 = ~ _T_466; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103733.4]
  assign _T_468 = io_addr < _T_467; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103734.4]
  assign _T_469 = _T_468 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103735.4]
  assign _T_475 = _T_469 & _T_380; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103741.4]
  assign _T_476 = _T_459 & _T_475; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103742.4]
  assign _T_477 = _T_450 ? _T_458 : _T_476; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103743.4]
  assign _T_478 = io_pmp_2_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103744.4]
  assign _T_531 = io_pmp_2_cfg_r | _T_478; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103799.4]
  assign _T_533 = io_pmp_2_cfg_w | _T_478; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103802.4]
  assign _T_535 = io_pmp_2_cfg_x | _T_478; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103805.4]
  assign _T_537_cfg_x = _T_477 ? _T_535 : _T_449_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  assign _T_537_cfg_w = _T_477 ? _T_533 : _T_449_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  assign _T_537_cfg_r = _T_477 ? _T_531 : _T_449_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103808.4]
  assign _T_538 = io_pmp_1_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103809.4]
  assign _T_543 = io_addr ^ _T_467; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103814.4]
  assign _T_544 = ~ io_pmp_1_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103815.4]
  assign _T_545 = _T_543 & _T_544; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103816.4]
  assign _T_546 = _T_545 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103817.4]
  assign _T_547 = io_pmp_1_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103818.4]
  assign _T_552 = {io_pmp_0_addr, 2'h0}; // @[PMP.scala 60:36:freechips.rocketchip.system.TinyConfig.fir@103823.4]
  assign _T_553 = ~ _T_552; // @[PMP.scala 60:29:freechips.rocketchip.system.TinyConfig.fir@103824.4]
  assign _T_554 = _T_553 | 32'h3; // @[PMP.scala 60:48:freechips.rocketchip.system.TinyConfig.fir@103825.4]
  assign _T_555 = ~ _T_554; // @[PMP.scala 60:27:freechips.rocketchip.system.TinyConfig.fir@103826.4]
  assign _T_556 = io_addr < _T_555; // @[PMP.scala 77:9:freechips.rocketchip.system.TinyConfig.fir@103827.4]
  assign _T_557 = _T_556 == 1'h0; // @[PMP.scala 88:5:freechips.rocketchip.system.TinyConfig.fir@103828.4]
  assign _T_563 = _T_557 & _T_468; // @[PMP.scala 94:48:freechips.rocketchip.system.TinyConfig.fir@103834.4]
  assign _T_564 = _T_547 & _T_563; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103835.4]
  assign _T_565 = _T_538 ? _T_546 : _T_564; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103836.4]
  assign _T_566 = io_pmp_1_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103837.4]
  assign _T_619 = io_pmp_1_cfg_r | _T_566; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103892.4]
  assign _T_621 = io_pmp_1_cfg_w | _T_566; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103895.4]
  assign _T_623 = io_pmp_1_cfg_x | _T_566; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103898.4]
  assign _T_625_cfg_x = _T_565 ? _T_623 : _T_537_cfg_x; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  assign _T_625_cfg_w = _T_565 ? _T_621 : _T_537_cfg_w; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  assign _T_625_cfg_r = _T_565 ? _T_619 : _T_537_cfg_r; // @[PMP.scala 184:8:freechips.rocketchip.system.TinyConfig.fir@103901.4]
  assign _T_626 = io_pmp_0_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@103902.4]
  assign _T_631 = io_addr ^ _T_555; // @[PMP.scala 63:47:freechips.rocketchip.system.TinyConfig.fir@103907.4]
  assign _T_632 = ~ io_pmp_0_mask; // @[PMP.scala 63:54:freechips.rocketchip.system.TinyConfig.fir@103908.4]
  assign _T_633 = _T_631 & _T_632; // @[PMP.scala 63:52:freechips.rocketchip.system.TinyConfig.fir@103909.4]
  assign _T_634 = _T_633 == 32'h0; // @[PMP.scala 63:58:freechips.rocketchip.system.TinyConfig.fir@103910.4]
  assign _T_635 = io_pmp_0_cfg_a[0]; // @[PMP.scala 46:26:freechips.rocketchip.system.TinyConfig.fir@103911.4]
  assign _T_652 = _T_635 & _T_556; // @[PMP.scala 132:61:freechips.rocketchip.system.TinyConfig.fir@103928.4]
  assign _T_653 = _T_626 ? _T_634 : _T_652; // @[PMP.scala 132:8:freechips.rocketchip.system.TinyConfig.fir@103929.4]
  assign _T_654 = io_pmp_0_cfg_l == 1'h0; // @[PMP.scala 163:29:freechips.rocketchip.system.TinyConfig.fir@103930.4]
  assign _T_707 = io_pmp_0_cfg_r | _T_654; // @[PMP.scala 181:40:freechips.rocketchip.system.TinyConfig.fir@103985.4]
  assign _T_709 = io_pmp_0_cfg_w | _T_654; // @[PMP.scala 182:40:freechips.rocketchip.system.TinyConfig.fir@103988.4]
  assign _T_711 = io_pmp_0_cfg_x | _T_654; // @[PMP.scala 183:40:freechips.rocketchip.system.TinyConfig.fir@103991.4]
  assign io_r = _T_653 ? _T_707 : _T_625_cfg_r; // @[PMP.scala 187:8:freechips.rocketchip.system.TinyConfig.fir@103995.4]
  assign io_w = _T_653 ? _T_709 : _T_625_cfg_w; // @[PMP.scala 188:8:freechips.rocketchip.system.TinyConfig.fir@103996.4]
  assign io_x = _T_653 ? _T_711 : _T_625_cfg_x; // @[PMP.scala 189:8:freechips.rocketchip.system.TinyConfig.fir@103997.4]
endmodule