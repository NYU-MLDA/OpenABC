module bp_accelerator_complex_05
(
  core_clk_i,
  core_reset_i,
  coh_clk_i,
  coh_reset_i,
  coh_req_link_i,
  coh_req_link_o,
  coh_cmd_link_i,
  coh_cmd_link_o,
  coh_resp_link_i,
  coh_resp_link_o
);

  input [259:0] coh_req_link_i;
  output [259:0] coh_req_link_o;
  input [259:0] coh_cmd_link_i;
  output [259:0] coh_cmd_link_o;
  input [259:0] coh_resp_link_i;
  output [259:0] coh_resp_link_o;
  input core_clk_i;
  input core_reset_i;
  input coh_clk_i;
  input coh_reset_i;
  wire [259:0] coh_req_link_o,coh_cmd_link_o,coh_resp_link_o;
  assign coh_resp_link_o[0] = 1'b0;
  assign coh_resp_link_o[1] = 1'b0;
  assign coh_resp_link_o[2] = 1'b0;
  assign coh_resp_link_o[3] = 1'b0;
  assign coh_resp_link_o[4] = 1'b0;
  assign coh_resp_link_o[5] = 1'b0;
  assign coh_resp_link_o[6] = 1'b0;
  assign coh_resp_link_o[7] = 1'b0;
  assign coh_resp_link_o[8] = 1'b0;
  assign coh_resp_link_o[9] = 1'b0;
  assign coh_resp_link_o[10] = 1'b0;
  assign coh_resp_link_o[11] = 1'b0;
  assign coh_resp_link_o[12] = 1'b0;
  assign coh_resp_link_o[13] = 1'b0;
  assign coh_resp_link_o[14] = 1'b0;
  assign coh_resp_link_o[15] = 1'b0;
  assign coh_resp_link_o[16] = 1'b0;
  assign coh_resp_link_o[17] = 1'b0;
  assign coh_resp_link_o[18] = 1'b0;
  assign coh_resp_link_o[19] = 1'b0;
  assign coh_resp_link_o[20] = 1'b0;
  assign coh_resp_link_o[21] = 1'b0;
  assign coh_resp_link_o[22] = 1'b0;
  assign coh_resp_link_o[23] = 1'b0;
  assign coh_resp_link_o[24] = 1'b0;
  assign coh_resp_link_o[25] = 1'b0;
  assign coh_resp_link_o[26] = 1'b0;
  assign coh_resp_link_o[27] = 1'b0;
  assign coh_resp_link_o[28] = 1'b0;
  assign coh_resp_link_o[29] = 1'b0;
  assign coh_resp_link_o[30] = 1'b0;
  assign coh_resp_link_o[31] = 1'b0;
  assign coh_resp_link_o[32] = 1'b0;
  assign coh_resp_link_o[33] = 1'b0;
  assign coh_resp_link_o[34] = 1'b0;
  assign coh_resp_link_o[35] = 1'b0;
  assign coh_resp_link_o[36] = 1'b0;
  assign coh_resp_link_o[37] = 1'b0;
  assign coh_resp_link_o[38] = 1'b0;
  assign coh_resp_link_o[39] = 1'b0;
  assign coh_resp_link_o[40] = 1'b0;
  assign coh_resp_link_o[41] = 1'b0;
  assign coh_resp_link_o[42] = 1'b0;
  assign coh_resp_link_o[43] = 1'b0;
  assign coh_resp_link_o[44] = 1'b0;
  assign coh_resp_link_o[45] = 1'b0;
  assign coh_resp_link_o[46] = 1'b0;
  assign coh_resp_link_o[47] = 1'b0;
  assign coh_resp_link_o[48] = 1'b0;
  assign coh_resp_link_o[49] = 1'b0;
  assign coh_resp_link_o[50] = 1'b0;
  assign coh_resp_link_o[51] = 1'b0;
  assign coh_resp_link_o[52] = 1'b0;
  assign coh_resp_link_o[53] = 1'b0;
  assign coh_resp_link_o[54] = 1'b0;
  assign coh_resp_link_o[55] = 1'b0;
  assign coh_resp_link_o[56] = 1'b0;
  assign coh_resp_link_o[57] = 1'b0;
  assign coh_resp_link_o[58] = 1'b0;
  assign coh_resp_link_o[59] = 1'b0;
  assign coh_resp_link_o[60] = 1'b0;
  assign coh_resp_link_o[61] = 1'b0;
  assign coh_resp_link_o[62] = 1'b0;
  assign coh_resp_link_o[63] = 1'b0;
  assign coh_resp_link_o[64] = 1'b0;
  assign coh_resp_link_o[65] = 1'b0;
  assign coh_resp_link_o[66] = 1'b0;
  assign coh_resp_link_o[67] = 1'b0;
  assign coh_resp_link_o[68] = 1'b0;
  assign coh_resp_link_o[69] = 1'b0;
  assign coh_resp_link_o[70] = 1'b0;
  assign coh_resp_link_o[71] = 1'b0;
  assign coh_resp_link_o[72] = 1'b0;
  assign coh_resp_link_o[73] = 1'b0;
  assign coh_resp_link_o[74] = 1'b0;
  assign coh_resp_link_o[75] = 1'b0;
  assign coh_resp_link_o[76] = 1'b0;
  assign coh_resp_link_o[77] = 1'b0;
  assign coh_resp_link_o[78] = 1'b0;
  assign coh_resp_link_o[79] = 1'b0;
  assign coh_resp_link_o[80] = 1'b0;
  assign coh_resp_link_o[81] = 1'b0;
  assign coh_resp_link_o[82] = 1'b0;
  assign coh_resp_link_o[83] = 1'b0;
  assign coh_resp_link_o[84] = 1'b0;
  assign coh_resp_link_o[85] = 1'b0;
  assign coh_resp_link_o[86] = 1'b0;
  assign coh_resp_link_o[87] = 1'b0;
  assign coh_resp_link_o[88] = 1'b0;
  assign coh_resp_link_o[89] = 1'b0;
  assign coh_resp_link_o[90] = 1'b0;
  assign coh_resp_link_o[91] = 1'b0;
  assign coh_resp_link_o[92] = 1'b0;
  assign coh_resp_link_o[93] = 1'b0;
  assign coh_resp_link_o[94] = 1'b0;
  assign coh_resp_link_o[95] = 1'b0;
  assign coh_resp_link_o[96] = 1'b0;
  assign coh_resp_link_o[97] = 1'b0;
  assign coh_resp_link_o[98] = 1'b0;
  assign coh_resp_link_o[99] = 1'b0;
  assign coh_resp_link_o[100] = 1'b0;
  assign coh_resp_link_o[101] = 1'b0;
  assign coh_resp_link_o[102] = 1'b0;
  assign coh_resp_link_o[103] = 1'b0;
  assign coh_resp_link_o[104] = 1'b0;
  assign coh_resp_link_o[105] = 1'b0;
  assign coh_resp_link_o[106] = 1'b0;
  assign coh_resp_link_o[107] = 1'b0;
  assign coh_resp_link_o[108] = 1'b0;
  assign coh_resp_link_o[109] = 1'b0;
  assign coh_resp_link_o[110] = 1'b0;
  assign coh_resp_link_o[111] = 1'b0;
  assign coh_resp_link_o[112] = 1'b0;
  assign coh_resp_link_o[113] = 1'b0;
  assign coh_resp_link_o[114] = 1'b0;
  assign coh_resp_link_o[115] = 1'b0;
  assign coh_resp_link_o[116] = 1'b0;
  assign coh_resp_link_o[117] = 1'b0;
  assign coh_resp_link_o[118] = 1'b0;
  assign coh_resp_link_o[119] = 1'b0;
  assign coh_resp_link_o[120] = 1'b0;
  assign coh_resp_link_o[121] = 1'b0;
  assign coh_resp_link_o[122] = 1'b0;
  assign coh_resp_link_o[123] = 1'b0;
  assign coh_resp_link_o[124] = 1'b0;
  assign coh_resp_link_o[125] = 1'b0;
  assign coh_resp_link_o[126] = 1'b0;
  assign coh_resp_link_o[127] = 1'b0;
  assign coh_resp_link_o[128] = 1'b0;
  assign coh_resp_link_o[129] = 1'b0;
  assign coh_resp_link_o[130] = 1'b0;
  assign coh_resp_link_o[131] = 1'b0;
  assign coh_resp_link_o[132] = 1'b0;
  assign coh_resp_link_o[133] = 1'b0;
  assign coh_resp_link_o[134] = 1'b0;
  assign coh_resp_link_o[135] = 1'b0;
  assign coh_resp_link_o[136] = 1'b0;
  assign coh_resp_link_o[137] = 1'b0;
  assign coh_resp_link_o[138] = 1'b0;
  assign coh_resp_link_o[139] = 1'b0;
  assign coh_resp_link_o[140] = 1'b0;
  assign coh_resp_link_o[141] = 1'b0;
  assign coh_resp_link_o[142] = 1'b0;
  assign coh_resp_link_o[143] = 1'b0;
  assign coh_resp_link_o[144] = 1'b0;
  assign coh_resp_link_o[145] = 1'b0;
  assign coh_resp_link_o[146] = 1'b0;
  assign coh_resp_link_o[147] = 1'b0;
  assign coh_resp_link_o[148] = 1'b0;
  assign coh_resp_link_o[149] = 1'b0;
  assign coh_resp_link_o[150] = 1'b0;
  assign coh_resp_link_o[151] = 1'b0;
  assign coh_resp_link_o[152] = 1'b0;
  assign coh_resp_link_o[153] = 1'b0;
  assign coh_resp_link_o[154] = 1'b0;
  assign coh_resp_link_o[155] = 1'b0;
  assign coh_resp_link_o[156] = 1'b0;
  assign coh_resp_link_o[157] = 1'b0;
  assign coh_resp_link_o[158] = 1'b0;
  assign coh_resp_link_o[159] = 1'b0;
  assign coh_resp_link_o[160] = 1'b0;
  assign coh_resp_link_o[161] = 1'b0;
  assign coh_resp_link_o[162] = 1'b0;
  assign coh_resp_link_o[163] = 1'b0;
  assign coh_resp_link_o[164] = 1'b0;
  assign coh_resp_link_o[165] = 1'b0;
  assign coh_resp_link_o[166] = 1'b0;
  assign coh_resp_link_o[167] = 1'b0;
  assign coh_resp_link_o[168] = 1'b0;
  assign coh_resp_link_o[169] = 1'b0;
  assign coh_resp_link_o[170] = 1'b0;
  assign coh_resp_link_o[171] = 1'b0;
  assign coh_resp_link_o[172] = 1'b0;
  assign coh_resp_link_o[173] = 1'b0;
  assign coh_resp_link_o[174] = 1'b0;
  assign coh_resp_link_o[175] = 1'b0;
  assign coh_resp_link_o[176] = 1'b0;
  assign coh_resp_link_o[177] = 1'b0;
  assign coh_resp_link_o[178] = 1'b0;
  assign coh_resp_link_o[179] = 1'b0;
  assign coh_resp_link_o[180] = 1'b0;
  assign coh_resp_link_o[181] = 1'b0;
  assign coh_resp_link_o[182] = 1'b0;
  assign coh_resp_link_o[183] = 1'b0;
  assign coh_resp_link_o[184] = 1'b0;
  assign coh_resp_link_o[185] = 1'b0;
  assign coh_resp_link_o[186] = 1'b0;
  assign coh_resp_link_o[187] = 1'b0;
  assign coh_resp_link_o[188] = 1'b0;
  assign coh_resp_link_o[189] = 1'b0;
  assign coh_resp_link_o[190] = 1'b0;
  assign coh_resp_link_o[191] = 1'b0;
  assign coh_resp_link_o[192] = 1'b0;
  assign coh_resp_link_o[193] = 1'b0;
  assign coh_resp_link_o[194] = 1'b0;
  assign coh_resp_link_o[195] = 1'b0;
  assign coh_resp_link_o[196] = 1'b0;
  assign coh_resp_link_o[197] = 1'b0;
  assign coh_resp_link_o[198] = 1'b0;
  assign coh_resp_link_o[199] = 1'b0;
  assign coh_resp_link_o[200] = 1'b0;
  assign coh_resp_link_o[201] = 1'b0;
  assign coh_resp_link_o[202] = 1'b0;
  assign coh_resp_link_o[203] = 1'b0;
  assign coh_resp_link_o[204] = 1'b0;
  assign coh_resp_link_o[205] = 1'b0;
  assign coh_resp_link_o[206] = 1'b0;
  assign coh_resp_link_o[207] = 1'b0;
  assign coh_resp_link_o[208] = 1'b0;
  assign coh_resp_link_o[209] = 1'b0;
  assign coh_resp_link_o[210] = 1'b0;
  assign coh_resp_link_o[211] = 1'b0;
  assign coh_resp_link_o[212] = 1'b0;
  assign coh_resp_link_o[213] = 1'b0;
  assign coh_resp_link_o[214] = 1'b0;
  assign coh_resp_link_o[215] = 1'b0;
  assign coh_resp_link_o[216] = 1'b0;
  assign coh_resp_link_o[217] = 1'b0;
  assign coh_resp_link_o[218] = 1'b0;
  assign coh_resp_link_o[219] = 1'b0;
  assign coh_resp_link_o[220] = 1'b0;
  assign coh_resp_link_o[221] = 1'b0;
  assign coh_resp_link_o[222] = 1'b0;
  assign coh_resp_link_o[223] = 1'b0;
  assign coh_resp_link_o[224] = 1'b0;
  assign coh_resp_link_o[225] = 1'b0;
  assign coh_resp_link_o[226] = 1'b0;
  assign coh_resp_link_o[227] = 1'b0;
  assign coh_resp_link_o[228] = 1'b0;
  assign coh_resp_link_o[229] = 1'b0;
  assign coh_resp_link_o[230] = 1'b0;
  assign coh_resp_link_o[231] = 1'b0;
  assign coh_resp_link_o[232] = 1'b0;
  assign coh_resp_link_o[233] = 1'b0;
  assign coh_resp_link_o[234] = 1'b0;
  assign coh_resp_link_o[235] = 1'b0;
  assign coh_resp_link_o[236] = 1'b0;
  assign coh_resp_link_o[237] = 1'b0;
  assign coh_resp_link_o[238] = 1'b0;
  assign coh_resp_link_o[239] = 1'b0;
  assign coh_resp_link_o[240] = 1'b0;
  assign coh_resp_link_o[241] = 1'b0;
  assign coh_resp_link_o[242] = 1'b0;
  assign coh_resp_link_o[243] = 1'b0;
  assign coh_resp_link_o[244] = 1'b0;
  assign coh_resp_link_o[245] = 1'b0;
  assign coh_resp_link_o[246] = 1'b0;
  assign coh_resp_link_o[247] = 1'b0;
  assign coh_resp_link_o[248] = 1'b0;
  assign coh_resp_link_o[249] = 1'b0;
  assign coh_resp_link_o[250] = 1'b0;
  assign coh_resp_link_o[251] = 1'b0;
  assign coh_resp_link_o[252] = 1'b0;
  assign coh_resp_link_o[253] = 1'b0;
  assign coh_resp_link_o[254] = 1'b0;
  assign coh_resp_link_o[255] = 1'b0;
  assign coh_resp_link_o[256] = 1'b0;
  assign coh_resp_link_o[257] = 1'b0;
  assign coh_resp_link_o[258] = 1'b0;
  assign coh_resp_link_o[259] = 1'b0;
  assign coh_cmd_link_o[0] = 1'b0;
  assign coh_cmd_link_o[1] = 1'b0;
  assign coh_cmd_link_o[2] = 1'b0;
  assign coh_cmd_link_o[3] = 1'b0;
  assign coh_cmd_link_o[4] = 1'b0;
  assign coh_cmd_link_o[5] = 1'b0;
  assign coh_cmd_link_o[6] = 1'b0;
  assign coh_cmd_link_o[7] = 1'b0;
  assign coh_cmd_link_o[8] = 1'b0;
  assign coh_cmd_link_o[9] = 1'b0;
  assign coh_cmd_link_o[10] = 1'b0;
  assign coh_cmd_link_o[11] = 1'b0;
  assign coh_cmd_link_o[12] = 1'b0;
  assign coh_cmd_link_o[13] = 1'b0;
  assign coh_cmd_link_o[14] = 1'b0;
  assign coh_cmd_link_o[15] = 1'b0;
  assign coh_cmd_link_o[16] = 1'b0;
  assign coh_cmd_link_o[17] = 1'b0;
  assign coh_cmd_link_o[18] = 1'b0;
  assign coh_cmd_link_o[19] = 1'b0;
  assign coh_cmd_link_o[20] = 1'b0;
  assign coh_cmd_link_o[21] = 1'b0;
  assign coh_cmd_link_o[22] = 1'b0;
  assign coh_cmd_link_o[23] = 1'b0;
  assign coh_cmd_link_o[24] = 1'b0;
  assign coh_cmd_link_o[25] = 1'b0;
  assign coh_cmd_link_o[26] = 1'b0;
  assign coh_cmd_link_o[27] = 1'b0;
  assign coh_cmd_link_o[28] = 1'b0;
  assign coh_cmd_link_o[29] = 1'b0;
  assign coh_cmd_link_o[30] = 1'b0;
  assign coh_cmd_link_o[31] = 1'b0;
  assign coh_cmd_link_o[32] = 1'b0;
  assign coh_cmd_link_o[33] = 1'b0;
  assign coh_cmd_link_o[34] = 1'b0;
  assign coh_cmd_link_o[35] = 1'b0;
  assign coh_cmd_link_o[36] = 1'b0;
  assign coh_cmd_link_o[37] = 1'b0;
  assign coh_cmd_link_o[38] = 1'b0;
  assign coh_cmd_link_o[39] = 1'b0;
  assign coh_cmd_link_o[40] = 1'b0;
  assign coh_cmd_link_o[41] = 1'b0;
  assign coh_cmd_link_o[42] = 1'b0;
  assign coh_cmd_link_o[43] = 1'b0;
  assign coh_cmd_link_o[44] = 1'b0;
  assign coh_cmd_link_o[45] = 1'b0;
  assign coh_cmd_link_o[46] = 1'b0;
  assign coh_cmd_link_o[47] = 1'b0;
  assign coh_cmd_link_o[48] = 1'b0;
  assign coh_cmd_link_o[49] = 1'b0;
  assign coh_cmd_link_o[50] = 1'b0;
  assign coh_cmd_link_o[51] = 1'b0;
  assign coh_cmd_link_o[52] = 1'b0;
  assign coh_cmd_link_o[53] = 1'b0;
  assign coh_cmd_link_o[54] = 1'b0;
  assign coh_cmd_link_o[55] = 1'b0;
  assign coh_cmd_link_o[56] = 1'b0;
  assign coh_cmd_link_o[57] = 1'b0;
  assign coh_cmd_link_o[58] = 1'b0;
  assign coh_cmd_link_o[59] = 1'b0;
  assign coh_cmd_link_o[60] = 1'b0;
  assign coh_cmd_link_o[61] = 1'b0;
  assign coh_cmd_link_o[62] = 1'b0;
  assign coh_cmd_link_o[63] = 1'b0;
  assign coh_cmd_link_o[64] = 1'b0;
  assign coh_cmd_link_o[65] = 1'b0;
  assign coh_cmd_link_o[66] = 1'b0;
  assign coh_cmd_link_o[67] = 1'b0;
  assign coh_cmd_link_o[68] = 1'b0;
  assign coh_cmd_link_o[69] = 1'b0;
  assign coh_cmd_link_o[70] = 1'b0;
  assign coh_cmd_link_o[71] = 1'b0;
  assign coh_cmd_link_o[72] = 1'b0;
  assign coh_cmd_link_o[73] = 1'b0;
  assign coh_cmd_link_o[74] = 1'b0;
  assign coh_cmd_link_o[75] = 1'b0;
  assign coh_cmd_link_o[76] = 1'b0;
  assign coh_cmd_link_o[77] = 1'b0;
  assign coh_cmd_link_o[78] = 1'b0;
  assign coh_cmd_link_o[79] = 1'b0;
  assign coh_cmd_link_o[80] = 1'b0;
  assign coh_cmd_link_o[81] = 1'b0;
  assign coh_cmd_link_o[82] = 1'b0;
  assign coh_cmd_link_o[83] = 1'b0;
  assign coh_cmd_link_o[84] = 1'b0;
  assign coh_cmd_link_o[85] = 1'b0;
  assign coh_cmd_link_o[86] = 1'b0;
  assign coh_cmd_link_o[87] = 1'b0;
  assign coh_cmd_link_o[88] = 1'b0;
  assign coh_cmd_link_o[89] = 1'b0;
  assign coh_cmd_link_o[90] = 1'b0;
  assign coh_cmd_link_o[91] = 1'b0;
  assign coh_cmd_link_o[92] = 1'b0;
  assign coh_cmd_link_o[93] = 1'b0;
  assign coh_cmd_link_o[94] = 1'b0;
  assign coh_cmd_link_o[95] = 1'b0;
  assign coh_cmd_link_o[96] = 1'b0;
  assign coh_cmd_link_o[97] = 1'b0;
  assign coh_cmd_link_o[98] = 1'b0;
  assign coh_cmd_link_o[99] = 1'b0;
  assign coh_cmd_link_o[100] = 1'b0;
  assign coh_cmd_link_o[101] = 1'b0;
  assign coh_cmd_link_o[102] = 1'b0;
  assign coh_cmd_link_o[103] = 1'b0;
  assign coh_cmd_link_o[104] = 1'b0;
  assign coh_cmd_link_o[105] = 1'b0;
  assign coh_cmd_link_o[106] = 1'b0;
  assign coh_cmd_link_o[107] = 1'b0;
  assign coh_cmd_link_o[108] = 1'b0;
  assign coh_cmd_link_o[109] = 1'b0;
  assign coh_cmd_link_o[110] = 1'b0;
  assign coh_cmd_link_o[111] = 1'b0;
  assign coh_cmd_link_o[112] = 1'b0;
  assign coh_cmd_link_o[113] = 1'b0;
  assign coh_cmd_link_o[114] = 1'b0;
  assign coh_cmd_link_o[115] = 1'b0;
  assign coh_cmd_link_o[116] = 1'b0;
  assign coh_cmd_link_o[117] = 1'b0;
  assign coh_cmd_link_o[118] = 1'b0;
  assign coh_cmd_link_o[119] = 1'b0;
  assign coh_cmd_link_o[120] = 1'b0;
  assign coh_cmd_link_o[121] = 1'b0;
  assign coh_cmd_link_o[122] = 1'b0;
  assign coh_cmd_link_o[123] = 1'b0;
  assign coh_cmd_link_o[124] = 1'b0;
  assign coh_cmd_link_o[125] = 1'b0;
  assign coh_cmd_link_o[126] = 1'b0;
  assign coh_cmd_link_o[127] = 1'b0;
  assign coh_cmd_link_o[128] = 1'b0;
  assign coh_cmd_link_o[129] = 1'b0;
  assign coh_cmd_link_o[130] = 1'b0;
  assign coh_cmd_link_o[131] = 1'b0;
  assign coh_cmd_link_o[132] = 1'b0;
  assign coh_cmd_link_o[133] = 1'b0;
  assign coh_cmd_link_o[134] = 1'b0;
  assign coh_cmd_link_o[135] = 1'b0;
  assign coh_cmd_link_o[136] = 1'b0;
  assign coh_cmd_link_o[137] = 1'b0;
  assign coh_cmd_link_o[138] = 1'b0;
  assign coh_cmd_link_o[139] = 1'b0;
  assign coh_cmd_link_o[140] = 1'b0;
  assign coh_cmd_link_o[141] = 1'b0;
  assign coh_cmd_link_o[142] = 1'b0;
  assign coh_cmd_link_o[143] = 1'b0;
  assign coh_cmd_link_o[144] = 1'b0;
  assign coh_cmd_link_o[145] = 1'b0;
  assign coh_cmd_link_o[146] = 1'b0;
  assign coh_cmd_link_o[147] = 1'b0;
  assign coh_cmd_link_o[148] = 1'b0;
  assign coh_cmd_link_o[149] = 1'b0;
  assign coh_cmd_link_o[150] = 1'b0;
  assign coh_cmd_link_o[151] = 1'b0;
  assign coh_cmd_link_o[152] = 1'b0;
  assign coh_cmd_link_o[153] = 1'b0;
  assign coh_cmd_link_o[154] = 1'b0;
  assign coh_cmd_link_o[155] = 1'b0;
  assign coh_cmd_link_o[156] = 1'b0;
  assign coh_cmd_link_o[157] = 1'b0;
  assign coh_cmd_link_o[158] = 1'b0;
  assign coh_cmd_link_o[159] = 1'b0;
  assign coh_cmd_link_o[160] = 1'b0;
  assign coh_cmd_link_o[161] = 1'b0;
  assign coh_cmd_link_o[162] = 1'b0;
  assign coh_cmd_link_o[163] = 1'b0;
  assign coh_cmd_link_o[164] = 1'b0;
  assign coh_cmd_link_o[165] = 1'b0;
  assign coh_cmd_link_o[166] = 1'b0;
  assign coh_cmd_link_o[167] = 1'b0;
  assign coh_cmd_link_o[168] = 1'b0;
  assign coh_cmd_link_o[169] = 1'b0;
  assign coh_cmd_link_o[170] = 1'b0;
  assign coh_cmd_link_o[171] = 1'b0;
  assign coh_cmd_link_o[172] = 1'b0;
  assign coh_cmd_link_o[173] = 1'b0;
  assign coh_cmd_link_o[174] = 1'b0;
  assign coh_cmd_link_o[175] = 1'b0;
  assign coh_cmd_link_o[176] = 1'b0;
  assign coh_cmd_link_o[177] = 1'b0;
  assign coh_cmd_link_o[178] = 1'b0;
  assign coh_cmd_link_o[179] = 1'b0;
  assign coh_cmd_link_o[180] = 1'b0;
  assign coh_cmd_link_o[181] = 1'b0;
  assign coh_cmd_link_o[182] = 1'b0;
  assign coh_cmd_link_o[183] = 1'b0;
  assign coh_cmd_link_o[184] = 1'b0;
  assign coh_cmd_link_o[185] = 1'b0;
  assign coh_cmd_link_o[186] = 1'b0;
  assign coh_cmd_link_o[187] = 1'b0;
  assign coh_cmd_link_o[188] = 1'b0;
  assign coh_cmd_link_o[189] = 1'b0;
  assign coh_cmd_link_o[190] = 1'b0;
  assign coh_cmd_link_o[191] = 1'b0;
  assign coh_cmd_link_o[192] = 1'b0;
  assign coh_cmd_link_o[193] = 1'b0;
  assign coh_cmd_link_o[194] = 1'b0;
  assign coh_cmd_link_o[195] = 1'b0;
  assign coh_cmd_link_o[196] = 1'b0;
  assign coh_cmd_link_o[197] = 1'b0;
  assign coh_cmd_link_o[198] = 1'b0;
  assign coh_cmd_link_o[199] = 1'b0;
  assign coh_cmd_link_o[200] = 1'b0;
  assign coh_cmd_link_o[201] = 1'b0;
  assign coh_cmd_link_o[202] = 1'b0;
  assign coh_cmd_link_o[203] = 1'b0;
  assign coh_cmd_link_o[204] = 1'b0;
  assign coh_cmd_link_o[205] = 1'b0;
  assign coh_cmd_link_o[206] = 1'b0;
  assign coh_cmd_link_o[207] = 1'b0;
  assign coh_cmd_link_o[208] = 1'b0;
  assign coh_cmd_link_o[209] = 1'b0;
  assign coh_cmd_link_o[210] = 1'b0;
  assign coh_cmd_link_o[211] = 1'b0;
  assign coh_cmd_link_o[212] = 1'b0;
  assign coh_cmd_link_o[213] = 1'b0;
  assign coh_cmd_link_o[214] = 1'b0;
  assign coh_cmd_link_o[215] = 1'b0;
  assign coh_cmd_link_o[216] = 1'b0;
  assign coh_cmd_link_o[217] = 1'b0;
  assign coh_cmd_link_o[218] = 1'b0;
  assign coh_cmd_link_o[219] = 1'b0;
  assign coh_cmd_link_o[220] = 1'b0;
  assign coh_cmd_link_o[221] = 1'b0;
  assign coh_cmd_link_o[222] = 1'b0;
  assign coh_cmd_link_o[223] = 1'b0;
  assign coh_cmd_link_o[224] = 1'b0;
  assign coh_cmd_link_o[225] = 1'b0;
  assign coh_cmd_link_o[226] = 1'b0;
  assign coh_cmd_link_o[227] = 1'b0;
  assign coh_cmd_link_o[228] = 1'b0;
  assign coh_cmd_link_o[229] = 1'b0;
  assign coh_cmd_link_o[230] = 1'b0;
  assign coh_cmd_link_o[231] = 1'b0;
  assign coh_cmd_link_o[232] = 1'b0;
  assign coh_cmd_link_o[233] = 1'b0;
  assign coh_cmd_link_o[234] = 1'b0;
  assign coh_cmd_link_o[235] = 1'b0;
  assign coh_cmd_link_o[236] = 1'b0;
  assign coh_cmd_link_o[237] = 1'b0;
  assign coh_cmd_link_o[238] = 1'b0;
  assign coh_cmd_link_o[239] = 1'b0;
  assign coh_cmd_link_o[240] = 1'b0;
  assign coh_cmd_link_o[241] = 1'b0;
  assign coh_cmd_link_o[242] = 1'b0;
  assign coh_cmd_link_o[243] = 1'b0;
  assign coh_cmd_link_o[244] = 1'b0;
  assign coh_cmd_link_o[245] = 1'b0;
  assign coh_cmd_link_o[246] = 1'b0;
  assign coh_cmd_link_o[247] = 1'b0;
  assign coh_cmd_link_o[248] = 1'b0;
  assign coh_cmd_link_o[249] = 1'b0;
  assign coh_cmd_link_o[250] = 1'b0;
  assign coh_cmd_link_o[251] = 1'b0;
  assign coh_cmd_link_o[252] = 1'b0;
  assign coh_cmd_link_o[253] = 1'b0;
  assign coh_cmd_link_o[254] = 1'b0;
  assign coh_cmd_link_o[255] = 1'b0;
  assign coh_cmd_link_o[256] = 1'b0;
  assign coh_cmd_link_o[257] = 1'b0;
  assign coh_cmd_link_o[258] = 1'b0;
  assign coh_cmd_link_o[259] = 1'b0;
  assign coh_req_link_o[0] = 1'b0;
  assign coh_req_link_o[1] = 1'b0;
  assign coh_req_link_o[2] = 1'b0;
  assign coh_req_link_o[3] = 1'b0;
  assign coh_req_link_o[4] = 1'b0;
  assign coh_req_link_o[5] = 1'b0;
  assign coh_req_link_o[6] = 1'b0;
  assign coh_req_link_o[7] = 1'b0;
  assign coh_req_link_o[8] = 1'b0;
  assign coh_req_link_o[9] = 1'b0;
  assign coh_req_link_o[10] = 1'b0;
  assign coh_req_link_o[11] = 1'b0;
  assign coh_req_link_o[12] = 1'b0;
  assign coh_req_link_o[13] = 1'b0;
  assign coh_req_link_o[14] = 1'b0;
  assign coh_req_link_o[15] = 1'b0;
  assign coh_req_link_o[16] = 1'b0;
  assign coh_req_link_o[17] = 1'b0;
  assign coh_req_link_o[18] = 1'b0;
  assign coh_req_link_o[19] = 1'b0;
  assign coh_req_link_o[20] = 1'b0;
  assign coh_req_link_o[21] = 1'b0;
  assign coh_req_link_o[22] = 1'b0;
  assign coh_req_link_o[23] = 1'b0;
  assign coh_req_link_o[24] = 1'b0;
  assign coh_req_link_o[25] = 1'b0;
  assign coh_req_link_o[26] = 1'b0;
  assign coh_req_link_o[27] = 1'b0;
  assign coh_req_link_o[28] = 1'b0;
  assign coh_req_link_o[29] = 1'b0;
  assign coh_req_link_o[30] = 1'b0;
  assign coh_req_link_o[31] = 1'b0;
  assign coh_req_link_o[32] = 1'b0;
  assign coh_req_link_o[33] = 1'b0;
  assign coh_req_link_o[34] = 1'b0;
  assign coh_req_link_o[35] = 1'b0;
  assign coh_req_link_o[36] = 1'b0;
  assign coh_req_link_o[37] = 1'b0;
  assign coh_req_link_o[38] = 1'b0;
  assign coh_req_link_o[39] = 1'b0;
  assign coh_req_link_o[40] = 1'b0;
  assign coh_req_link_o[41] = 1'b0;
  assign coh_req_link_o[42] = 1'b0;
  assign coh_req_link_o[43] = 1'b0;
  assign coh_req_link_o[44] = 1'b0;
  assign coh_req_link_o[45] = 1'b0;
  assign coh_req_link_o[46] = 1'b0;
  assign coh_req_link_o[47] = 1'b0;
  assign coh_req_link_o[48] = 1'b0;
  assign coh_req_link_o[49] = 1'b0;
  assign coh_req_link_o[50] = 1'b0;
  assign coh_req_link_o[51] = 1'b0;
  assign coh_req_link_o[52] = 1'b0;
  assign coh_req_link_o[53] = 1'b0;
  assign coh_req_link_o[54] = 1'b0;
  assign coh_req_link_o[55] = 1'b0;
  assign coh_req_link_o[56] = 1'b0;
  assign coh_req_link_o[57] = 1'b0;
  assign coh_req_link_o[58] = 1'b0;
  assign coh_req_link_o[59] = 1'b0;
  assign coh_req_link_o[60] = 1'b0;
  assign coh_req_link_o[61] = 1'b0;
  assign coh_req_link_o[62] = 1'b0;
  assign coh_req_link_o[63] = 1'b0;
  assign coh_req_link_o[64] = 1'b0;
  assign coh_req_link_o[65] = 1'b0;
  assign coh_req_link_o[66] = 1'b0;
  assign coh_req_link_o[67] = 1'b0;
  assign coh_req_link_o[68] = 1'b0;
  assign coh_req_link_o[69] = 1'b0;
  assign coh_req_link_o[70] = 1'b0;
  assign coh_req_link_o[71] = 1'b0;
  assign coh_req_link_o[72] = 1'b0;
  assign coh_req_link_o[73] = 1'b0;
  assign coh_req_link_o[74] = 1'b0;
  assign coh_req_link_o[75] = 1'b0;
  assign coh_req_link_o[76] = 1'b0;
  assign coh_req_link_o[77] = 1'b0;
  assign coh_req_link_o[78] = 1'b0;
  assign coh_req_link_o[79] = 1'b0;
  assign coh_req_link_o[80] = 1'b0;
  assign coh_req_link_o[81] = 1'b0;
  assign coh_req_link_o[82] = 1'b0;
  assign coh_req_link_o[83] = 1'b0;
  assign coh_req_link_o[84] = 1'b0;
  assign coh_req_link_o[85] = 1'b0;
  assign coh_req_link_o[86] = 1'b0;
  assign coh_req_link_o[87] = 1'b0;
  assign coh_req_link_o[88] = 1'b0;
  assign coh_req_link_o[89] = 1'b0;
  assign coh_req_link_o[90] = 1'b0;
  assign coh_req_link_o[91] = 1'b0;
  assign coh_req_link_o[92] = 1'b0;
  assign coh_req_link_o[93] = 1'b0;
  assign coh_req_link_o[94] = 1'b0;
  assign coh_req_link_o[95] = 1'b0;
  assign coh_req_link_o[96] = 1'b0;
  assign coh_req_link_o[97] = 1'b0;
  assign coh_req_link_o[98] = 1'b0;
  assign coh_req_link_o[99] = 1'b0;
  assign coh_req_link_o[100] = 1'b0;
  assign coh_req_link_o[101] = 1'b0;
  assign coh_req_link_o[102] = 1'b0;
  assign coh_req_link_o[103] = 1'b0;
  assign coh_req_link_o[104] = 1'b0;
  assign coh_req_link_o[105] = 1'b0;
  assign coh_req_link_o[106] = 1'b0;
  assign coh_req_link_o[107] = 1'b0;
  assign coh_req_link_o[108] = 1'b0;
  assign coh_req_link_o[109] = 1'b0;
  assign coh_req_link_o[110] = 1'b0;
  assign coh_req_link_o[111] = 1'b0;
  assign coh_req_link_o[112] = 1'b0;
  assign coh_req_link_o[113] = 1'b0;
  assign coh_req_link_o[114] = 1'b0;
  assign coh_req_link_o[115] = 1'b0;
  assign coh_req_link_o[116] = 1'b0;
  assign coh_req_link_o[117] = 1'b0;
  assign coh_req_link_o[118] = 1'b0;
  assign coh_req_link_o[119] = 1'b0;
  assign coh_req_link_o[120] = 1'b0;
  assign coh_req_link_o[121] = 1'b0;
  assign coh_req_link_o[122] = 1'b0;
  assign coh_req_link_o[123] = 1'b0;
  assign coh_req_link_o[124] = 1'b0;
  assign coh_req_link_o[125] = 1'b0;
  assign coh_req_link_o[126] = 1'b0;
  assign coh_req_link_o[127] = 1'b0;
  assign coh_req_link_o[128] = 1'b0;
  assign coh_req_link_o[129] = 1'b0;
  assign coh_req_link_o[130] = 1'b0;
  assign coh_req_link_o[131] = 1'b0;
  assign coh_req_link_o[132] = 1'b0;
  assign coh_req_link_o[133] = 1'b0;
  assign coh_req_link_o[134] = 1'b0;
  assign coh_req_link_o[135] = 1'b0;
  assign coh_req_link_o[136] = 1'b0;
  assign coh_req_link_o[137] = 1'b0;
  assign coh_req_link_o[138] = 1'b0;
  assign coh_req_link_o[139] = 1'b0;
  assign coh_req_link_o[140] = 1'b0;
  assign coh_req_link_o[141] = 1'b0;
  assign coh_req_link_o[142] = 1'b0;
  assign coh_req_link_o[143] = 1'b0;
  assign coh_req_link_o[144] = 1'b0;
  assign coh_req_link_o[145] = 1'b0;
  assign coh_req_link_o[146] = 1'b0;
  assign coh_req_link_o[147] = 1'b0;
  assign coh_req_link_o[148] = 1'b0;
  assign coh_req_link_o[149] = 1'b0;
  assign coh_req_link_o[150] = 1'b0;
  assign coh_req_link_o[151] = 1'b0;
  assign coh_req_link_o[152] = 1'b0;
  assign coh_req_link_o[153] = 1'b0;
  assign coh_req_link_o[154] = 1'b0;
  assign coh_req_link_o[155] = 1'b0;
  assign coh_req_link_o[156] = 1'b0;
  assign coh_req_link_o[157] = 1'b0;
  assign coh_req_link_o[158] = 1'b0;
  assign coh_req_link_o[159] = 1'b0;
  assign coh_req_link_o[160] = 1'b0;
  assign coh_req_link_o[161] = 1'b0;
  assign coh_req_link_o[162] = 1'b0;
  assign coh_req_link_o[163] = 1'b0;
  assign coh_req_link_o[164] = 1'b0;
  assign coh_req_link_o[165] = 1'b0;
  assign coh_req_link_o[166] = 1'b0;
  assign coh_req_link_o[167] = 1'b0;
  assign coh_req_link_o[168] = 1'b0;
  assign coh_req_link_o[169] = 1'b0;
  assign coh_req_link_o[170] = 1'b0;
  assign coh_req_link_o[171] = 1'b0;
  assign coh_req_link_o[172] = 1'b0;
  assign coh_req_link_o[173] = 1'b0;
  assign coh_req_link_o[174] = 1'b0;
  assign coh_req_link_o[175] = 1'b0;
  assign coh_req_link_o[176] = 1'b0;
  assign coh_req_link_o[177] = 1'b0;
  assign coh_req_link_o[178] = 1'b0;
  assign coh_req_link_o[179] = 1'b0;
  assign coh_req_link_o[180] = 1'b0;
  assign coh_req_link_o[181] = 1'b0;
  assign coh_req_link_o[182] = 1'b0;
  assign coh_req_link_o[183] = 1'b0;
  assign coh_req_link_o[184] = 1'b0;
  assign coh_req_link_o[185] = 1'b0;
  assign coh_req_link_o[186] = 1'b0;
  assign coh_req_link_o[187] = 1'b0;
  assign coh_req_link_o[188] = 1'b0;
  assign coh_req_link_o[189] = 1'b0;
  assign coh_req_link_o[190] = 1'b0;
  assign coh_req_link_o[191] = 1'b0;
  assign coh_req_link_o[192] = 1'b0;
  assign coh_req_link_o[193] = 1'b0;
  assign coh_req_link_o[194] = 1'b0;
  assign coh_req_link_o[195] = 1'b0;
  assign coh_req_link_o[196] = 1'b0;
  assign coh_req_link_o[197] = 1'b0;
  assign coh_req_link_o[198] = 1'b0;
  assign coh_req_link_o[199] = 1'b0;
  assign coh_req_link_o[200] = 1'b0;
  assign coh_req_link_o[201] = 1'b0;
  assign coh_req_link_o[202] = 1'b0;
  assign coh_req_link_o[203] = 1'b0;
  assign coh_req_link_o[204] = 1'b0;
  assign coh_req_link_o[205] = 1'b0;
  assign coh_req_link_o[206] = 1'b0;
  assign coh_req_link_o[207] = 1'b0;
  assign coh_req_link_o[208] = 1'b0;
  assign coh_req_link_o[209] = 1'b0;
  assign coh_req_link_o[210] = 1'b0;
  assign coh_req_link_o[211] = 1'b0;
  assign coh_req_link_o[212] = 1'b0;
  assign coh_req_link_o[213] = 1'b0;
  assign coh_req_link_o[214] = 1'b0;
  assign coh_req_link_o[215] = 1'b0;
  assign coh_req_link_o[216] = 1'b0;
  assign coh_req_link_o[217] = 1'b0;
  assign coh_req_link_o[218] = 1'b0;
  assign coh_req_link_o[219] = 1'b0;
  assign coh_req_link_o[220] = 1'b0;
  assign coh_req_link_o[221] = 1'b0;
  assign coh_req_link_o[222] = 1'b0;
  assign coh_req_link_o[223] = 1'b0;
  assign coh_req_link_o[224] = 1'b0;
  assign coh_req_link_o[225] = 1'b0;
  assign coh_req_link_o[226] = 1'b0;
  assign coh_req_link_o[227] = 1'b0;
  assign coh_req_link_o[228] = 1'b0;
  assign coh_req_link_o[229] = 1'b0;
  assign coh_req_link_o[230] = 1'b0;
  assign coh_req_link_o[231] = 1'b0;
  assign coh_req_link_o[232] = 1'b0;
  assign coh_req_link_o[233] = 1'b0;
  assign coh_req_link_o[234] = 1'b0;
  assign coh_req_link_o[235] = 1'b0;
  assign coh_req_link_o[236] = 1'b0;
  assign coh_req_link_o[237] = 1'b0;
  assign coh_req_link_o[238] = 1'b0;
  assign coh_req_link_o[239] = 1'b0;
  assign coh_req_link_o[240] = 1'b0;
  assign coh_req_link_o[241] = 1'b0;
  assign coh_req_link_o[242] = 1'b0;
  assign coh_req_link_o[243] = 1'b0;
  assign coh_req_link_o[244] = 1'b0;
  assign coh_req_link_o[245] = 1'b0;
  assign coh_req_link_o[246] = 1'b0;
  assign coh_req_link_o[247] = 1'b0;
  assign coh_req_link_o[248] = 1'b0;
  assign coh_req_link_o[249] = 1'b0;
  assign coh_req_link_o[250] = 1'b0;
  assign coh_req_link_o[251] = 1'b0;
  assign coh_req_link_o[252] = 1'b0;
  assign coh_req_link_o[253] = 1'b0;
  assign coh_req_link_o[254] = 1'b0;
  assign coh_req_link_o[255] = 1'b0;
  assign coh_req_link_o[256] = 1'b0;
  assign coh_req_link_o[257] = 1'b0;
  assign coh_req_link_o[258] = 1'b0;
  assign coh_req_link_o[259] = 1'b0;

endmodule