module tlb_00000010_00000001
(
  clk_i,
  rst_ni,
  flush_i,
  update_i,
  lu_access_i,
  lu_asid_i,
  lu_vaddr_i,
  lu_content_o,
  lu_is_2M_o,
  lu_is_1G_o,
  lu_hit_o
);

  input [94:0] update_i;
  input [0:0] lu_asid_i;
  input [63:0] lu_vaddr_i;
  output [63:0] lu_content_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input lu_access_i;
  output lu_is_2M_o;
  output lu_is_1G_o;
  output lu_hit_o;
  wire [63:0] lu_content_o;
  wire lu_is_2M_o,lu_is_1G_o,lu_hit_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,
  N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,
  N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,
  N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,
  N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,
  N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,
  N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,
  N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,
  N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,
  N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,
  N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,
  N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,
  N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,
  N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,
  N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,
  N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,
  N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,
  N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,
  N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,
  N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,
  N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,
  N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,
  N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,
  N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,
  N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,
  N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,
  N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,
  N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,
  N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,
  N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,
  N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,
  N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,
  N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,
  N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,
  N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,
  N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,
  N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,
  N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,
  N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,
  N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,
  N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,
  N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,
  N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,
  N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,
  N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,
  N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,
  N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,
  N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,
  N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,
  N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,
  N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,
  N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,
  N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,
  N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,
  N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,
  N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,
  N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,
  N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,
  N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,
  N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,
  N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,
  N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,
  N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,
  N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,
  N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,
  N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,
  N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,
  N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,
  N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,
  N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,
  N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
  N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,
  N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,
  N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,
  N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,
  N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,
  N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
  N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,
  N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,
  N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,
  N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,
  N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,
  N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,
  N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,
  N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,
  N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,
  N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,
  N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,
  N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,
  N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,
  N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,
  N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,
  N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,
  N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,
  N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,
  N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,
  N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,
  N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,
  N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,
  N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,
  N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,
  N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,
  N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,
  N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,
  N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,
  N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,
  N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,
  N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,
  N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,
  N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,
  N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,
  N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,
  N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,
  N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,
  N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,
  N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,
  N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,
  N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,
  N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,
  N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,
  N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,
  N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,
  N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,
  N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,
  N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,
  N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,
  N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
  N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,
  N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,
  N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
  N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,
  N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,
  N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
  N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,
  N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,
  N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
  N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,
  N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,
  N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
  N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,
  N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,
  N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
  N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,
  N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,
  N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
  N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,
  N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,
  N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
  N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,
  N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,
  N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
  N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,
  N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,
  N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
  N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,
  N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,
  N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
  N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,
  N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,
  N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
  N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,
  N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,
  N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
  N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,
  N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,
  N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
  N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,
  N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,
  N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
  N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,
  N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,
  N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
  N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,
  N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,
  N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
  N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,
  N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,
  N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
  N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,
  N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,
  N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
  N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,
  N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,
  N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
  N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,
  N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,
  N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
  N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,
  N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,
  N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
  N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,
  N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,
  N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
  N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,
  N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,
  N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
  N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,
  N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,
  N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
  N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,
  N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,
  N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
  N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,
  N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,
  N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
  N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,
  N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,
  N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
  N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,
  N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,
  N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
  N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,
  N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,
  N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
  N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,
  N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
  N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
  N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,
  N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,
  N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
  N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,
  N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,
  N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
  N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,
  N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,
  N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
  N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,
  N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,
  N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
  N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,
  N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,
  N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
  N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,
  N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,
  N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
  N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,
  N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,
  N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
  N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,
  N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,
  N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
  N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,
  N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,
  N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
  N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,
  N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,
  N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
  N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,
  N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,
  N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
  N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,
  N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,
  N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
  N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,
  N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,
  N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
  N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,
  N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,
  N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
  N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,
  N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,
  N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
  N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,
  N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,
  N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
  N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,
  N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,
  N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
  N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,
  N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,
  N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
  N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,
  N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,
  N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
  N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,
  N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,
  N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
  N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,
  N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,
  N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
  N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,
  N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,
  N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
  N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,
  N4553,tags_n_15__valid_,tags_n_14__valid_,tags_n_13__valid_,tags_n_12__valid_,
  tags_n_11__valid_,tags_n_10__valid_,tags_n_9__valid_,tags_n_8__valid_,
  tags_n_7__asid__0_,tags_n_7__vpn2__8_,tags_n_7__vpn2__7_,tags_n_7__vpn2__6_,
  tags_n_7__vpn2__5_,tags_n_7__vpn2__4_,tags_n_7__vpn2__3_,tags_n_7__vpn2__2_,tags_n_7__vpn2__1_,
  tags_n_7__vpn2__0_,tags_n_7__vpn1__8_,tags_n_7__vpn1__7_,tags_n_7__vpn1__6_,
  tags_n_7__vpn1__5_,tags_n_7__vpn1__4_,tags_n_7__vpn1__3_,tags_n_7__vpn1__2_,
  tags_n_7__vpn1__1_,tags_n_7__vpn1__0_,tags_n_7__vpn0__8_,tags_n_7__vpn0__7_,
  tags_n_7__vpn0__6_,tags_n_7__vpn0__5_,tags_n_7__vpn0__4_,tags_n_7__vpn0__3_,
  tags_n_7__vpn0__2_,tags_n_7__vpn0__1_,tags_n_7__vpn0__0_,tags_n_7__is_2M_,tags_n_7__is_1G_,
  tags_n_7__valid_,tags_n_6__asid__0_,tags_n_6__vpn2__8_,tags_n_6__vpn2__7_,
  tags_n_6__vpn2__6_,tags_n_6__vpn2__5_,tags_n_6__vpn2__4_,tags_n_6__vpn2__3_,
  tags_n_6__vpn2__2_,tags_n_6__vpn2__1_,tags_n_6__vpn2__0_,tags_n_6__vpn1__8_,tags_n_6__vpn1__7_,
  tags_n_6__vpn1__6_,tags_n_6__vpn1__5_,tags_n_6__vpn1__4_,tags_n_6__vpn1__3_,
  tags_n_6__vpn1__2_,tags_n_6__vpn1__1_,tags_n_6__vpn1__0_,tags_n_6__vpn0__8_,
  tags_n_6__vpn0__7_,tags_n_6__vpn0__6_,tags_n_6__vpn0__5_,tags_n_6__vpn0__4_,
  tags_n_6__vpn0__3_,tags_n_6__vpn0__2_,tags_n_6__vpn0__1_,tags_n_6__vpn0__0_,tags_n_6__is_2M_,
  tags_n_6__is_1G_,tags_n_6__valid_,tags_n_5__asid__0_,tags_n_5__vpn2__8_,
  tags_n_5__vpn2__7_,tags_n_5__vpn2__6_,tags_n_5__vpn2__5_,tags_n_5__vpn2__4_,
  tags_n_5__vpn2__3_,tags_n_5__vpn2__2_,tags_n_5__vpn2__1_,tags_n_5__vpn2__0_,
  tags_n_5__vpn1__8_,tags_n_5__vpn1__7_,tags_n_5__vpn1__6_,tags_n_5__vpn1__5_,tags_n_5__vpn1__4_,
  tags_n_5__vpn1__3_,tags_n_5__vpn1__2_,tags_n_5__vpn1__1_,tags_n_5__vpn1__0_,
  tags_n_5__vpn0__8_,tags_n_5__vpn0__7_,tags_n_5__vpn0__6_,tags_n_5__vpn0__5_,
  tags_n_5__vpn0__4_,tags_n_5__vpn0__3_,tags_n_5__vpn0__2_,tags_n_5__vpn0__1_,
  tags_n_5__vpn0__0_,tags_n_5__is_2M_,tags_n_5__is_1G_,tags_n_5__valid_,tags_n_4__asid__0_,
  tags_n_4__vpn2__8_,tags_n_4__vpn2__7_,tags_n_4__vpn2__6_,tags_n_4__vpn2__5_,
  tags_n_4__vpn2__4_,tags_n_4__vpn2__3_,tags_n_4__vpn2__2_,tags_n_4__vpn2__1_,
  tags_n_4__vpn2__0_,tags_n_4__vpn1__8_,tags_n_4__vpn1__7_,tags_n_4__vpn1__6_,
  tags_n_4__vpn1__5_,tags_n_4__vpn1__4_,tags_n_4__vpn1__3_,tags_n_4__vpn1__2_,tags_n_4__vpn1__1_,
  tags_n_4__vpn1__0_,tags_n_4__vpn0__8_,tags_n_4__vpn0__7_,tags_n_4__vpn0__6_,
  tags_n_4__vpn0__5_,tags_n_4__vpn0__4_,tags_n_4__vpn0__3_,tags_n_4__vpn0__2_,
  tags_n_4__vpn0__1_,tags_n_4__vpn0__0_,tags_n_4__is_2M_,tags_n_4__is_1G_,tags_n_4__valid_,
  tags_n_3__asid__0_,tags_n_3__vpn2__8_,tags_n_3__vpn2__7_,tags_n_3__vpn2__6_,
  tags_n_3__vpn2__5_,tags_n_3__vpn2__4_,tags_n_3__vpn2__3_,tags_n_3__vpn2__2_,
  tags_n_3__vpn2__1_,tags_n_3__vpn2__0_,tags_n_3__vpn1__8_,tags_n_3__vpn1__7_,
  tags_n_3__vpn1__6_,tags_n_3__vpn1__5_,tags_n_3__vpn1__4_,tags_n_3__vpn1__3_,
  tags_n_3__vpn1__2_,tags_n_3__vpn1__1_,tags_n_3__vpn1__0_,tags_n_3__vpn0__8_,tags_n_3__vpn0__7_,
  tags_n_3__vpn0__6_,tags_n_3__vpn0__5_,tags_n_3__vpn0__4_,tags_n_3__vpn0__3_,
  tags_n_3__vpn0__2_,tags_n_3__vpn0__1_,tags_n_3__vpn0__0_,tags_n_3__is_2M_,
  tags_n_3__is_1G_,tags_n_3__valid_,tags_n_2__asid__0_,tags_n_2__vpn2__8_,tags_n_2__vpn2__7_,
  tags_n_2__vpn2__6_,tags_n_2__vpn2__5_,tags_n_2__vpn2__4_,tags_n_2__vpn2__3_,
  tags_n_2__vpn2__2_,tags_n_2__vpn2__1_,tags_n_2__vpn2__0_,tags_n_2__vpn1__8_,
  tags_n_2__vpn1__7_,tags_n_2__vpn1__6_,tags_n_2__vpn1__5_,tags_n_2__vpn1__4_,
  tags_n_2__vpn1__3_,tags_n_2__vpn1__2_,tags_n_2__vpn1__1_,tags_n_2__vpn1__0_,
  tags_n_2__vpn0__8_,tags_n_2__vpn0__7_,tags_n_2__vpn0__6_,tags_n_2__vpn0__5_,tags_n_2__vpn0__4_,
  tags_n_2__vpn0__3_,tags_n_2__vpn0__2_,tags_n_2__vpn0__1_,tags_n_2__vpn0__0_,
  tags_n_2__is_2M_,tags_n_2__is_1G_,tags_n_2__valid_,tags_n_1__asid__0_,
  tags_n_1__vpn2__8_,tags_n_1__vpn2__7_,tags_n_1__vpn2__6_,tags_n_1__vpn2__5_,tags_n_1__vpn2__4_,
  tags_n_1__vpn2__3_,tags_n_1__vpn2__2_,tags_n_1__vpn2__1_,tags_n_1__vpn2__0_,
  tags_n_1__vpn1__8_,tags_n_1__vpn1__7_,tags_n_1__vpn1__6_,tags_n_1__vpn1__5_,
  tags_n_1__vpn1__4_,tags_n_1__vpn1__3_,tags_n_1__vpn1__2_,tags_n_1__vpn1__1_,
  tags_n_1__vpn1__0_,tags_n_1__vpn0__8_,tags_n_1__vpn0__7_,tags_n_1__vpn0__6_,
  tags_n_1__vpn0__5_,tags_n_1__vpn0__4_,tags_n_1__vpn0__3_,tags_n_1__vpn0__2_,tags_n_1__vpn0__1_,
  tags_n_1__vpn0__0_,tags_n_1__is_2M_,tags_n_1__is_1G_,tags_n_1__valid_,
  tags_n_0__asid__0_,tags_n_0__vpn2__8_,tags_n_0__vpn2__7_,tags_n_0__vpn2__6_,
  tags_n_0__vpn2__5_,tags_n_0__vpn2__4_,tags_n_0__vpn2__3_,tags_n_0__vpn2__2_,tags_n_0__vpn2__1_,
  tags_n_0__vpn2__0_,tags_n_0__vpn1__8_,tags_n_0__vpn1__7_,tags_n_0__vpn1__6_,
  tags_n_0__vpn1__5_,tags_n_0__vpn1__4_,tags_n_0__vpn1__3_,tags_n_0__vpn1__2_,
  tags_n_0__vpn1__1_,tags_n_0__vpn1__0_,tags_n_0__vpn0__8_,tags_n_0__vpn0__7_,
  tags_n_0__vpn0__6_,tags_n_0__vpn0__5_,tags_n_0__vpn0__4_,tags_n_0__vpn0__3_,
  tags_n_0__vpn0__2_,tags_n_0__vpn0__1_,tags_n_0__vpn0__0_,tags_n_0__is_2M_,tags_n_0__is_1G_,
  tags_n_0__valid_,content_n_7__reserved__9_,content_n_7__reserved__8_,
  content_n_7__reserved__7_,content_n_7__reserved__6_,content_n_7__reserved__5_,
  content_n_7__reserved__4_,content_n_7__reserved__3_,content_n_7__reserved__2_,
  content_n_7__reserved__1_,content_n_7__reserved__0_,content_n_7__ppn__43_,content_n_7__ppn__42_,
  content_n_7__ppn__41_,content_n_7__ppn__40_,content_n_7__ppn__39_,
  content_n_7__ppn__38_,content_n_7__ppn__37_,content_n_7__ppn__36_,content_n_7__ppn__35_,
  content_n_7__ppn__34_,content_n_7__ppn__33_,content_n_7__ppn__32_,content_n_7__ppn__31_,
  content_n_7__ppn__30_,content_n_7__ppn__29_,content_n_7__ppn__28_,
  content_n_7__ppn__27_,content_n_7__ppn__26_,content_n_7__ppn__25_,content_n_7__ppn__24_,
  content_n_7__ppn__23_,content_n_7__ppn__22_,content_n_7__ppn__21_,content_n_7__ppn__20_,
  content_n_7__ppn__19_,content_n_7__ppn__18_,content_n_7__ppn__17_,
  content_n_7__ppn__16_,content_n_7__ppn__15_,content_n_7__ppn__14_,content_n_7__ppn__13_,
  content_n_7__ppn__12_,content_n_7__ppn__11_,content_n_7__ppn__10_,content_n_7__ppn__9_,
  content_n_7__ppn__8_,content_n_7__ppn__7_,content_n_7__ppn__6_,
  content_n_7__ppn__5_,content_n_7__ppn__4_,content_n_7__ppn__3_,content_n_7__ppn__2_,
  content_n_7__ppn__1_,content_n_7__ppn__0_,content_n_7__rsw__1_,content_n_7__rsw__0_,
  content_n_7__d_,content_n_7__a_,content_n_7__g_,content_n_7__u_,content_n_7__x_,
  content_n_7__w_,content_n_7__r_,content_n_7__v_,content_n_6__reserved__9_,
  content_n_6__reserved__8_,content_n_6__reserved__7_,content_n_6__reserved__6_,
  content_n_6__reserved__5_,content_n_6__reserved__4_,content_n_6__reserved__3_,
  content_n_6__reserved__2_,content_n_6__reserved__1_,content_n_6__reserved__0_,
  content_n_6__ppn__43_,content_n_6__ppn__42_,content_n_6__ppn__41_,content_n_6__ppn__40_,
  content_n_6__ppn__39_,content_n_6__ppn__38_,content_n_6__ppn__37_,content_n_6__ppn__36_,
  content_n_6__ppn__35_,content_n_6__ppn__34_,content_n_6__ppn__33_,
  content_n_6__ppn__32_,content_n_6__ppn__31_,content_n_6__ppn__30_,content_n_6__ppn__29_,
  content_n_6__ppn__28_,content_n_6__ppn__27_,content_n_6__ppn__26_,content_n_6__ppn__25_,
  content_n_6__ppn__24_,content_n_6__ppn__23_,content_n_6__ppn__22_,
  content_n_6__ppn__21_,content_n_6__ppn__20_,content_n_6__ppn__19_,content_n_6__ppn__18_,
  content_n_6__ppn__17_,content_n_6__ppn__16_,content_n_6__ppn__15_,content_n_6__ppn__14_,
  content_n_6__ppn__13_,content_n_6__ppn__12_,content_n_6__ppn__11_,
  content_n_6__ppn__10_,content_n_6__ppn__9_,content_n_6__ppn__8_,content_n_6__ppn__7_,
  content_n_6__ppn__6_,content_n_6__ppn__5_,content_n_6__ppn__4_,content_n_6__ppn__3_,
  content_n_6__ppn__2_,content_n_6__ppn__1_,content_n_6__ppn__0_,content_n_6__rsw__1_,
  content_n_6__rsw__0_,content_n_6__d_,content_n_6__a_,content_n_6__g_,
  content_n_6__u_,content_n_6__x_,content_n_6__w_,content_n_6__r_,content_n_6__v_,
  content_n_5__reserved__9_,content_n_5__reserved__8_,content_n_5__reserved__7_,
  content_n_5__reserved__6_,content_n_5__reserved__5_,content_n_5__reserved__4_,
  content_n_5__reserved__3_,content_n_5__reserved__2_,content_n_5__reserved__1_,
  content_n_5__reserved__0_,content_n_5__ppn__43_,content_n_5__ppn__42_,content_n_5__ppn__41_,
  content_n_5__ppn__40_,content_n_5__ppn__39_,content_n_5__ppn__38_,
  content_n_5__ppn__37_,content_n_5__ppn__36_,content_n_5__ppn__35_,content_n_5__ppn__34_,
  content_n_5__ppn__33_,content_n_5__ppn__32_,content_n_5__ppn__31_,content_n_5__ppn__30_,
  content_n_5__ppn__29_,content_n_5__ppn__28_,content_n_5__ppn__27_,
  content_n_5__ppn__26_,content_n_5__ppn__25_,content_n_5__ppn__24_,content_n_5__ppn__23_,
  content_n_5__ppn__22_,content_n_5__ppn__21_,content_n_5__ppn__20_,content_n_5__ppn__19_,
  content_n_5__ppn__18_,content_n_5__ppn__17_,content_n_5__ppn__16_,
  content_n_5__ppn__15_,content_n_5__ppn__14_,content_n_5__ppn__13_,content_n_5__ppn__12_,
  content_n_5__ppn__11_,content_n_5__ppn__10_,content_n_5__ppn__9_,content_n_5__ppn__8_,
  content_n_5__ppn__7_,content_n_5__ppn__6_,content_n_5__ppn__5_,
  content_n_5__ppn__4_,content_n_5__ppn__3_,content_n_5__ppn__2_,content_n_5__ppn__1_,
  content_n_5__ppn__0_,content_n_5__rsw__1_,content_n_5__rsw__0_,content_n_5__d_,content_n_5__a_,
  content_n_5__g_,content_n_5__u_,content_n_5__x_,content_n_5__w_,content_n_5__r_,
  content_n_5__v_,content_n_4__reserved__9_,content_n_4__reserved__8_,
  content_n_4__reserved__7_,content_n_4__reserved__6_,content_n_4__reserved__5_,
  content_n_4__reserved__4_,content_n_4__reserved__3_,content_n_4__reserved__2_,
  content_n_4__reserved__1_,content_n_4__reserved__0_,content_n_4__ppn__43_,content_n_4__ppn__42_,
  content_n_4__ppn__41_,content_n_4__ppn__40_,content_n_4__ppn__39_,
  content_n_4__ppn__38_,content_n_4__ppn__37_,content_n_4__ppn__36_,content_n_4__ppn__35_,
  content_n_4__ppn__34_,content_n_4__ppn__33_,content_n_4__ppn__32_,
  content_n_4__ppn__31_,content_n_4__ppn__30_,content_n_4__ppn__29_,content_n_4__ppn__28_,
  content_n_4__ppn__27_,content_n_4__ppn__26_,content_n_4__ppn__25_,content_n_4__ppn__24_,
  content_n_4__ppn__23_,content_n_4__ppn__22_,content_n_4__ppn__21_,
  content_n_4__ppn__20_,content_n_4__ppn__19_,content_n_4__ppn__18_,content_n_4__ppn__17_,
  content_n_4__ppn__16_,content_n_4__ppn__15_,content_n_4__ppn__14_,content_n_4__ppn__13_,
  content_n_4__ppn__12_,content_n_4__ppn__11_,content_n_4__ppn__10_,
  content_n_4__ppn__9_,content_n_4__ppn__8_,content_n_4__ppn__7_,content_n_4__ppn__6_,
  content_n_4__ppn__5_,content_n_4__ppn__4_,content_n_4__ppn__3_,content_n_4__ppn__2_,
  content_n_4__ppn__1_,content_n_4__ppn__0_,content_n_4__rsw__1_,content_n_4__rsw__0_,
  content_n_4__d_,content_n_4__a_,content_n_4__g_,content_n_4__u_,content_n_4__x_,
  content_n_4__w_,content_n_4__r_,content_n_4__v_,content_n_3__reserved__9_,
  content_n_3__reserved__8_,content_n_3__reserved__7_,content_n_3__reserved__6_,
  content_n_3__reserved__5_,content_n_3__reserved__4_,content_n_3__reserved__3_,
  content_n_3__reserved__2_,content_n_3__reserved__1_,content_n_3__reserved__0_,
  content_n_3__ppn__43_,content_n_3__ppn__42_,content_n_3__ppn__41_,content_n_3__ppn__40_,
  content_n_3__ppn__39_,content_n_3__ppn__38_,content_n_3__ppn__37_,content_n_3__ppn__36_,
  content_n_3__ppn__35_,content_n_3__ppn__34_,content_n_3__ppn__33_,
  content_n_3__ppn__32_,content_n_3__ppn__31_,content_n_3__ppn__30_,content_n_3__ppn__29_,
  content_n_3__ppn__28_,content_n_3__ppn__27_,content_n_3__ppn__26_,
  content_n_3__ppn__25_,content_n_3__ppn__24_,content_n_3__ppn__23_,content_n_3__ppn__22_,
  content_n_3__ppn__21_,content_n_3__ppn__20_,content_n_3__ppn__19_,content_n_3__ppn__18_,
  content_n_3__ppn__17_,content_n_3__ppn__16_,content_n_3__ppn__15_,
  content_n_3__ppn__14_,content_n_3__ppn__13_,content_n_3__ppn__12_,content_n_3__ppn__11_,
  content_n_3__ppn__10_,content_n_3__ppn__9_,content_n_3__ppn__8_,content_n_3__ppn__7_,
  content_n_3__ppn__6_,content_n_3__ppn__5_,content_n_3__ppn__4_,content_n_3__ppn__3_,
  content_n_3__ppn__2_,content_n_3__ppn__1_,content_n_3__ppn__0_,
  content_n_3__rsw__1_,content_n_3__rsw__0_,content_n_3__d_,content_n_3__a_,content_n_3__g_,
  content_n_3__u_,content_n_3__x_,content_n_3__w_,content_n_3__r_,content_n_3__v_,
  content_n_2__reserved__9_,content_n_2__reserved__8_,content_n_2__reserved__7_,
  content_n_2__reserved__6_,content_n_2__reserved__5_,content_n_2__reserved__4_,
  content_n_2__reserved__3_,content_n_2__reserved__2_,content_n_2__reserved__1_,
  content_n_2__reserved__0_,content_n_2__ppn__43_,content_n_2__ppn__42_,content_n_2__ppn__41_,
  content_n_2__ppn__40_,content_n_2__ppn__39_,content_n_2__ppn__38_,
  content_n_2__ppn__37_,content_n_2__ppn__36_,content_n_2__ppn__35_,content_n_2__ppn__34_,
  content_n_2__ppn__33_,content_n_2__ppn__32_,content_n_2__ppn__31_,content_n_2__ppn__30_,
  content_n_2__ppn__29_,content_n_2__ppn__28_,content_n_2__ppn__27_,
  content_n_2__ppn__26_,content_n_2__ppn__25_,content_n_2__ppn__24_,content_n_2__ppn__23_,
  content_n_2__ppn__22_,content_n_2__ppn__21_,content_n_2__ppn__20_,
  content_n_2__ppn__19_,content_n_2__ppn__18_,content_n_2__ppn__17_,content_n_2__ppn__16_,
  content_n_2__ppn__15_,content_n_2__ppn__14_,content_n_2__ppn__13_,content_n_2__ppn__12_,
  content_n_2__ppn__11_,content_n_2__ppn__10_,content_n_2__ppn__9_,
  content_n_2__ppn__8_,content_n_2__ppn__7_,content_n_2__ppn__6_,content_n_2__ppn__5_,
  content_n_2__ppn__4_,content_n_2__ppn__3_,content_n_2__ppn__2_,content_n_2__ppn__1_,
  content_n_2__ppn__0_,content_n_2__rsw__1_,content_n_2__rsw__0_,content_n_2__d_,
  content_n_2__a_,content_n_2__g_,content_n_2__u_,content_n_2__x_,content_n_2__w_,
  content_n_2__r_,content_n_2__v_,content_n_1__reserved__9_,content_n_1__reserved__8_,
  content_n_1__reserved__7_,content_n_1__reserved__6_,content_n_1__reserved__5_,
  content_n_1__reserved__4_,content_n_1__reserved__3_,content_n_1__reserved__2_,
  content_n_1__reserved__1_,content_n_1__reserved__0_,content_n_1__ppn__43_,
  content_n_1__ppn__42_,content_n_1__ppn__41_,content_n_1__ppn__40_,content_n_1__ppn__39_,
  content_n_1__ppn__38_,content_n_1__ppn__37_,content_n_1__ppn__36_,content_n_1__ppn__35_,
  content_n_1__ppn__34_,content_n_1__ppn__33_,content_n_1__ppn__32_,
  content_n_1__ppn__31_,content_n_1__ppn__30_,content_n_1__ppn__29_,content_n_1__ppn__28_,
  content_n_1__ppn__27_,content_n_1__ppn__26_,content_n_1__ppn__25_,content_n_1__ppn__24_,
  content_n_1__ppn__23_,content_n_1__ppn__22_,content_n_1__ppn__21_,
  content_n_1__ppn__20_,content_n_1__ppn__19_,content_n_1__ppn__18_,content_n_1__ppn__17_,
  content_n_1__ppn__16_,content_n_1__ppn__15_,content_n_1__ppn__14_,
  content_n_1__ppn__13_,content_n_1__ppn__12_,content_n_1__ppn__11_,content_n_1__ppn__10_,
  content_n_1__ppn__9_,content_n_1__ppn__8_,content_n_1__ppn__7_,content_n_1__ppn__6_,
  content_n_1__ppn__5_,content_n_1__ppn__4_,content_n_1__ppn__3_,content_n_1__ppn__2_,
  content_n_1__ppn__1_,content_n_1__ppn__0_,content_n_1__rsw__1_,content_n_1__rsw__0_,
  content_n_1__d_,content_n_1__a_,content_n_1__g_,content_n_1__u_,content_n_1__x_,
  content_n_1__w_,content_n_1__r_,content_n_1__v_,content_n_0__reserved__9_,
  content_n_0__reserved__8_,content_n_0__reserved__7_,content_n_0__reserved__6_,
  content_n_0__reserved__5_,content_n_0__reserved__4_,content_n_0__reserved__3_,
  content_n_0__reserved__2_,content_n_0__reserved__1_,content_n_0__reserved__0_,
  content_n_0__ppn__43_,content_n_0__ppn__42_,content_n_0__ppn__41_,content_n_0__ppn__40_,
  content_n_0__ppn__39_,content_n_0__ppn__38_,content_n_0__ppn__37_,
  content_n_0__ppn__36_,content_n_0__ppn__35_,content_n_0__ppn__34_,content_n_0__ppn__33_,
  content_n_0__ppn__32_,content_n_0__ppn__31_,content_n_0__ppn__30_,content_n_0__ppn__29_,
  content_n_0__ppn__28_,content_n_0__ppn__27_,content_n_0__ppn__26_,
  content_n_0__ppn__25_,content_n_0__ppn__24_,content_n_0__ppn__23_,content_n_0__ppn__22_,
  content_n_0__ppn__21_,content_n_0__ppn__20_,content_n_0__ppn__19_,content_n_0__ppn__18_,
  content_n_0__ppn__17_,content_n_0__ppn__16_,content_n_0__ppn__15_,
  content_n_0__ppn__14_,content_n_0__ppn__13_,content_n_0__ppn__12_,content_n_0__ppn__11_,
  content_n_0__ppn__10_,content_n_0__ppn__9_,content_n_0__ppn__8_,content_n_0__ppn__7_,
  content_n_0__ppn__6_,content_n_0__ppn__5_,content_n_0__ppn__4_,
  content_n_0__ppn__3_,content_n_0__ppn__2_,content_n_0__ppn__1_,content_n_0__ppn__0_,
  content_n_0__rsw__1_,content_n_0__rsw__0_,content_n_0__d_,content_n_0__a_,content_n_0__g_,
  content_n_0__u_,content_n_0__x_,content_n_0__w_,content_n_0__r_,content_n_0__v_,
  N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,
  N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,
  N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,
  N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,
  N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,
  N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,
  N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,
  N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,
  N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,
  N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,
  N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,
  N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,
  N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,
  N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,
  N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,
  N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,
  N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,
  N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,
  N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,
  N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,
  N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,
  N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,
  N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,
  N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868;
  wire [15:0] lu_hit,replace_en;
  wire [14:0] plru_tree_n;
  reg [14:0] plru_tree_q;
  reg [495:0] tags_q;
  reg [1023:0] content_q;
  assign N0 = lu_asid_i[0] ^ tags_q[30];
  assign N145 = ~N0;
  assign N146 = lu_vaddr_i[38:30] == tags_q[29:21];
  assign N152 = lu_vaddr_i[29:21] == tags_q[20:12];
  assign N154 = lu_vaddr_i[20:12] == tags_q[11:3];
  assign N1 = lu_asid_i[0] ^ tags_q[61];
  assign N421 = ~N1;
  assign N422 = lu_vaddr_i[38:30] == tags_q[60:52];
  assign N428 = lu_vaddr_i[29:21] == tags_q[51:43];
  assign N430 = lu_vaddr_i[20:12] == tags_q[42:34];
  assign N2 = lu_asid_i[0] ^ tags_q[92];
  assign N701 = ~N2;
  assign N702 = lu_vaddr_i[38:30] == tags_q[91:83];
  assign N708 = lu_vaddr_i[29:21] == tags_q[82:74];
  assign N710 = lu_vaddr_i[20:12] == tags_q[73:65];
  assign N3 = lu_asid_i[0] ^ tags_q[123];
  assign N981 = ~N3;
  assign N982 = lu_vaddr_i[38:30] == tags_q[122:114];
  assign N988 = lu_vaddr_i[29:21] == tags_q[113:105];
  assign N990 = lu_vaddr_i[20:12] == tags_q[104:96];
  assign N4 = lu_asid_i[0] ^ tags_q[154];
  assign N1261 = ~N4;
  assign N1262 = lu_vaddr_i[38:30] == tags_q[153:145];
  assign N1268 = lu_vaddr_i[29:21] == tags_q[144:136];
  assign N1270 = lu_vaddr_i[20:12] == tags_q[135:127];
  assign N5 = lu_asid_i[0] ^ tags_q[185];
  assign N1541 = ~N5;
  assign N1542 = lu_vaddr_i[38:30] == tags_q[184:176];
  assign N1548 = lu_vaddr_i[29:21] == tags_q[175:167];
  assign N1550 = lu_vaddr_i[20:12] == tags_q[166:158];
  assign N6 = lu_asid_i[0] ^ tags_q[216];
  assign N1821 = ~N6;
  assign N1822 = lu_vaddr_i[38:30] == tags_q[215:207];
  assign N1828 = lu_vaddr_i[29:21] == tags_q[206:198];
  assign N1830 = lu_vaddr_i[20:12] == tags_q[197:189];
  assign N7 = lu_asid_i[0] ^ tags_q[247];
  assign N2101 = ~N7;
  assign N2102 = lu_vaddr_i[38:30] == tags_q[246:238];
  assign N2108 = lu_vaddr_i[29:21] == tags_q[237:229];
  assign N2110 = lu_vaddr_i[20:12] == tags_q[228:220];
  assign N8 = lu_asid_i[0] ^ tags_q[278];
  assign N2381 = ~N8;
  assign N2382 = lu_vaddr_i[38:30] == tags_q[277:269];
  assign N2388 = lu_vaddr_i[29:21] == tags_q[268:260];
  assign N2390 = lu_vaddr_i[20:12] == tags_q[259:251];
  assign N9 = lu_asid_i[0] ^ tags_q[309];
  assign N2661 = ~N9;
  assign N2662 = lu_vaddr_i[38:30] == tags_q[308:300];
  assign N2668 = lu_vaddr_i[29:21] == tags_q[299:291];
  assign N2670 = lu_vaddr_i[20:12] == tags_q[290:282];
  assign N10 = lu_asid_i[0] ^ tags_q[340];
  assign N2941 = ~N10;
  assign N2942 = lu_vaddr_i[38:30] == tags_q[339:331];
  assign N2948 = lu_vaddr_i[29:21] == tags_q[330:322];
  assign N2950 = lu_vaddr_i[20:12] == tags_q[321:313];
  assign N11 = lu_asid_i[0] ^ tags_q[371];
  assign N3221 = ~N11;
  assign N3222 = lu_vaddr_i[38:30] == tags_q[370:362];
  assign N3228 = lu_vaddr_i[29:21] == tags_q[361:353];
  assign N3230 = lu_vaddr_i[20:12] == tags_q[352:344];
  assign N12 = lu_asid_i[0] ^ tags_q[402];
  assign N3501 = ~N12;
  assign N3502 = lu_vaddr_i[38:30] == tags_q[401:393];
  assign N3508 = lu_vaddr_i[29:21] == tags_q[392:384];
  assign N3510 = lu_vaddr_i[20:12] == tags_q[383:375];
  assign N13 = lu_asid_i[0] ^ tags_q[433];
  assign N3781 = ~N13;
  assign N3782 = lu_vaddr_i[38:30] == tags_q[432:424];
  assign N3788 = lu_vaddr_i[29:21] == tags_q[423:415];
  assign N3790 = lu_vaddr_i[20:12] == tags_q[414:406];
  assign N14 = lu_asid_i[0] ^ tags_q[464];
  assign N4061 = ~N14;
  assign N4062 = lu_vaddr_i[38:30] == tags_q[463:455];
  assign N4068 = lu_vaddr_i[29:21] == tags_q[454:446];
  assign N4070 = lu_vaddr_i[20:12] == tags_q[445:437];
  assign N15 = lu_asid_i[0] ^ tags_q[495];
  assign N4341 = ~N15;
  assign N4342 = lu_vaddr_i[38:30] == tags_q[494:486];
  assign N4348 = lu_vaddr_i[29:21] == tags_q[485:477];
  assign N4350 = lu_vaddr_i[20:12] == tags_q[476:468];
  assign N16 = lu_asid_i[0] ^ tags_q[30];
  assign N4557 = ~N16;
  assign N17 = lu_asid_i[0] ^ tags_q[61];
  assign N4563 = ~N17;
  assign N18 = lu_asid_i[0] ^ tags_q[92];
  assign N4569 = ~N18;
  assign N19 = lu_asid_i[0] ^ tags_q[123];
  assign N4575 = ~N19;
  assign N20 = lu_asid_i[0] ^ tags_q[154];
  assign N4581 = ~N20;
  assign N21 = lu_asid_i[0] ^ tags_q[185];
  assign N4587 = ~N21;
  assign N22 = lu_asid_i[0] ^ tags_q[216];
  assign N4593 = ~N22;
  assign N23 = lu_asid_i[0] ^ tags_q[247];
  assign N4599 = ~N23;
  assign N24 = lu_asid_i[0] ^ tags_q[278];
  assign N4605 = ~N24;
  assign N25 = lu_asid_i[0] ^ tags_q[309];
  assign N4611 = ~N25;
  assign N26 = lu_asid_i[0] ^ tags_q[340];
  assign N4617 = ~N26;
  assign N27 = lu_asid_i[0] ^ tags_q[371];
  assign N4623 = ~N27;
  assign N28 = lu_asid_i[0] ^ tags_q[402];
  assign N4629 = ~N28;
  assign N29 = lu_asid_i[0] ^ tags_q[433];
  assign N4635 = ~N29;
  assign N30 = lu_asid_i[0] ^ tags_q[464];
  assign N4641 = ~N30;
  assign N31 = lu_asid_i[0] ^ tags_q[495];
  assign N4647 = ~N31;

  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[14] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[14] <= plru_tree_n[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[13] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[13] <= plru_tree_n[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[12] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[12] <= plru_tree_n[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[11] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[11] <= plru_tree_n[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[10] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[10] <= plru_tree_n[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[9] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[9] <= plru_tree_n[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[8] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[8] <= plru_tree_n[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[7] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[7] <= plru_tree_n[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[6] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[6] <= plru_tree_n[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[5] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[5] <= plru_tree_n[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[4] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[4] <= plru_tree_n[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[3] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[3] <= plru_tree_n[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[2] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[2] <= plru_tree_n[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[1] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[1] <= plru_tree_n[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      plru_tree_q[0] <= 1'b0;
    end else if(1'b1) begin
      plru_tree_q[0] <= plru_tree_n[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[495] <= 1'b0;
    end else if(N4783) begin
      tags_q[495] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[494] <= 1'b0;
    end else if(N4783) begin
      tags_q[494] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[493] <= 1'b0;
    end else if(N4783) begin
      tags_q[493] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[492] <= 1'b0;
    end else if(N4783) begin
      tags_q[492] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[491] <= 1'b0;
    end else if(N4783) begin
      tags_q[491] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[490] <= 1'b0;
    end else if(N4783) begin
      tags_q[490] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[489] <= 1'b0;
    end else if(N4783) begin
      tags_q[489] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[488] <= 1'b0;
    end else if(N4783) begin
      tags_q[488] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[487] <= 1'b0;
    end else if(N4783) begin
      tags_q[487] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[486] <= 1'b0;
    end else if(N4783) begin
      tags_q[486] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[485] <= 1'b0;
    end else if(N4783) begin
      tags_q[485] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[484] <= 1'b0;
    end else if(N4783) begin
      tags_q[484] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[483] <= 1'b0;
    end else if(N4783) begin
      tags_q[483] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[482] <= 1'b0;
    end else if(N4783) begin
      tags_q[482] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[481] <= 1'b0;
    end else if(N4783) begin
      tags_q[481] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[480] <= 1'b0;
    end else if(N4783) begin
      tags_q[480] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[479] <= 1'b0;
    end else if(N4783) begin
      tags_q[479] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[478] <= 1'b0;
    end else if(N4783) begin
      tags_q[478] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[477] <= 1'b0;
    end else if(N4783) begin
      tags_q[477] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[476] <= 1'b0;
    end else if(N4783) begin
      tags_q[476] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[475] <= 1'b0;
    end else if(N4783) begin
      tags_q[475] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[474] <= 1'b0;
    end else if(N4783) begin
      tags_q[474] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[473] <= 1'b0;
    end else if(N4783) begin
      tags_q[473] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[472] <= 1'b0;
    end else if(N4783) begin
      tags_q[472] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[471] <= 1'b0;
    end else if(N4783) begin
      tags_q[471] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[470] <= 1'b0;
    end else if(N4783) begin
      tags_q[470] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[469] <= 1'b0;
    end else if(N4783) begin
      tags_q[469] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[468] <= 1'b0;
    end else if(N4783) begin
      tags_q[468] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[467] <= 1'b0;
    end else if(N4783) begin
      tags_q[467] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[466] <= 1'b0;
    end else if(N4783) begin
      tags_q[466] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[465] <= 1'b0;
    end else if(N4786) begin
      tags_q[465] <= tags_n_15__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[464] <= 1'b0;
    end else if(N4788) begin
      tags_q[464] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[463] <= 1'b0;
    end else if(N4788) begin
      tags_q[463] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[462] <= 1'b0;
    end else if(N4788) begin
      tags_q[462] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[461] <= 1'b0;
    end else if(N4788) begin
      tags_q[461] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[460] <= 1'b0;
    end else if(N4788) begin
      tags_q[460] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[459] <= 1'b0;
    end else if(N4788) begin
      tags_q[459] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[458] <= 1'b0;
    end else if(N4788) begin
      tags_q[458] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[457] <= 1'b0;
    end else if(N4788) begin
      tags_q[457] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[456] <= 1'b0;
    end else if(N4788) begin
      tags_q[456] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[455] <= 1'b0;
    end else if(N4788) begin
      tags_q[455] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[454] <= 1'b0;
    end else if(N4788) begin
      tags_q[454] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[453] <= 1'b0;
    end else if(N4788) begin
      tags_q[453] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[452] <= 1'b0;
    end else if(N4788) begin
      tags_q[452] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[451] <= 1'b0;
    end else if(N4788) begin
      tags_q[451] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[450] <= 1'b0;
    end else if(N4788) begin
      tags_q[450] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[449] <= 1'b0;
    end else if(N4788) begin
      tags_q[449] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[448] <= 1'b0;
    end else if(N4788) begin
      tags_q[448] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[447] <= 1'b0;
    end else if(N4788) begin
      tags_q[447] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[446] <= 1'b0;
    end else if(N4788) begin
      tags_q[446] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[445] <= 1'b0;
    end else if(N4788) begin
      tags_q[445] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[444] <= 1'b0;
    end else if(N4788) begin
      tags_q[444] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[443] <= 1'b0;
    end else if(N4788) begin
      tags_q[443] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[442] <= 1'b0;
    end else if(N4788) begin
      tags_q[442] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[441] <= 1'b0;
    end else if(N4788) begin
      tags_q[441] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[440] <= 1'b0;
    end else if(N4788) begin
      tags_q[440] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[439] <= 1'b0;
    end else if(N4788) begin
      tags_q[439] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[438] <= 1'b0;
    end else if(N4788) begin
      tags_q[438] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[437] <= 1'b0;
    end else if(N4788) begin
      tags_q[437] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[436] <= 1'b0;
    end else if(N4788) begin
      tags_q[436] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[435] <= 1'b0;
    end else if(N4788) begin
      tags_q[435] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[434] <= 1'b0;
    end else if(N4791) begin
      tags_q[434] <= tags_n_14__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[433] <= 1'b0;
    end else if(N4793) begin
      tags_q[433] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[432] <= 1'b0;
    end else if(N4793) begin
      tags_q[432] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[431] <= 1'b0;
    end else if(N4793) begin
      tags_q[431] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[430] <= 1'b0;
    end else if(N4793) begin
      tags_q[430] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[429] <= 1'b0;
    end else if(N4793) begin
      tags_q[429] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[428] <= 1'b0;
    end else if(N4793) begin
      tags_q[428] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[427] <= 1'b0;
    end else if(N4793) begin
      tags_q[427] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[426] <= 1'b0;
    end else if(N4793) begin
      tags_q[426] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[425] <= 1'b0;
    end else if(N4793) begin
      tags_q[425] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[424] <= 1'b0;
    end else if(N4793) begin
      tags_q[424] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[423] <= 1'b0;
    end else if(N4793) begin
      tags_q[423] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[422] <= 1'b0;
    end else if(N4793) begin
      tags_q[422] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[421] <= 1'b0;
    end else if(N4793) begin
      tags_q[421] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[420] <= 1'b0;
    end else if(N4793) begin
      tags_q[420] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[419] <= 1'b0;
    end else if(N4793) begin
      tags_q[419] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[418] <= 1'b0;
    end else if(N4793) begin
      tags_q[418] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[417] <= 1'b0;
    end else if(N4793) begin
      tags_q[417] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[416] <= 1'b0;
    end else if(N4793) begin
      tags_q[416] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[415] <= 1'b0;
    end else if(N4793) begin
      tags_q[415] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[414] <= 1'b0;
    end else if(N4793) begin
      tags_q[414] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[413] <= 1'b0;
    end else if(N4793) begin
      tags_q[413] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[412] <= 1'b0;
    end else if(N4793) begin
      tags_q[412] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[411] <= 1'b0;
    end else if(N4793) begin
      tags_q[411] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[410] <= 1'b0;
    end else if(N4793) begin
      tags_q[410] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[409] <= 1'b0;
    end else if(N4793) begin
      tags_q[409] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[408] <= 1'b0;
    end else if(N4793) begin
      tags_q[408] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[407] <= 1'b0;
    end else if(N4793) begin
      tags_q[407] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[406] <= 1'b0;
    end else if(N4793) begin
      tags_q[406] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[405] <= 1'b0;
    end else if(N4793) begin
      tags_q[405] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[404] <= 1'b0;
    end else if(N4793) begin
      tags_q[404] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[403] <= 1'b0;
    end else if(N4796) begin
      tags_q[403] <= tags_n_13__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[402] <= 1'b0;
    end else if(N4798) begin
      tags_q[402] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[401] <= 1'b0;
    end else if(N4798) begin
      tags_q[401] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[400] <= 1'b0;
    end else if(N4798) begin
      tags_q[400] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[399] <= 1'b0;
    end else if(N4798) begin
      tags_q[399] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[398] <= 1'b0;
    end else if(N4798) begin
      tags_q[398] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[397] <= 1'b0;
    end else if(N4798) begin
      tags_q[397] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[396] <= 1'b0;
    end else if(N4798) begin
      tags_q[396] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[395] <= 1'b0;
    end else if(N4798) begin
      tags_q[395] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[394] <= 1'b0;
    end else if(N4798) begin
      tags_q[394] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[393] <= 1'b0;
    end else if(N4798) begin
      tags_q[393] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[392] <= 1'b0;
    end else if(N4798) begin
      tags_q[392] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[391] <= 1'b0;
    end else if(N4798) begin
      tags_q[391] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[390] <= 1'b0;
    end else if(N4798) begin
      tags_q[390] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[389] <= 1'b0;
    end else if(N4798) begin
      tags_q[389] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[388] <= 1'b0;
    end else if(N4798) begin
      tags_q[388] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[387] <= 1'b0;
    end else if(N4798) begin
      tags_q[387] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[386] <= 1'b0;
    end else if(N4798) begin
      tags_q[386] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[385] <= 1'b0;
    end else if(N4798) begin
      tags_q[385] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[384] <= 1'b0;
    end else if(N4798) begin
      tags_q[384] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[383] <= 1'b0;
    end else if(N4798) begin
      tags_q[383] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[382] <= 1'b0;
    end else if(N4798) begin
      tags_q[382] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[381] <= 1'b0;
    end else if(N4798) begin
      tags_q[381] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[380] <= 1'b0;
    end else if(N4798) begin
      tags_q[380] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[379] <= 1'b0;
    end else if(N4798) begin
      tags_q[379] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[378] <= 1'b0;
    end else if(N4798) begin
      tags_q[378] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[377] <= 1'b0;
    end else if(N4798) begin
      tags_q[377] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[376] <= 1'b0;
    end else if(N4798) begin
      tags_q[376] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[375] <= 1'b0;
    end else if(N4798) begin
      tags_q[375] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[374] <= 1'b0;
    end else if(N4798) begin
      tags_q[374] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[373] <= 1'b0;
    end else if(N4798) begin
      tags_q[373] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[372] <= 1'b0;
    end else if(N4801) begin
      tags_q[372] <= tags_n_12__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[371] <= 1'b0;
    end else if(N4803) begin
      tags_q[371] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[370] <= 1'b0;
    end else if(N4803) begin
      tags_q[370] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[369] <= 1'b0;
    end else if(N4803) begin
      tags_q[369] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[368] <= 1'b0;
    end else if(N4803) begin
      tags_q[368] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[367] <= 1'b0;
    end else if(N4803) begin
      tags_q[367] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[366] <= 1'b0;
    end else if(N4803) begin
      tags_q[366] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[365] <= 1'b0;
    end else if(N4803) begin
      tags_q[365] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[364] <= 1'b0;
    end else if(N4803) begin
      tags_q[364] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[363] <= 1'b0;
    end else if(N4803) begin
      tags_q[363] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[362] <= 1'b0;
    end else if(N4803) begin
      tags_q[362] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[361] <= 1'b0;
    end else if(N4803) begin
      tags_q[361] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[360] <= 1'b0;
    end else if(N4803) begin
      tags_q[360] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[359] <= 1'b0;
    end else if(N4803) begin
      tags_q[359] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[358] <= 1'b0;
    end else if(N4803) begin
      tags_q[358] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[357] <= 1'b0;
    end else if(N4803) begin
      tags_q[357] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[356] <= 1'b0;
    end else if(N4803) begin
      tags_q[356] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[355] <= 1'b0;
    end else if(N4803) begin
      tags_q[355] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[354] <= 1'b0;
    end else if(N4803) begin
      tags_q[354] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[353] <= 1'b0;
    end else if(N4803) begin
      tags_q[353] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[352] <= 1'b0;
    end else if(N4803) begin
      tags_q[352] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[351] <= 1'b0;
    end else if(N4803) begin
      tags_q[351] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[350] <= 1'b0;
    end else if(N4803) begin
      tags_q[350] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[349] <= 1'b0;
    end else if(N4803) begin
      tags_q[349] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[348] <= 1'b0;
    end else if(N4803) begin
      tags_q[348] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[347] <= 1'b0;
    end else if(N4803) begin
      tags_q[347] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[346] <= 1'b0;
    end else if(N4803) begin
      tags_q[346] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[345] <= 1'b0;
    end else if(N4803) begin
      tags_q[345] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[344] <= 1'b0;
    end else if(N4803) begin
      tags_q[344] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[343] <= 1'b0;
    end else if(N4803) begin
      tags_q[343] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[342] <= 1'b0;
    end else if(N4803) begin
      tags_q[342] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[341] <= 1'b0;
    end else if(N4806) begin
      tags_q[341] <= tags_n_11__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[340] <= 1'b0;
    end else if(N4808) begin
      tags_q[340] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[339] <= 1'b0;
    end else if(N4808) begin
      tags_q[339] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[338] <= 1'b0;
    end else if(N4808) begin
      tags_q[338] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[337] <= 1'b0;
    end else if(N4808) begin
      tags_q[337] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[336] <= 1'b0;
    end else if(N4808) begin
      tags_q[336] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[335] <= 1'b0;
    end else if(N4808) begin
      tags_q[335] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[334] <= 1'b0;
    end else if(N4808) begin
      tags_q[334] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[333] <= 1'b0;
    end else if(N4808) begin
      tags_q[333] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[332] <= 1'b0;
    end else if(N4808) begin
      tags_q[332] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[331] <= 1'b0;
    end else if(N4808) begin
      tags_q[331] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[330] <= 1'b0;
    end else if(N4808) begin
      tags_q[330] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[329] <= 1'b0;
    end else if(N4808) begin
      tags_q[329] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[328] <= 1'b0;
    end else if(N4808) begin
      tags_q[328] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[327] <= 1'b0;
    end else if(N4808) begin
      tags_q[327] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[326] <= 1'b0;
    end else if(N4808) begin
      tags_q[326] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[325] <= 1'b0;
    end else if(N4808) begin
      tags_q[325] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[324] <= 1'b0;
    end else if(N4808) begin
      tags_q[324] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[323] <= 1'b0;
    end else if(N4808) begin
      tags_q[323] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[322] <= 1'b0;
    end else if(N4808) begin
      tags_q[322] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[321] <= 1'b0;
    end else if(N4808) begin
      tags_q[321] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[320] <= 1'b0;
    end else if(N4808) begin
      tags_q[320] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[319] <= 1'b0;
    end else if(N4808) begin
      tags_q[319] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[318] <= 1'b0;
    end else if(N4808) begin
      tags_q[318] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[317] <= 1'b0;
    end else if(N4808) begin
      tags_q[317] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[316] <= 1'b0;
    end else if(N4808) begin
      tags_q[316] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[315] <= 1'b0;
    end else if(N4808) begin
      tags_q[315] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[314] <= 1'b0;
    end else if(N4808) begin
      tags_q[314] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[313] <= 1'b0;
    end else if(N4808) begin
      tags_q[313] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[312] <= 1'b0;
    end else if(N4808) begin
      tags_q[312] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[311] <= 1'b0;
    end else if(N4808) begin
      tags_q[311] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[310] <= 1'b0;
    end else if(N4811) begin
      tags_q[310] <= tags_n_10__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[309] <= 1'b0;
    end else if(N4813) begin
      tags_q[309] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[308] <= 1'b0;
    end else if(N4813) begin
      tags_q[308] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[307] <= 1'b0;
    end else if(N4813) begin
      tags_q[307] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[306] <= 1'b0;
    end else if(N4813) begin
      tags_q[306] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[305] <= 1'b0;
    end else if(N4813) begin
      tags_q[305] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[304] <= 1'b0;
    end else if(N4813) begin
      tags_q[304] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[303] <= 1'b0;
    end else if(N4813) begin
      tags_q[303] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[302] <= 1'b0;
    end else if(N4813) begin
      tags_q[302] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[301] <= 1'b0;
    end else if(N4813) begin
      tags_q[301] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[300] <= 1'b0;
    end else if(N4813) begin
      tags_q[300] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[299] <= 1'b0;
    end else if(N4813) begin
      tags_q[299] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[298] <= 1'b0;
    end else if(N4813) begin
      tags_q[298] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[297] <= 1'b0;
    end else if(N4813) begin
      tags_q[297] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[296] <= 1'b0;
    end else if(N4813) begin
      tags_q[296] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[295] <= 1'b0;
    end else if(N4813) begin
      tags_q[295] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[294] <= 1'b0;
    end else if(N4813) begin
      tags_q[294] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[293] <= 1'b0;
    end else if(N4813) begin
      tags_q[293] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[292] <= 1'b0;
    end else if(N4813) begin
      tags_q[292] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[291] <= 1'b0;
    end else if(N4813) begin
      tags_q[291] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[290] <= 1'b0;
    end else if(N4813) begin
      tags_q[290] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[289] <= 1'b0;
    end else if(N4813) begin
      tags_q[289] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[288] <= 1'b0;
    end else if(N4813) begin
      tags_q[288] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[287] <= 1'b0;
    end else if(N4813) begin
      tags_q[287] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[286] <= 1'b0;
    end else if(N4813) begin
      tags_q[286] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[285] <= 1'b0;
    end else if(N4813) begin
      tags_q[285] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[284] <= 1'b0;
    end else if(N4813) begin
      tags_q[284] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[283] <= 1'b0;
    end else if(N4813) begin
      tags_q[283] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[282] <= 1'b0;
    end else if(N4813) begin
      tags_q[282] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[281] <= 1'b0;
    end else if(N4813) begin
      tags_q[281] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[280] <= 1'b0;
    end else if(N4813) begin
      tags_q[280] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[279] <= 1'b0;
    end else if(N4816) begin
      tags_q[279] <= tags_n_9__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[278] <= 1'b0;
    end else if(N4818) begin
      tags_q[278] <= update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[277] <= 1'b0;
    end else if(N4818) begin
      tags_q[277] <= update_i[91];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[276] <= 1'b0;
    end else if(N4818) begin
      tags_q[276] <= update_i[90];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[275] <= 1'b0;
    end else if(N4818) begin
      tags_q[275] <= update_i[89];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[274] <= 1'b0;
    end else if(N4818) begin
      tags_q[274] <= update_i[88];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[273] <= 1'b0;
    end else if(N4818) begin
      tags_q[273] <= update_i[87];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[272] <= 1'b0;
    end else if(N4818) begin
      tags_q[272] <= update_i[86];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[271] <= 1'b0;
    end else if(N4818) begin
      tags_q[271] <= update_i[85];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[270] <= 1'b0;
    end else if(N4818) begin
      tags_q[270] <= update_i[84];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[269] <= 1'b0;
    end else if(N4818) begin
      tags_q[269] <= update_i[83];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[268] <= 1'b0;
    end else if(N4818) begin
      tags_q[268] <= update_i[82];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[267] <= 1'b0;
    end else if(N4818) begin
      tags_q[267] <= update_i[81];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[266] <= 1'b0;
    end else if(N4818) begin
      tags_q[266] <= update_i[80];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[265] <= 1'b0;
    end else if(N4818) begin
      tags_q[265] <= update_i[79];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[264] <= 1'b0;
    end else if(N4818) begin
      tags_q[264] <= update_i[78];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[263] <= 1'b0;
    end else if(N4818) begin
      tags_q[263] <= update_i[77];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[262] <= 1'b0;
    end else if(N4818) begin
      tags_q[262] <= update_i[76];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[261] <= 1'b0;
    end else if(N4818) begin
      tags_q[261] <= update_i[75];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[260] <= 1'b0;
    end else if(N4818) begin
      tags_q[260] <= update_i[74];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[259] <= 1'b0;
    end else if(N4818) begin
      tags_q[259] <= update_i[73];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[258] <= 1'b0;
    end else if(N4818) begin
      tags_q[258] <= update_i[72];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[257] <= 1'b0;
    end else if(N4818) begin
      tags_q[257] <= update_i[71];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[256] <= 1'b0;
    end else if(N4818) begin
      tags_q[256] <= update_i[70];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[255] <= 1'b0;
    end else if(N4818) begin
      tags_q[255] <= update_i[69];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[254] <= 1'b0;
    end else if(N4818) begin
      tags_q[254] <= update_i[68];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[253] <= 1'b0;
    end else if(N4818) begin
      tags_q[253] <= update_i[67];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[252] <= 1'b0;
    end else if(N4818) begin
      tags_q[252] <= update_i[66];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[251] <= 1'b0;
    end else if(N4818) begin
      tags_q[251] <= update_i[65];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[250] <= 1'b0;
    end else if(N4818) begin
      tags_q[250] <= update_i[93];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[249] <= 1'b0;
    end else if(N4818) begin
      tags_q[249] <= update_i[92];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[248] <= 1'b0;
    end else if(N4821) begin
      tags_q[248] <= tags_n_8__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[247] <= 1'b0;
    end else if(N4650) begin
      tags_q[247] <= tags_n_7__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[246] <= 1'b0;
    end else if(N4650) begin
      tags_q[246] <= tags_n_7__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[245] <= 1'b0;
    end else if(N4650) begin
      tags_q[245] <= tags_n_7__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[244] <= 1'b0;
    end else if(N4650) begin
      tags_q[244] <= tags_n_7__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[243] <= 1'b0;
    end else if(N4650) begin
      tags_q[243] <= tags_n_7__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[242] <= 1'b0;
    end else if(N4650) begin
      tags_q[242] <= tags_n_7__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[241] <= 1'b0;
    end else if(N4650) begin
      tags_q[241] <= tags_n_7__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[240] <= 1'b0;
    end else if(N4650) begin
      tags_q[240] <= tags_n_7__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[239] <= 1'b0;
    end else if(N4650) begin
      tags_q[239] <= tags_n_7__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[238] <= 1'b0;
    end else if(N4650) begin
      tags_q[238] <= tags_n_7__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[237] <= 1'b0;
    end else if(N4650) begin
      tags_q[237] <= tags_n_7__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[236] <= 1'b0;
    end else if(N4650) begin
      tags_q[236] <= tags_n_7__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[235] <= 1'b0;
    end else if(N4650) begin
      tags_q[235] <= tags_n_7__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[234] <= 1'b0;
    end else if(N4650) begin
      tags_q[234] <= tags_n_7__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[233] <= 1'b0;
    end else if(N4650) begin
      tags_q[233] <= tags_n_7__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[232] <= 1'b0;
    end else if(N4650) begin
      tags_q[232] <= tags_n_7__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[231] <= 1'b0;
    end else if(N4650) begin
      tags_q[231] <= tags_n_7__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[230] <= 1'b0;
    end else if(N4650) begin
      tags_q[230] <= tags_n_7__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[229] <= 1'b0;
    end else if(N4650) begin
      tags_q[229] <= tags_n_7__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[228] <= 1'b0;
    end else if(N4650) begin
      tags_q[228] <= tags_n_7__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[227] <= 1'b0;
    end else if(N4650) begin
      tags_q[227] <= tags_n_7__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[226] <= 1'b0;
    end else if(N4650) begin
      tags_q[226] <= tags_n_7__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[225] <= 1'b0;
    end else if(N4650) begin
      tags_q[225] <= tags_n_7__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[224] <= 1'b0;
    end else if(N4650) begin
      tags_q[224] <= tags_n_7__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[223] <= 1'b0;
    end else if(N4650) begin
      tags_q[223] <= tags_n_7__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[222] <= 1'b0;
    end else if(N4650) begin
      tags_q[222] <= tags_n_7__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[221] <= 1'b0;
    end else if(N4650) begin
      tags_q[221] <= tags_n_7__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[220] <= 1'b0;
    end else if(N4650) begin
      tags_q[220] <= tags_n_7__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[219] <= 1'b0;
    end else if(N4650) begin
      tags_q[219] <= tags_n_7__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[218] <= 1'b0;
    end else if(N4650) begin
      tags_q[218] <= tags_n_7__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[217] <= 1'b0;
    end else if(N4823) begin
      tags_q[217] <= tags_n_7__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[216] <= 1'b0;
    end else if(N4650) begin
      tags_q[216] <= tags_n_6__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[215] <= 1'b0;
    end else if(N4650) begin
      tags_q[215] <= tags_n_6__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[214] <= 1'b0;
    end else if(N4650) begin
      tags_q[214] <= tags_n_6__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[213] <= 1'b0;
    end else if(N4650) begin
      tags_q[213] <= tags_n_6__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[212] <= 1'b0;
    end else if(N4650) begin
      tags_q[212] <= tags_n_6__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[211] <= 1'b0;
    end else if(N4650) begin
      tags_q[211] <= tags_n_6__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[210] <= 1'b0;
    end else if(N4650) begin
      tags_q[210] <= tags_n_6__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[209] <= 1'b0;
    end else if(N4650) begin
      tags_q[209] <= tags_n_6__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[208] <= 1'b0;
    end else if(N4650) begin
      tags_q[208] <= tags_n_6__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[207] <= 1'b0;
    end else if(N4650) begin
      tags_q[207] <= tags_n_6__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[206] <= 1'b0;
    end else if(N4650) begin
      tags_q[206] <= tags_n_6__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[205] <= 1'b0;
    end else if(N4650) begin
      tags_q[205] <= tags_n_6__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[204] <= 1'b0;
    end else if(N4650) begin
      tags_q[204] <= tags_n_6__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[203] <= 1'b0;
    end else if(N4650) begin
      tags_q[203] <= tags_n_6__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[202] <= 1'b0;
    end else if(N4650) begin
      tags_q[202] <= tags_n_6__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[201] <= 1'b0;
    end else if(N4650) begin
      tags_q[201] <= tags_n_6__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[200] <= 1'b0;
    end else if(N4650) begin
      tags_q[200] <= tags_n_6__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[199] <= 1'b0;
    end else if(N4650) begin
      tags_q[199] <= tags_n_6__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[198] <= 1'b0;
    end else if(N4650) begin
      tags_q[198] <= tags_n_6__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[197] <= 1'b0;
    end else if(N4650) begin
      tags_q[197] <= tags_n_6__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[196] <= 1'b0;
    end else if(N4650) begin
      tags_q[196] <= tags_n_6__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[195] <= 1'b0;
    end else if(N4650) begin
      tags_q[195] <= tags_n_6__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[194] <= 1'b0;
    end else if(N4650) begin
      tags_q[194] <= tags_n_6__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[193] <= 1'b0;
    end else if(N4650) begin
      tags_q[193] <= tags_n_6__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[192] <= 1'b0;
    end else if(N4650) begin
      tags_q[192] <= tags_n_6__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[191] <= 1'b0;
    end else if(N4650) begin
      tags_q[191] <= tags_n_6__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[190] <= 1'b0;
    end else if(N4650) begin
      tags_q[190] <= tags_n_6__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[189] <= 1'b0;
    end else if(N4650) begin
      tags_q[189] <= tags_n_6__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[188] <= 1'b0;
    end else if(N4650) begin
      tags_q[188] <= tags_n_6__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[187] <= 1'b0;
    end else if(N4650) begin
      tags_q[187] <= tags_n_6__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[186] <= 1'b0;
    end else if(N4825) begin
      tags_q[186] <= tags_n_6__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[185] <= 1'b0;
    end else if(N4650) begin
      tags_q[185] <= tags_n_5__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[184] <= 1'b0;
    end else if(N4650) begin
      tags_q[184] <= tags_n_5__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[183] <= 1'b0;
    end else if(N4650) begin
      tags_q[183] <= tags_n_5__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[182] <= 1'b0;
    end else if(N4650) begin
      tags_q[182] <= tags_n_5__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[181] <= 1'b0;
    end else if(N4650) begin
      tags_q[181] <= tags_n_5__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[180] <= 1'b0;
    end else if(N4650) begin
      tags_q[180] <= tags_n_5__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[179] <= 1'b0;
    end else if(N4650) begin
      tags_q[179] <= tags_n_5__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[178] <= 1'b0;
    end else if(N4650) begin
      tags_q[178] <= tags_n_5__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[177] <= 1'b0;
    end else if(N4650) begin
      tags_q[177] <= tags_n_5__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[176] <= 1'b0;
    end else if(N4650) begin
      tags_q[176] <= tags_n_5__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[175] <= 1'b0;
    end else if(N4650) begin
      tags_q[175] <= tags_n_5__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[174] <= 1'b0;
    end else if(N4650) begin
      tags_q[174] <= tags_n_5__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[173] <= 1'b0;
    end else if(N4650) begin
      tags_q[173] <= tags_n_5__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[172] <= 1'b0;
    end else if(N4650) begin
      tags_q[172] <= tags_n_5__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[171] <= 1'b0;
    end else if(N4650) begin
      tags_q[171] <= tags_n_5__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[170] <= 1'b0;
    end else if(N4650) begin
      tags_q[170] <= tags_n_5__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[169] <= 1'b0;
    end else if(N4650) begin
      tags_q[169] <= tags_n_5__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[168] <= 1'b0;
    end else if(N4650) begin
      tags_q[168] <= tags_n_5__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[167] <= 1'b0;
    end else if(N4650) begin
      tags_q[167] <= tags_n_5__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[166] <= 1'b0;
    end else if(N4650) begin
      tags_q[166] <= tags_n_5__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[165] <= 1'b0;
    end else if(N4650) begin
      tags_q[165] <= tags_n_5__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[164] <= 1'b0;
    end else if(N4650) begin
      tags_q[164] <= tags_n_5__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[163] <= 1'b0;
    end else if(N4650) begin
      tags_q[163] <= tags_n_5__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[162] <= 1'b0;
    end else if(N4650) begin
      tags_q[162] <= tags_n_5__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[161] <= 1'b0;
    end else if(N4650) begin
      tags_q[161] <= tags_n_5__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[160] <= 1'b0;
    end else if(N4650) begin
      tags_q[160] <= tags_n_5__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[159] <= 1'b0;
    end else if(N4650) begin
      tags_q[159] <= tags_n_5__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[158] <= 1'b0;
    end else if(N4650) begin
      tags_q[158] <= tags_n_5__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[157] <= 1'b0;
    end else if(N4650) begin
      tags_q[157] <= tags_n_5__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[156] <= 1'b0;
    end else if(N4650) begin
      tags_q[156] <= tags_n_5__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[155] <= 1'b0;
    end else if(N4827) begin
      tags_q[155] <= tags_n_5__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[154] <= 1'b0;
    end else if(N4650) begin
      tags_q[154] <= tags_n_4__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[153] <= 1'b0;
    end else if(N4650) begin
      tags_q[153] <= tags_n_4__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[152] <= 1'b0;
    end else if(N4650) begin
      tags_q[152] <= tags_n_4__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[151] <= 1'b0;
    end else if(N4650) begin
      tags_q[151] <= tags_n_4__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[150] <= 1'b0;
    end else if(N4650) begin
      tags_q[150] <= tags_n_4__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[149] <= 1'b0;
    end else if(N4650) begin
      tags_q[149] <= tags_n_4__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[148] <= 1'b0;
    end else if(N4650) begin
      tags_q[148] <= tags_n_4__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[147] <= 1'b0;
    end else if(N4650) begin
      tags_q[147] <= tags_n_4__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[146] <= 1'b0;
    end else if(N4650) begin
      tags_q[146] <= tags_n_4__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[145] <= 1'b0;
    end else if(N4650) begin
      tags_q[145] <= tags_n_4__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[144] <= 1'b0;
    end else if(N4650) begin
      tags_q[144] <= tags_n_4__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[143] <= 1'b0;
    end else if(N4650) begin
      tags_q[143] <= tags_n_4__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[142] <= 1'b0;
    end else if(N4650) begin
      tags_q[142] <= tags_n_4__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[141] <= 1'b0;
    end else if(N4650) begin
      tags_q[141] <= tags_n_4__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[140] <= 1'b0;
    end else if(N4650) begin
      tags_q[140] <= tags_n_4__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[139] <= 1'b0;
    end else if(N4650) begin
      tags_q[139] <= tags_n_4__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[138] <= 1'b0;
    end else if(N4650) begin
      tags_q[138] <= tags_n_4__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[137] <= 1'b0;
    end else if(N4650) begin
      tags_q[137] <= tags_n_4__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[136] <= 1'b0;
    end else if(N4650) begin
      tags_q[136] <= tags_n_4__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[135] <= 1'b0;
    end else if(N4650) begin
      tags_q[135] <= tags_n_4__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[134] <= 1'b0;
    end else if(N4650) begin
      tags_q[134] <= tags_n_4__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[133] <= 1'b0;
    end else if(N4650) begin
      tags_q[133] <= tags_n_4__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[132] <= 1'b0;
    end else if(N4650) begin
      tags_q[132] <= tags_n_4__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[131] <= 1'b0;
    end else if(N4650) begin
      tags_q[131] <= tags_n_4__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[130] <= 1'b0;
    end else if(N4650) begin
      tags_q[130] <= tags_n_4__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[129] <= 1'b0;
    end else if(N4650) begin
      tags_q[129] <= tags_n_4__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[128] <= 1'b0;
    end else if(N4650) begin
      tags_q[128] <= tags_n_4__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[127] <= 1'b0;
    end else if(N4650) begin
      tags_q[127] <= tags_n_4__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[126] <= 1'b0;
    end else if(N4650) begin
      tags_q[126] <= tags_n_4__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[125] <= 1'b0;
    end else if(N4650) begin
      tags_q[125] <= tags_n_4__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[124] <= 1'b0;
    end else if(N4829) begin
      tags_q[124] <= tags_n_4__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[123] <= 1'b0;
    end else if(N4650) begin
      tags_q[123] <= tags_n_3__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[122] <= 1'b0;
    end else if(N4650) begin
      tags_q[122] <= tags_n_3__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[121] <= 1'b0;
    end else if(N4650) begin
      tags_q[121] <= tags_n_3__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[120] <= 1'b0;
    end else if(N4650) begin
      tags_q[120] <= tags_n_3__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[119] <= 1'b0;
    end else if(N4650) begin
      tags_q[119] <= tags_n_3__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[118] <= 1'b0;
    end else if(N4650) begin
      tags_q[118] <= tags_n_3__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[117] <= 1'b0;
    end else if(N4650) begin
      tags_q[117] <= tags_n_3__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[116] <= 1'b0;
    end else if(N4650) begin
      tags_q[116] <= tags_n_3__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[115] <= 1'b0;
    end else if(N4650) begin
      tags_q[115] <= tags_n_3__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[114] <= 1'b0;
    end else if(N4650) begin
      tags_q[114] <= tags_n_3__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[113] <= 1'b0;
    end else if(N4650) begin
      tags_q[113] <= tags_n_3__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[112] <= 1'b0;
    end else if(N4650) begin
      tags_q[112] <= tags_n_3__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[111] <= 1'b0;
    end else if(N4650) begin
      tags_q[111] <= tags_n_3__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[110] <= 1'b0;
    end else if(N4650) begin
      tags_q[110] <= tags_n_3__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[109] <= 1'b0;
    end else if(N4650) begin
      tags_q[109] <= tags_n_3__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[108] <= 1'b0;
    end else if(N4650) begin
      tags_q[108] <= tags_n_3__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[107] <= 1'b0;
    end else if(N4650) begin
      tags_q[107] <= tags_n_3__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[106] <= 1'b0;
    end else if(N4650) begin
      tags_q[106] <= tags_n_3__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[105] <= 1'b0;
    end else if(N4650) begin
      tags_q[105] <= tags_n_3__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[104] <= 1'b0;
    end else if(N4650) begin
      tags_q[104] <= tags_n_3__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[103] <= 1'b0;
    end else if(N4650) begin
      tags_q[103] <= tags_n_3__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[102] <= 1'b0;
    end else if(N4650) begin
      tags_q[102] <= tags_n_3__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[101] <= 1'b0;
    end else if(N4650) begin
      tags_q[101] <= tags_n_3__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[100] <= 1'b0;
    end else if(N4650) begin
      tags_q[100] <= tags_n_3__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[99] <= 1'b0;
    end else if(N4650) begin
      tags_q[99] <= tags_n_3__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[98] <= 1'b0;
    end else if(N4650) begin
      tags_q[98] <= tags_n_3__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[97] <= 1'b0;
    end else if(N4650) begin
      tags_q[97] <= tags_n_3__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[96] <= 1'b0;
    end else if(N4650) begin
      tags_q[96] <= tags_n_3__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[95] <= 1'b0;
    end else if(N4650) begin
      tags_q[95] <= tags_n_3__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[94] <= 1'b0;
    end else if(N4650) begin
      tags_q[94] <= tags_n_3__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[93] <= 1'b0;
    end else if(N4831) begin
      tags_q[93] <= tags_n_3__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[92] <= 1'b0;
    end else if(N4650) begin
      tags_q[92] <= tags_n_2__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[91] <= 1'b0;
    end else if(N4650) begin
      tags_q[91] <= tags_n_2__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[90] <= 1'b0;
    end else if(N4650) begin
      tags_q[90] <= tags_n_2__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[89] <= 1'b0;
    end else if(N4650) begin
      tags_q[89] <= tags_n_2__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[88] <= 1'b0;
    end else if(N4650) begin
      tags_q[88] <= tags_n_2__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[87] <= 1'b0;
    end else if(N4650) begin
      tags_q[87] <= tags_n_2__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[86] <= 1'b0;
    end else if(N4650) begin
      tags_q[86] <= tags_n_2__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[85] <= 1'b0;
    end else if(N4650) begin
      tags_q[85] <= tags_n_2__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[84] <= 1'b0;
    end else if(N4650) begin
      tags_q[84] <= tags_n_2__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[83] <= 1'b0;
    end else if(N4650) begin
      tags_q[83] <= tags_n_2__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[82] <= 1'b0;
    end else if(N4650) begin
      tags_q[82] <= tags_n_2__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[81] <= 1'b0;
    end else if(N4650) begin
      tags_q[81] <= tags_n_2__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[80] <= 1'b0;
    end else if(N4650) begin
      tags_q[80] <= tags_n_2__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[79] <= 1'b0;
    end else if(N4650) begin
      tags_q[79] <= tags_n_2__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[78] <= 1'b0;
    end else if(N4650) begin
      tags_q[78] <= tags_n_2__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[77] <= 1'b0;
    end else if(N4650) begin
      tags_q[77] <= tags_n_2__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[76] <= 1'b0;
    end else if(N4650) begin
      tags_q[76] <= tags_n_2__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[75] <= 1'b0;
    end else if(N4650) begin
      tags_q[75] <= tags_n_2__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[74] <= 1'b0;
    end else if(N4650) begin
      tags_q[74] <= tags_n_2__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[73] <= 1'b0;
    end else if(N4650) begin
      tags_q[73] <= tags_n_2__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[72] <= 1'b0;
    end else if(N4650) begin
      tags_q[72] <= tags_n_2__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[71] <= 1'b0;
    end else if(N4650) begin
      tags_q[71] <= tags_n_2__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[70] <= 1'b0;
    end else if(N4650) begin
      tags_q[70] <= tags_n_2__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[69] <= 1'b0;
    end else if(N4650) begin
      tags_q[69] <= tags_n_2__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[68] <= 1'b0;
    end else if(N4650) begin
      tags_q[68] <= tags_n_2__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[67] <= 1'b0;
    end else if(N4650) begin
      tags_q[67] <= tags_n_2__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[66] <= 1'b0;
    end else if(N4650) begin
      tags_q[66] <= tags_n_2__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[65] <= 1'b0;
    end else if(N4650) begin
      tags_q[65] <= tags_n_2__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[64] <= 1'b0;
    end else if(N4650) begin
      tags_q[64] <= tags_n_2__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[63] <= 1'b0;
    end else if(N4650) begin
      tags_q[63] <= tags_n_2__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[62] <= 1'b0;
    end else if(N4833) begin
      tags_q[62] <= tags_n_2__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[61] <= 1'b0;
    end else if(N4650) begin
      tags_q[61] <= tags_n_1__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[60] <= 1'b0;
    end else if(N4650) begin
      tags_q[60] <= tags_n_1__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[59] <= 1'b0;
    end else if(N4650) begin
      tags_q[59] <= tags_n_1__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[58] <= 1'b0;
    end else if(N4650) begin
      tags_q[58] <= tags_n_1__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[57] <= 1'b0;
    end else if(N4650) begin
      tags_q[57] <= tags_n_1__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[56] <= 1'b0;
    end else if(N4650) begin
      tags_q[56] <= tags_n_1__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[55] <= 1'b0;
    end else if(N4650) begin
      tags_q[55] <= tags_n_1__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[54] <= 1'b0;
    end else if(N4650) begin
      tags_q[54] <= tags_n_1__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[53] <= 1'b0;
    end else if(N4650) begin
      tags_q[53] <= tags_n_1__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[52] <= 1'b0;
    end else if(N4650) begin
      tags_q[52] <= tags_n_1__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[51] <= 1'b0;
    end else if(N4650) begin
      tags_q[51] <= tags_n_1__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[50] <= 1'b0;
    end else if(N4650) begin
      tags_q[50] <= tags_n_1__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[49] <= 1'b0;
    end else if(N4650) begin
      tags_q[49] <= tags_n_1__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[48] <= 1'b0;
    end else if(N4650) begin
      tags_q[48] <= tags_n_1__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[47] <= 1'b0;
    end else if(N4650) begin
      tags_q[47] <= tags_n_1__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[46] <= 1'b0;
    end else if(N4650) begin
      tags_q[46] <= tags_n_1__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[45] <= 1'b0;
    end else if(N4650) begin
      tags_q[45] <= tags_n_1__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[44] <= 1'b0;
    end else if(N4650) begin
      tags_q[44] <= tags_n_1__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[43] <= 1'b0;
    end else if(N4650) begin
      tags_q[43] <= tags_n_1__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[42] <= 1'b0;
    end else if(N4650) begin
      tags_q[42] <= tags_n_1__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[41] <= 1'b0;
    end else if(N4650) begin
      tags_q[41] <= tags_n_1__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[40] <= 1'b0;
    end else if(N4650) begin
      tags_q[40] <= tags_n_1__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[39] <= 1'b0;
    end else if(N4650) begin
      tags_q[39] <= tags_n_1__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[38] <= 1'b0;
    end else if(N4650) begin
      tags_q[38] <= tags_n_1__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[37] <= 1'b0;
    end else if(N4650) begin
      tags_q[37] <= tags_n_1__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[36] <= 1'b0;
    end else if(N4650) begin
      tags_q[36] <= tags_n_1__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[35] <= 1'b0;
    end else if(N4650) begin
      tags_q[35] <= tags_n_1__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[34] <= 1'b0;
    end else if(N4650) begin
      tags_q[34] <= tags_n_1__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[33] <= 1'b0;
    end else if(N4650) begin
      tags_q[33] <= tags_n_1__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[32] <= 1'b0;
    end else if(N4650) begin
      tags_q[32] <= tags_n_1__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[31] <= 1'b0;
    end else if(N4835) begin
      tags_q[31] <= tags_n_1__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[30] <= 1'b0;
    end else if(N4650) begin
      tags_q[30] <= tags_n_0__asid__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[29] <= 1'b0;
    end else if(N4650) begin
      tags_q[29] <= tags_n_0__vpn2__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[28] <= 1'b0;
    end else if(N4650) begin
      tags_q[28] <= tags_n_0__vpn2__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[27] <= 1'b0;
    end else if(N4650) begin
      tags_q[27] <= tags_n_0__vpn2__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[26] <= 1'b0;
    end else if(N4650) begin
      tags_q[26] <= tags_n_0__vpn2__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[25] <= 1'b0;
    end else if(N4650) begin
      tags_q[25] <= tags_n_0__vpn2__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[24] <= 1'b0;
    end else if(N4650) begin
      tags_q[24] <= tags_n_0__vpn2__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[23] <= 1'b0;
    end else if(N4650) begin
      tags_q[23] <= tags_n_0__vpn2__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[22] <= 1'b0;
    end else if(N4650) begin
      tags_q[22] <= tags_n_0__vpn2__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[21] <= 1'b0;
    end else if(N4650) begin
      tags_q[21] <= tags_n_0__vpn2__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[20] <= 1'b0;
    end else if(N4650) begin
      tags_q[20] <= tags_n_0__vpn1__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[19] <= 1'b0;
    end else if(N4650) begin
      tags_q[19] <= tags_n_0__vpn1__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[18] <= 1'b0;
    end else if(N4650) begin
      tags_q[18] <= tags_n_0__vpn1__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[17] <= 1'b0;
    end else if(N4650) begin
      tags_q[17] <= tags_n_0__vpn1__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[16] <= 1'b0;
    end else if(N4650) begin
      tags_q[16] <= tags_n_0__vpn1__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[15] <= 1'b0;
    end else if(N4650) begin
      tags_q[15] <= tags_n_0__vpn1__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[14] <= 1'b0;
    end else if(N4650) begin
      tags_q[14] <= tags_n_0__vpn1__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[13] <= 1'b0;
    end else if(N4650) begin
      tags_q[13] <= tags_n_0__vpn1__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[12] <= 1'b0;
    end else if(N4650) begin
      tags_q[12] <= tags_n_0__vpn1__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[11] <= 1'b0;
    end else if(N4650) begin
      tags_q[11] <= tags_n_0__vpn0__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[10] <= 1'b0;
    end else if(N4650) begin
      tags_q[10] <= tags_n_0__vpn0__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[9] <= 1'b0;
    end else if(N4650) begin
      tags_q[9] <= tags_n_0__vpn0__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[8] <= 1'b0;
    end else if(N4650) begin
      tags_q[8] <= tags_n_0__vpn0__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[7] <= 1'b0;
    end else if(N4650) begin
      tags_q[7] <= tags_n_0__vpn0__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[6] <= 1'b0;
    end else if(N4650) begin
      tags_q[6] <= tags_n_0__vpn0__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[5] <= 1'b0;
    end else if(N4650) begin
      tags_q[5] <= tags_n_0__vpn0__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[4] <= 1'b0;
    end else if(N4650) begin
      tags_q[4] <= tags_n_0__vpn0__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[3] <= 1'b0;
    end else if(N4650) begin
      tags_q[3] <= tags_n_0__vpn0__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[2] <= 1'b0;
    end else if(N4650) begin
      tags_q[2] <= tags_n_0__is_2M_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[1] <= 1'b0;
    end else if(N4650) begin
      tags_q[1] <= tags_n_0__is_1G_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      tags_q[0] <= 1'b0;
    end else if(N4837) begin
      tags_q[0] <= tags_n_0__valid_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1023] <= 1'b0;
    end else if(N4783) begin
      content_q[1023] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1022] <= 1'b0;
    end else if(N4783) begin
      content_q[1022] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1021] <= 1'b0;
    end else if(N4783) begin
      content_q[1021] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1020] <= 1'b0;
    end else if(N4783) begin
      content_q[1020] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1019] <= 1'b0;
    end else if(N4783) begin
      content_q[1019] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1018] <= 1'b0;
    end else if(N4783) begin
      content_q[1018] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1017] <= 1'b0;
    end else if(N4783) begin
      content_q[1017] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1016] <= 1'b0;
    end else if(N4783) begin
      content_q[1016] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1015] <= 1'b0;
    end else if(N4783) begin
      content_q[1015] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1014] <= 1'b0;
    end else if(N4783) begin
      content_q[1014] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1013] <= 1'b0;
    end else if(N4783) begin
      content_q[1013] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1012] <= 1'b0;
    end else if(N4783) begin
      content_q[1012] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1011] <= 1'b0;
    end else if(N4783) begin
      content_q[1011] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1010] <= 1'b0;
    end else if(N4783) begin
      content_q[1010] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1009] <= 1'b0;
    end else if(N4783) begin
      content_q[1009] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1008] <= 1'b0;
    end else if(N4783) begin
      content_q[1008] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1007] <= 1'b0;
    end else if(N4783) begin
      content_q[1007] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1006] <= 1'b0;
    end else if(N4783) begin
      content_q[1006] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1005] <= 1'b0;
    end else if(N4783) begin
      content_q[1005] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1004] <= 1'b0;
    end else if(N4783) begin
      content_q[1004] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1003] <= 1'b0;
    end else if(N4783) begin
      content_q[1003] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1002] <= 1'b0;
    end else if(N4783) begin
      content_q[1002] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1001] <= 1'b0;
    end else if(N4783) begin
      content_q[1001] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1000] <= 1'b0;
    end else if(N4783) begin
      content_q[1000] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[999] <= 1'b0;
    end else if(N4783) begin
      content_q[999] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[998] <= 1'b0;
    end else if(N4783) begin
      content_q[998] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[997] <= 1'b0;
    end else if(N4783) begin
      content_q[997] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[996] <= 1'b0;
    end else if(N4783) begin
      content_q[996] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[995] <= 1'b0;
    end else if(N4783) begin
      content_q[995] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[994] <= 1'b0;
    end else if(N4783) begin
      content_q[994] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[993] <= 1'b0;
    end else if(N4783) begin
      content_q[993] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[992] <= 1'b0;
    end else if(N4783) begin
      content_q[992] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[991] <= 1'b0;
    end else if(N4783) begin
      content_q[991] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[990] <= 1'b0;
    end else if(N4783) begin
      content_q[990] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[989] <= 1'b0;
    end else if(N4783) begin
      content_q[989] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[988] <= 1'b0;
    end else if(N4783) begin
      content_q[988] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[987] <= 1'b0;
    end else if(N4783) begin
      content_q[987] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[986] <= 1'b0;
    end else if(N4783) begin
      content_q[986] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[985] <= 1'b0;
    end else if(N4783) begin
      content_q[985] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[984] <= 1'b0;
    end else if(N4783) begin
      content_q[984] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[983] <= 1'b0;
    end else if(N4783) begin
      content_q[983] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[982] <= 1'b0;
    end else if(N4783) begin
      content_q[982] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[981] <= 1'b0;
    end else if(N4783) begin
      content_q[981] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[980] <= 1'b0;
    end else if(N4783) begin
      content_q[980] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[979] <= 1'b0;
    end else if(N4783) begin
      content_q[979] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[978] <= 1'b0;
    end else if(N4783) begin
      content_q[978] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[977] <= 1'b0;
    end else if(N4783) begin
      content_q[977] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[976] <= 1'b0;
    end else if(N4783) begin
      content_q[976] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[975] <= 1'b0;
    end else if(N4783) begin
      content_q[975] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[974] <= 1'b0;
    end else if(N4783) begin
      content_q[974] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[973] <= 1'b0;
    end else if(N4783) begin
      content_q[973] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[972] <= 1'b0;
    end else if(N4783) begin
      content_q[972] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[971] <= 1'b0;
    end else if(N4783) begin
      content_q[971] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[970] <= 1'b0;
    end else if(N4783) begin
      content_q[970] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[969] <= 1'b0;
    end else if(N4783) begin
      content_q[969] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[968] <= 1'b0;
    end else if(N4783) begin
      content_q[968] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[967] <= 1'b0;
    end else if(N4783) begin
      content_q[967] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[966] <= 1'b0;
    end else if(N4783) begin
      content_q[966] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[965] <= 1'b0;
    end else if(N4783) begin
      content_q[965] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[964] <= 1'b0;
    end else if(N4783) begin
      content_q[964] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[963] <= 1'b0;
    end else if(N4783) begin
      content_q[963] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[962] <= 1'b0;
    end else if(N4783) begin
      content_q[962] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[961] <= 1'b0;
    end else if(N4783) begin
      content_q[961] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[960] <= 1'b0;
    end else if(N4783) begin
      content_q[960] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[959] <= 1'b0;
    end else if(N4788) begin
      content_q[959] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[958] <= 1'b0;
    end else if(N4788) begin
      content_q[958] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[957] <= 1'b0;
    end else if(N4788) begin
      content_q[957] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[956] <= 1'b0;
    end else if(N4788) begin
      content_q[956] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[955] <= 1'b0;
    end else if(N4788) begin
      content_q[955] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[954] <= 1'b0;
    end else if(N4788) begin
      content_q[954] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[953] <= 1'b0;
    end else if(N4788) begin
      content_q[953] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[952] <= 1'b0;
    end else if(N4788) begin
      content_q[952] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[951] <= 1'b0;
    end else if(N4788) begin
      content_q[951] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[950] <= 1'b0;
    end else if(N4788) begin
      content_q[950] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[949] <= 1'b0;
    end else if(N4788) begin
      content_q[949] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[948] <= 1'b0;
    end else if(N4788) begin
      content_q[948] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[947] <= 1'b0;
    end else if(N4788) begin
      content_q[947] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[946] <= 1'b0;
    end else if(N4788) begin
      content_q[946] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[945] <= 1'b0;
    end else if(N4788) begin
      content_q[945] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[944] <= 1'b0;
    end else if(N4788) begin
      content_q[944] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[943] <= 1'b0;
    end else if(N4788) begin
      content_q[943] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[942] <= 1'b0;
    end else if(N4788) begin
      content_q[942] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[941] <= 1'b0;
    end else if(N4788) begin
      content_q[941] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[940] <= 1'b0;
    end else if(N4788) begin
      content_q[940] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[939] <= 1'b0;
    end else if(N4788) begin
      content_q[939] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[938] <= 1'b0;
    end else if(N4788) begin
      content_q[938] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[937] <= 1'b0;
    end else if(N4788) begin
      content_q[937] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[936] <= 1'b0;
    end else if(N4788) begin
      content_q[936] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[935] <= 1'b0;
    end else if(N4788) begin
      content_q[935] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[934] <= 1'b0;
    end else if(N4788) begin
      content_q[934] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[933] <= 1'b0;
    end else if(N4788) begin
      content_q[933] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[932] <= 1'b0;
    end else if(N4788) begin
      content_q[932] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[931] <= 1'b0;
    end else if(N4788) begin
      content_q[931] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[930] <= 1'b0;
    end else if(N4788) begin
      content_q[930] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[929] <= 1'b0;
    end else if(N4788) begin
      content_q[929] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[928] <= 1'b0;
    end else if(N4788) begin
      content_q[928] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[927] <= 1'b0;
    end else if(N4788) begin
      content_q[927] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[926] <= 1'b0;
    end else if(N4788) begin
      content_q[926] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[925] <= 1'b0;
    end else if(N4788) begin
      content_q[925] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[924] <= 1'b0;
    end else if(N4788) begin
      content_q[924] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[923] <= 1'b0;
    end else if(N4788) begin
      content_q[923] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[922] <= 1'b0;
    end else if(N4788) begin
      content_q[922] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[921] <= 1'b0;
    end else if(N4788) begin
      content_q[921] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[920] <= 1'b0;
    end else if(N4788) begin
      content_q[920] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[919] <= 1'b0;
    end else if(N4788) begin
      content_q[919] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[918] <= 1'b0;
    end else if(N4788) begin
      content_q[918] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[917] <= 1'b0;
    end else if(N4788) begin
      content_q[917] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[916] <= 1'b0;
    end else if(N4788) begin
      content_q[916] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[915] <= 1'b0;
    end else if(N4788) begin
      content_q[915] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[914] <= 1'b0;
    end else if(N4788) begin
      content_q[914] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[913] <= 1'b0;
    end else if(N4788) begin
      content_q[913] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[912] <= 1'b0;
    end else if(N4788) begin
      content_q[912] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[911] <= 1'b0;
    end else if(N4788) begin
      content_q[911] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[910] <= 1'b0;
    end else if(N4788) begin
      content_q[910] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[909] <= 1'b0;
    end else if(N4788) begin
      content_q[909] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[908] <= 1'b0;
    end else if(N4788) begin
      content_q[908] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[907] <= 1'b0;
    end else if(N4788) begin
      content_q[907] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[906] <= 1'b0;
    end else if(N4788) begin
      content_q[906] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[905] <= 1'b0;
    end else if(N4788) begin
      content_q[905] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[904] <= 1'b0;
    end else if(N4788) begin
      content_q[904] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[903] <= 1'b0;
    end else if(N4788) begin
      content_q[903] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[902] <= 1'b0;
    end else if(N4788) begin
      content_q[902] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[901] <= 1'b0;
    end else if(N4788) begin
      content_q[901] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[900] <= 1'b0;
    end else if(N4788) begin
      content_q[900] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[899] <= 1'b0;
    end else if(N4788) begin
      content_q[899] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[898] <= 1'b0;
    end else if(N4788) begin
      content_q[898] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[897] <= 1'b0;
    end else if(N4788) begin
      content_q[897] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[896] <= 1'b0;
    end else if(N4788) begin
      content_q[896] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[895] <= 1'b0;
    end else if(N4793) begin
      content_q[895] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[894] <= 1'b0;
    end else if(N4793) begin
      content_q[894] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[893] <= 1'b0;
    end else if(N4793) begin
      content_q[893] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[892] <= 1'b0;
    end else if(N4793) begin
      content_q[892] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[891] <= 1'b0;
    end else if(N4793) begin
      content_q[891] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[890] <= 1'b0;
    end else if(N4793) begin
      content_q[890] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[889] <= 1'b0;
    end else if(N4793) begin
      content_q[889] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[888] <= 1'b0;
    end else if(N4793) begin
      content_q[888] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[887] <= 1'b0;
    end else if(N4793) begin
      content_q[887] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[886] <= 1'b0;
    end else if(N4793) begin
      content_q[886] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[885] <= 1'b0;
    end else if(N4793) begin
      content_q[885] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[884] <= 1'b0;
    end else if(N4793) begin
      content_q[884] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[883] <= 1'b0;
    end else if(N4793) begin
      content_q[883] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[882] <= 1'b0;
    end else if(N4793) begin
      content_q[882] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[881] <= 1'b0;
    end else if(N4793) begin
      content_q[881] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[880] <= 1'b0;
    end else if(N4793) begin
      content_q[880] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[879] <= 1'b0;
    end else if(N4793) begin
      content_q[879] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[878] <= 1'b0;
    end else if(N4793) begin
      content_q[878] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[877] <= 1'b0;
    end else if(N4793) begin
      content_q[877] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[876] <= 1'b0;
    end else if(N4793) begin
      content_q[876] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[875] <= 1'b0;
    end else if(N4793) begin
      content_q[875] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[874] <= 1'b0;
    end else if(N4793) begin
      content_q[874] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[873] <= 1'b0;
    end else if(N4793) begin
      content_q[873] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[872] <= 1'b0;
    end else if(N4793) begin
      content_q[872] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[871] <= 1'b0;
    end else if(N4793) begin
      content_q[871] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[870] <= 1'b0;
    end else if(N4793) begin
      content_q[870] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[869] <= 1'b0;
    end else if(N4793) begin
      content_q[869] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[868] <= 1'b0;
    end else if(N4793) begin
      content_q[868] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[867] <= 1'b0;
    end else if(N4793) begin
      content_q[867] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[866] <= 1'b0;
    end else if(N4793) begin
      content_q[866] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[865] <= 1'b0;
    end else if(N4793) begin
      content_q[865] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[864] <= 1'b0;
    end else if(N4793) begin
      content_q[864] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[863] <= 1'b0;
    end else if(N4793) begin
      content_q[863] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[862] <= 1'b0;
    end else if(N4793) begin
      content_q[862] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[861] <= 1'b0;
    end else if(N4793) begin
      content_q[861] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[860] <= 1'b0;
    end else if(N4793) begin
      content_q[860] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[859] <= 1'b0;
    end else if(N4793) begin
      content_q[859] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[858] <= 1'b0;
    end else if(N4793) begin
      content_q[858] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[857] <= 1'b0;
    end else if(N4793) begin
      content_q[857] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[856] <= 1'b0;
    end else if(N4793) begin
      content_q[856] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[855] <= 1'b0;
    end else if(N4793) begin
      content_q[855] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[854] <= 1'b0;
    end else if(N4793) begin
      content_q[854] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[853] <= 1'b0;
    end else if(N4793) begin
      content_q[853] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[852] <= 1'b0;
    end else if(N4793) begin
      content_q[852] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[851] <= 1'b0;
    end else if(N4793) begin
      content_q[851] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[850] <= 1'b0;
    end else if(N4793) begin
      content_q[850] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[849] <= 1'b0;
    end else if(N4793) begin
      content_q[849] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[848] <= 1'b0;
    end else if(N4793) begin
      content_q[848] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[847] <= 1'b0;
    end else if(N4793) begin
      content_q[847] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[846] <= 1'b0;
    end else if(N4793) begin
      content_q[846] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[845] <= 1'b0;
    end else if(N4793) begin
      content_q[845] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[844] <= 1'b0;
    end else if(N4793) begin
      content_q[844] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[843] <= 1'b0;
    end else if(N4793) begin
      content_q[843] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[842] <= 1'b0;
    end else if(N4793) begin
      content_q[842] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[841] <= 1'b0;
    end else if(N4793) begin
      content_q[841] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[840] <= 1'b0;
    end else if(N4793) begin
      content_q[840] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[839] <= 1'b0;
    end else if(N4793) begin
      content_q[839] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[838] <= 1'b0;
    end else if(N4793) begin
      content_q[838] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[837] <= 1'b0;
    end else if(N4793) begin
      content_q[837] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[836] <= 1'b0;
    end else if(N4793) begin
      content_q[836] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[835] <= 1'b0;
    end else if(N4793) begin
      content_q[835] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[834] <= 1'b0;
    end else if(N4793) begin
      content_q[834] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[833] <= 1'b0;
    end else if(N4793) begin
      content_q[833] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[832] <= 1'b0;
    end else if(N4793) begin
      content_q[832] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[831] <= 1'b0;
    end else if(N4798) begin
      content_q[831] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[830] <= 1'b0;
    end else if(N4798) begin
      content_q[830] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[829] <= 1'b0;
    end else if(N4798) begin
      content_q[829] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[828] <= 1'b0;
    end else if(N4798) begin
      content_q[828] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[827] <= 1'b0;
    end else if(N4798) begin
      content_q[827] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[826] <= 1'b0;
    end else if(N4798) begin
      content_q[826] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[825] <= 1'b0;
    end else if(N4798) begin
      content_q[825] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[824] <= 1'b0;
    end else if(N4798) begin
      content_q[824] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[823] <= 1'b0;
    end else if(N4798) begin
      content_q[823] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[822] <= 1'b0;
    end else if(N4798) begin
      content_q[822] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[821] <= 1'b0;
    end else if(N4798) begin
      content_q[821] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[820] <= 1'b0;
    end else if(N4798) begin
      content_q[820] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[819] <= 1'b0;
    end else if(N4798) begin
      content_q[819] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[818] <= 1'b0;
    end else if(N4798) begin
      content_q[818] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[817] <= 1'b0;
    end else if(N4798) begin
      content_q[817] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[816] <= 1'b0;
    end else if(N4798) begin
      content_q[816] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[815] <= 1'b0;
    end else if(N4798) begin
      content_q[815] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[814] <= 1'b0;
    end else if(N4798) begin
      content_q[814] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[813] <= 1'b0;
    end else if(N4798) begin
      content_q[813] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[812] <= 1'b0;
    end else if(N4798) begin
      content_q[812] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[811] <= 1'b0;
    end else if(N4798) begin
      content_q[811] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[810] <= 1'b0;
    end else if(N4798) begin
      content_q[810] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[809] <= 1'b0;
    end else if(N4798) begin
      content_q[809] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[808] <= 1'b0;
    end else if(N4798) begin
      content_q[808] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[807] <= 1'b0;
    end else if(N4798) begin
      content_q[807] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[806] <= 1'b0;
    end else if(N4798) begin
      content_q[806] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[805] <= 1'b0;
    end else if(N4798) begin
      content_q[805] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[804] <= 1'b0;
    end else if(N4798) begin
      content_q[804] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[803] <= 1'b0;
    end else if(N4798) begin
      content_q[803] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[802] <= 1'b0;
    end else if(N4798) begin
      content_q[802] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[801] <= 1'b0;
    end else if(N4798) begin
      content_q[801] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[800] <= 1'b0;
    end else if(N4798) begin
      content_q[800] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[799] <= 1'b0;
    end else if(N4798) begin
      content_q[799] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[798] <= 1'b0;
    end else if(N4798) begin
      content_q[798] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[797] <= 1'b0;
    end else if(N4798) begin
      content_q[797] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[796] <= 1'b0;
    end else if(N4798) begin
      content_q[796] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[795] <= 1'b0;
    end else if(N4798) begin
      content_q[795] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[794] <= 1'b0;
    end else if(N4798) begin
      content_q[794] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[793] <= 1'b0;
    end else if(N4798) begin
      content_q[793] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[792] <= 1'b0;
    end else if(N4798) begin
      content_q[792] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[791] <= 1'b0;
    end else if(N4798) begin
      content_q[791] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[790] <= 1'b0;
    end else if(N4798) begin
      content_q[790] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[789] <= 1'b0;
    end else if(N4798) begin
      content_q[789] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[788] <= 1'b0;
    end else if(N4798) begin
      content_q[788] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[787] <= 1'b0;
    end else if(N4798) begin
      content_q[787] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[786] <= 1'b0;
    end else if(N4798) begin
      content_q[786] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[785] <= 1'b0;
    end else if(N4798) begin
      content_q[785] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[784] <= 1'b0;
    end else if(N4798) begin
      content_q[784] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[783] <= 1'b0;
    end else if(N4798) begin
      content_q[783] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[782] <= 1'b0;
    end else if(N4798) begin
      content_q[782] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[781] <= 1'b0;
    end else if(N4798) begin
      content_q[781] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[780] <= 1'b0;
    end else if(N4798) begin
      content_q[780] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[779] <= 1'b0;
    end else if(N4798) begin
      content_q[779] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[778] <= 1'b0;
    end else if(N4798) begin
      content_q[778] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[777] <= 1'b0;
    end else if(N4798) begin
      content_q[777] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[776] <= 1'b0;
    end else if(N4798) begin
      content_q[776] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[775] <= 1'b0;
    end else if(N4798) begin
      content_q[775] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[774] <= 1'b0;
    end else if(N4798) begin
      content_q[774] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[773] <= 1'b0;
    end else if(N4798) begin
      content_q[773] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[772] <= 1'b0;
    end else if(N4798) begin
      content_q[772] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[771] <= 1'b0;
    end else if(N4798) begin
      content_q[771] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[770] <= 1'b0;
    end else if(N4798) begin
      content_q[770] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[769] <= 1'b0;
    end else if(N4798) begin
      content_q[769] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[768] <= 1'b0;
    end else if(N4798) begin
      content_q[768] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[767] <= 1'b0;
    end else if(N4803) begin
      content_q[767] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[766] <= 1'b0;
    end else if(N4803) begin
      content_q[766] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[765] <= 1'b0;
    end else if(N4803) begin
      content_q[765] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[764] <= 1'b0;
    end else if(N4803) begin
      content_q[764] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[763] <= 1'b0;
    end else if(N4803) begin
      content_q[763] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[762] <= 1'b0;
    end else if(N4803) begin
      content_q[762] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[761] <= 1'b0;
    end else if(N4803) begin
      content_q[761] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[760] <= 1'b0;
    end else if(N4803) begin
      content_q[760] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[759] <= 1'b0;
    end else if(N4803) begin
      content_q[759] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[758] <= 1'b0;
    end else if(N4803) begin
      content_q[758] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[757] <= 1'b0;
    end else if(N4803) begin
      content_q[757] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[756] <= 1'b0;
    end else if(N4803) begin
      content_q[756] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[755] <= 1'b0;
    end else if(N4803) begin
      content_q[755] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[754] <= 1'b0;
    end else if(N4803) begin
      content_q[754] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[753] <= 1'b0;
    end else if(N4803) begin
      content_q[753] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[752] <= 1'b0;
    end else if(N4803) begin
      content_q[752] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[751] <= 1'b0;
    end else if(N4803) begin
      content_q[751] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[750] <= 1'b0;
    end else if(N4803) begin
      content_q[750] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[749] <= 1'b0;
    end else if(N4803) begin
      content_q[749] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[748] <= 1'b0;
    end else if(N4803) begin
      content_q[748] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[747] <= 1'b0;
    end else if(N4803) begin
      content_q[747] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[746] <= 1'b0;
    end else if(N4803) begin
      content_q[746] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[745] <= 1'b0;
    end else if(N4803) begin
      content_q[745] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[744] <= 1'b0;
    end else if(N4803) begin
      content_q[744] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[743] <= 1'b0;
    end else if(N4803) begin
      content_q[743] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[742] <= 1'b0;
    end else if(N4803) begin
      content_q[742] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[741] <= 1'b0;
    end else if(N4803) begin
      content_q[741] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[740] <= 1'b0;
    end else if(N4803) begin
      content_q[740] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[739] <= 1'b0;
    end else if(N4803) begin
      content_q[739] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[738] <= 1'b0;
    end else if(N4803) begin
      content_q[738] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[737] <= 1'b0;
    end else if(N4803) begin
      content_q[737] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[736] <= 1'b0;
    end else if(N4803) begin
      content_q[736] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[735] <= 1'b0;
    end else if(N4803) begin
      content_q[735] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[734] <= 1'b0;
    end else if(N4803) begin
      content_q[734] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[733] <= 1'b0;
    end else if(N4803) begin
      content_q[733] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[732] <= 1'b0;
    end else if(N4803) begin
      content_q[732] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[731] <= 1'b0;
    end else if(N4803) begin
      content_q[731] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[730] <= 1'b0;
    end else if(N4803) begin
      content_q[730] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[729] <= 1'b0;
    end else if(N4803) begin
      content_q[729] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[728] <= 1'b0;
    end else if(N4803) begin
      content_q[728] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[727] <= 1'b0;
    end else if(N4803) begin
      content_q[727] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[726] <= 1'b0;
    end else if(N4803) begin
      content_q[726] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[725] <= 1'b0;
    end else if(N4803) begin
      content_q[725] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[724] <= 1'b0;
    end else if(N4803) begin
      content_q[724] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[723] <= 1'b0;
    end else if(N4803) begin
      content_q[723] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[722] <= 1'b0;
    end else if(N4803) begin
      content_q[722] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[721] <= 1'b0;
    end else if(N4803) begin
      content_q[721] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[720] <= 1'b0;
    end else if(N4803) begin
      content_q[720] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[719] <= 1'b0;
    end else if(N4803) begin
      content_q[719] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[718] <= 1'b0;
    end else if(N4803) begin
      content_q[718] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[717] <= 1'b0;
    end else if(N4803) begin
      content_q[717] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[716] <= 1'b0;
    end else if(N4803) begin
      content_q[716] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[715] <= 1'b0;
    end else if(N4803) begin
      content_q[715] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[714] <= 1'b0;
    end else if(N4803) begin
      content_q[714] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[713] <= 1'b0;
    end else if(N4803) begin
      content_q[713] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[712] <= 1'b0;
    end else if(N4803) begin
      content_q[712] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[711] <= 1'b0;
    end else if(N4803) begin
      content_q[711] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[710] <= 1'b0;
    end else if(N4803) begin
      content_q[710] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[709] <= 1'b0;
    end else if(N4803) begin
      content_q[709] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[708] <= 1'b0;
    end else if(N4803) begin
      content_q[708] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[707] <= 1'b0;
    end else if(N4803) begin
      content_q[707] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[706] <= 1'b0;
    end else if(N4803) begin
      content_q[706] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[705] <= 1'b0;
    end else if(N4803) begin
      content_q[705] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[704] <= 1'b0;
    end else if(N4803) begin
      content_q[704] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[703] <= 1'b0;
    end else if(N4808) begin
      content_q[703] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[702] <= 1'b0;
    end else if(N4808) begin
      content_q[702] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[701] <= 1'b0;
    end else if(N4808) begin
      content_q[701] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[700] <= 1'b0;
    end else if(N4808) begin
      content_q[700] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[699] <= 1'b0;
    end else if(N4808) begin
      content_q[699] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[698] <= 1'b0;
    end else if(N4808) begin
      content_q[698] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[697] <= 1'b0;
    end else if(N4808) begin
      content_q[697] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[696] <= 1'b0;
    end else if(N4808) begin
      content_q[696] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[695] <= 1'b0;
    end else if(N4808) begin
      content_q[695] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[694] <= 1'b0;
    end else if(N4808) begin
      content_q[694] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[693] <= 1'b0;
    end else if(N4808) begin
      content_q[693] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[692] <= 1'b0;
    end else if(N4808) begin
      content_q[692] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[691] <= 1'b0;
    end else if(N4808) begin
      content_q[691] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[690] <= 1'b0;
    end else if(N4808) begin
      content_q[690] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[689] <= 1'b0;
    end else if(N4808) begin
      content_q[689] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[688] <= 1'b0;
    end else if(N4808) begin
      content_q[688] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[687] <= 1'b0;
    end else if(N4808) begin
      content_q[687] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[686] <= 1'b0;
    end else if(N4808) begin
      content_q[686] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[685] <= 1'b0;
    end else if(N4808) begin
      content_q[685] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[684] <= 1'b0;
    end else if(N4808) begin
      content_q[684] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[683] <= 1'b0;
    end else if(N4808) begin
      content_q[683] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[682] <= 1'b0;
    end else if(N4808) begin
      content_q[682] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[681] <= 1'b0;
    end else if(N4808) begin
      content_q[681] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[680] <= 1'b0;
    end else if(N4808) begin
      content_q[680] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[679] <= 1'b0;
    end else if(N4808) begin
      content_q[679] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[678] <= 1'b0;
    end else if(N4808) begin
      content_q[678] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[677] <= 1'b0;
    end else if(N4808) begin
      content_q[677] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[676] <= 1'b0;
    end else if(N4808) begin
      content_q[676] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[675] <= 1'b0;
    end else if(N4808) begin
      content_q[675] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[674] <= 1'b0;
    end else if(N4808) begin
      content_q[674] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[673] <= 1'b0;
    end else if(N4808) begin
      content_q[673] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[672] <= 1'b0;
    end else if(N4808) begin
      content_q[672] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[671] <= 1'b0;
    end else if(N4808) begin
      content_q[671] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[670] <= 1'b0;
    end else if(N4808) begin
      content_q[670] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[669] <= 1'b0;
    end else if(N4808) begin
      content_q[669] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[668] <= 1'b0;
    end else if(N4808) begin
      content_q[668] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[667] <= 1'b0;
    end else if(N4808) begin
      content_q[667] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[666] <= 1'b0;
    end else if(N4808) begin
      content_q[666] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[665] <= 1'b0;
    end else if(N4808) begin
      content_q[665] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[664] <= 1'b0;
    end else if(N4808) begin
      content_q[664] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[663] <= 1'b0;
    end else if(N4808) begin
      content_q[663] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[662] <= 1'b0;
    end else if(N4808) begin
      content_q[662] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[661] <= 1'b0;
    end else if(N4808) begin
      content_q[661] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[660] <= 1'b0;
    end else if(N4808) begin
      content_q[660] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[659] <= 1'b0;
    end else if(N4808) begin
      content_q[659] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[658] <= 1'b0;
    end else if(N4808) begin
      content_q[658] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[657] <= 1'b0;
    end else if(N4808) begin
      content_q[657] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[656] <= 1'b0;
    end else if(N4808) begin
      content_q[656] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[655] <= 1'b0;
    end else if(N4808) begin
      content_q[655] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[654] <= 1'b0;
    end else if(N4808) begin
      content_q[654] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[653] <= 1'b0;
    end else if(N4808) begin
      content_q[653] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[652] <= 1'b0;
    end else if(N4808) begin
      content_q[652] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[651] <= 1'b0;
    end else if(N4808) begin
      content_q[651] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[650] <= 1'b0;
    end else if(N4808) begin
      content_q[650] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[649] <= 1'b0;
    end else if(N4808) begin
      content_q[649] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[648] <= 1'b0;
    end else if(N4808) begin
      content_q[648] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[647] <= 1'b0;
    end else if(N4808) begin
      content_q[647] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[646] <= 1'b0;
    end else if(N4808) begin
      content_q[646] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[645] <= 1'b0;
    end else if(N4808) begin
      content_q[645] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[644] <= 1'b0;
    end else if(N4808) begin
      content_q[644] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[643] <= 1'b0;
    end else if(N4808) begin
      content_q[643] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[642] <= 1'b0;
    end else if(N4808) begin
      content_q[642] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[641] <= 1'b0;
    end else if(N4808) begin
      content_q[641] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[640] <= 1'b0;
    end else if(N4808) begin
      content_q[640] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[639] <= 1'b0;
    end else if(N4813) begin
      content_q[639] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[638] <= 1'b0;
    end else if(N4813) begin
      content_q[638] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[637] <= 1'b0;
    end else if(N4813) begin
      content_q[637] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[636] <= 1'b0;
    end else if(N4813) begin
      content_q[636] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[635] <= 1'b0;
    end else if(N4813) begin
      content_q[635] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[634] <= 1'b0;
    end else if(N4813) begin
      content_q[634] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[633] <= 1'b0;
    end else if(N4813) begin
      content_q[633] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[632] <= 1'b0;
    end else if(N4813) begin
      content_q[632] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[631] <= 1'b0;
    end else if(N4813) begin
      content_q[631] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[630] <= 1'b0;
    end else if(N4813) begin
      content_q[630] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[629] <= 1'b0;
    end else if(N4813) begin
      content_q[629] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[628] <= 1'b0;
    end else if(N4813) begin
      content_q[628] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[627] <= 1'b0;
    end else if(N4813) begin
      content_q[627] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[626] <= 1'b0;
    end else if(N4813) begin
      content_q[626] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[625] <= 1'b0;
    end else if(N4813) begin
      content_q[625] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[624] <= 1'b0;
    end else if(N4813) begin
      content_q[624] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[623] <= 1'b0;
    end else if(N4813) begin
      content_q[623] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[622] <= 1'b0;
    end else if(N4813) begin
      content_q[622] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[621] <= 1'b0;
    end else if(N4813) begin
      content_q[621] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[620] <= 1'b0;
    end else if(N4813) begin
      content_q[620] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[619] <= 1'b0;
    end else if(N4813) begin
      content_q[619] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[618] <= 1'b0;
    end else if(N4813) begin
      content_q[618] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[617] <= 1'b0;
    end else if(N4813) begin
      content_q[617] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[616] <= 1'b0;
    end else if(N4813) begin
      content_q[616] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[615] <= 1'b0;
    end else if(N4813) begin
      content_q[615] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[614] <= 1'b0;
    end else if(N4813) begin
      content_q[614] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[613] <= 1'b0;
    end else if(N4813) begin
      content_q[613] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[612] <= 1'b0;
    end else if(N4813) begin
      content_q[612] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[611] <= 1'b0;
    end else if(N4813) begin
      content_q[611] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[610] <= 1'b0;
    end else if(N4813) begin
      content_q[610] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[609] <= 1'b0;
    end else if(N4813) begin
      content_q[609] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[608] <= 1'b0;
    end else if(N4813) begin
      content_q[608] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[607] <= 1'b0;
    end else if(N4813) begin
      content_q[607] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[606] <= 1'b0;
    end else if(N4813) begin
      content_q[606] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[605] <= 1'b0;
    end else if(N4813) begin
      content_q[605] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[604] <= 1'b0;
    end else if(N4813) begin
      content_q[604] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[603] <= 1'b0;
    end else if(N4813) begin
      content_q[603] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[602] <= 1'b0;
    end else if(N4813) begin
      content_q[602] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[601] <= 1'b0;
    end else if(N4813) begin
      content_q[601] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[600] <= 1'b0;
    end else if(N4813) begin
      content_q[600] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[599] <= 1'b0;
    end else if(N4813) begin
      content_q[599] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[598] <= 1'b0;
    end else if(N4813) begin
      content_q[598] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[597] <= 1'b0;
    end else if(N4813) begin
      content_q[597] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[596] <= 1'b0;
    end else if(N4813) begin
      content_q[596] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[595] <= 1'b0;
    end else if(N4813) begin
      content_q[595] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[594] <= 1'b0;
    end else if(N4813) begin
      content_q[594] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[593] <= 1'b0;
    end else if(N4813) begin
      content_q[593] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[592] <= 1'b0;
    end else if(N4813) begin
      content_q[592] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[591] <= 1'b0;
    end else if(N4813) begin
      content_q[591] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[590] <= 1'b0;
    end else if(N4813) begin
      content_q[590] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[589] <= 1'b0;
    end else if(N4813) begin
      content_q[589] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[588] <= 1'b0;
    end else if(N4813) begin
      content_q[588] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[587] <= 1'b0;
    end else if(N4813) begin
      content_q[587] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[586] <= 1'b0;
    end else if(N4813) begin
      content_q[586] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[585] <= 1'b0;
    end else if(N4813) begin
      content_q[585] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[584] <= 1'b0;
    end else if(N4813) begin
      content_q[584] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[583] <= 1'b0;
    end else if(N4813) begin
      content_q[583] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[582] <= 1'b0;
    end else if(N4813) begin
      content_q[582] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[581] <= 1'b0;
    end else if(N4813) begin
      content_q[581] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[580] <= 1'b0;
    end else if(N4813) begin
      content_q[580] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[579] <= 1'b0;
    end else if(N4813) begin
      content_q[579] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[578] <= 1'b0;
    end else if(N4813) begin
      content_q[578] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[577] <= 1'b0;
    end else if(N4813) begin
      content_q[577] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[576] <= 1'b0;
    end else if(N4813) begin
      content_q[576] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[575] <= 1'b0;
    end else if(N4818) begin
      content_q[575] <= update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[574] <= 1'b0;
    end else if(N4818) begin
      content_q[574] <= update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[573] <= 1'b0;
    end else if(N4818) begin
      content_q[573] <= update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[572] <= 1'b0;
    end else if(N4818) begin
      content_q[572] <= update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[571] <= 1'b0;
    end else if(N4818) begin
      content_q[571] <= update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[570] <= 1'b0;
    end else if(N4818) begin
      content_q[570] <= update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[569] <= 1'b0;
    end else if(N4818) begin
      content_q[569] <= update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[568] <= 1'b0;
    end else if(N4818) begin
      content_q[568] <= update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[567] <= 1'b0;
    end else if(N4818) begin
      content_q[567] <= update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[566] <= 1'b0;
    end else if(N4818) begin
      content_q[566] <= update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[565] <= 1'b0;
    end else if(N4818) begin
      content_q[565] <= update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[564] <= 1'b0;
    end else if(N4818) begin
      content_q[564] <= update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[563] <= 1'b0;
    end else if(N4818) begin
      content_q[563] <= update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[562] <= 1'b0;
    end else if(N4818) begin
      content_q[562] <= update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[561] <= 1'b0;
    end else if(N4818) begin
      content_q[561] <= update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[560] <= 1'b0;
    end else if(N4818) begin
      content_q[560] <= update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[559] <= 1'b0;
    end else if(N4818) begin
      content_q[559] <= update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[558] <= 1'b0;
    end else if(N4818) begin
      content_q[558] <= update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[557] <= 1'b0;
    end else if(N4818) begin
      content_q[557] <= update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[556] <= 1'b0;
    end else if(N4818) begin
      content_q[556] <= update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[555] <= 1'b0;
    end else if(N4818) begin
      content_q[555] <= update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[554] <= 1'b0;
    end else if(N4818) begin
      content_q[554] <= update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[553] <= 1'b0;
    end else if(N4818) begin
      content_q[553] <= update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[552] <= 1'b0;
    end else if(N4818) begin
      content_q[552] <= update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[551] <= 1'b0;
    end else if(N4818) begin
      content_q[551] <= update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[550] <= 1'b0;
    end else if(N4818) begin
      content_q[550] <= update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[549] <= 1'b0;
    end else if(N4818) begin
      content_q[549] <= update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[548] <= 1'b0;
    end else if(N4818) begin
      content_q[548] <= update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[547] <= 1'b0;
    end else if(N4818) begin
      content_q[547] <= update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[546] <= 1'b0;
    end else if(N4818) begin
      content_q[546] <= update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[545] <= 1'b0;
    end else if(N4818) begin
      content_q[545] <= update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[544] <= 1'b0;
    end else if(N4818) begin
      content_q[544] <= update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[543] <= 1'b0;
    end else if(N4818) begin
      content_q[543] <= update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[542] <= 1'b0;
    end else if(N4818) begin
      content_q[542] <= update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[541] <= 1'b0;
    end else if(N4818) begin
      content_q[541] <= update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[540] <= 1'b0;
    end else if(N4818) begin
      content_q[540] <= update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[539] <= 1'b0;
    end else if(N4818) begin
      content_q[539] <= update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[538] <= 1'b0;
    end else if(N4818) begin
      content_q[538] <= update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[537] <= 1'b0;
    end else if(N4818) begin
      content_q[537] <= update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[536] <= 1'b0;
    end else if(N4818) begin
      content_q[536] <= update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[535] <= 1'b0;
    end else if(N4818) begin
      content_q[535] <= update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[534] <= 1'b0;
    end else if(N4818) begin
      content_q[534] <= update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[533] <= 1'b0;
    end else if(N4818) begin
      content_q[533] <= update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[532] <= 1'b0;
    end else if(N4818) begin
      content_q[532] <= update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[531] <= 1'b0;
    end else if(N4818) begin
      content_q[531] <= update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[530] <= 1'b0;
    end else if(N4818) begin
      content_q[530] <= update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[529] <= 1'b0;
    end else if(N4818) begin
      content_q[529] <= update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[528] <= 1'b0;
    end else if(N4818) begin
      content_q[528] <= update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[527] <= 1'b0;
    end else if(N4818) begin
      content_q[527] <= update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[526] <= 1'b0;
    end else if(N4818) begin
      content_q[526] <= update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[525] <= 1'b0;
    end else if(N4818) begin
      content_q[525] <= update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[524] <= 1'b0;
    end else if(N4818) begin
      content_q[524] <= update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[523] <= 1'b0;
    end else if(N4818) begin
      content_q[523] <= update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[522] <= 1'b0;
    end else if(N4818) begin
      content_q[522] <= update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[521] <= 1'b0;
    end else if(N4818) begin
      content_q[521] <= update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[520] <= 1'b0;
    end else if(N4818) begin
      content_q[520] <= update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[519] <= 1'b0;
    end else if(N4818) begin
      content_q[519] <= update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[518] <= 1'b0;
    end else if(N4818) begin
      content_q[518] <= update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[517] <= 1'b0;
    end else if(N4818) begin
      content_q[517] <= update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[516] <= 1'b0;
    end else if(N4818) begin
      content_q[516] <= update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[515] <= 1'b0;
    end else if(N4818) begin
      content_q[515] <= update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[514] <= 1'b0;
    end else if(N4818) begin
      content_q[514] <= update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[513] <= 1'b0;
    end else if(N4818) begin
      content_q[513] <= update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[512] <= 1'b0;
    end else if(N4818) begin
      content_q[512] <= update_i[0];
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[511] <= 1'b0;
    end else if(N4650) begin
      content_q[511] <= content_n_7__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[510] <= 1'b0;
    end else if(N4650) begin
      content_q[510] <= content_n_7__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[509] <= 1'b0;
    end else if(N4650) begin
      content_q[509] <= content_n_7__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[508] <= 1'b0;
    end else if(N4650) begin
      content_q[508] <= content_n_7__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[507] <= 1'b0;
    end else if(N4650) begin
      content_q[507] <= content_n_7__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[506] <= 1'b0;
    end else if(N4650) begin
      content_q[506] <= content_n_7__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[505] <= 1'b0;
    end else if(N4650) begin
      content_q[505] <= content_n_7__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[504] <= 1'b0;
    end else if(N4650) begin
      content_q[504] <= content_n_7__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[503] <= 1'b0;
    end else if(N4650) begin
      content_q[503] <= content_n_7__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[502] <= 1'b0;
    end else if(N4650) begin
      content_q[502] <= content_n_7__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[501] <= 1'b0;
    end else if(N4650) begin
      content_q[501] <= content_n_7__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[500] <= 1'b0;
    end else if(N4650) begin
      content_q[500] <= content_n_7__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[499] <= 1'b0;
    end else if(N4650) begin
      content_q[499] <= content_n_7__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[498] <= 1'b0;
    end else if(N4650) begin
      content_q[498] <= content_n_7__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[497] <= 1'b0;
    end else if(N4650) begin
      content_q[497] <= content_n_7__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[496] <= 1'b0;
    end else if(N4650) begin
      content_q[496] <= content_n_7__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[495] <= 1'b0;
    end else if(N4650) begin
      content_q[495] <= content_n_7__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[494] <= 1'b0;
    end else if(N4650) begin
      content_q[494] <= content_n_7__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[493] <= 1'b0;
    end else if(N4650) begin
      content_q[493] <= content_n_7__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[492] <= 1'b0;
    end else if(N4650) begin
      content_q[492] <= content_n_7__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[491] <= 1'b0;
    end else if(N4650) begin
      content_q[491] <= content_n_7__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[490] <= 1'b0;
    end else if(N4650) begin
      content_q[490] <= content_n_7__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[489] <= 1'b0;
    end else if(N4650) begin
      content_q[489] <= content_n_7__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[488] <= 1'b0;
    end else if(N4650) begin
      content_q[488] <= content_n_7__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[487] <= 1'b0;
    end else if(N4650) begin
      content_q[487] <= content_n_7__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[486] <= 1'b0;
    end else if(N4650) begin
      content_q[486] <= content_n_7__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[485] <= 1'b0;
    end else if(N4650) begin
      content_q[485] <= content_n_7__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[484] <= 1'b0;
    end else if(N4650) begin
      content_q[484] <= content_n_7__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[483] <= 1'b0;
    end else if(N4650) begin
      content_q[483] <= content_n_7__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[482] <= 1'b0;
    end else if(N4650) begin
      content_q[482] <= content_n_7__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[481] <= 1'b0;
    end else if(N4650) begin
      content_q[481] <= content_n_7__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[480] <= 1'b0;
    end else if(N4650) begin
      content_q[480] <= content_n_7__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[479] <= 1'b0;
    end else if(N4650) begin
      content_q[479] <= content_n_7__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[478] <= 1'b0;
    end else if(N4650) begin
      content_q[478] <= content_n_7__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[477] <= 1'b0;
    end else if(N4650) begin
      content_q[477] <= content_n_7__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[476] <= 1'b0;
    end else if(N4650) begin
      content_q[476] <= content_n_7__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[475] <= 1'b0;
    end else if(N4650) begin
      content_q[475] <= content_n_7__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[474] <= 1'b0;
    end else if(N4650) begin
      content_q[474] <= content_n_7__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[473] <= 1'b0;
    end else if(N4650) begin
      content_q[473] <= content_n_7__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[472] <= 1'b0;
    end else if(N4650) begin
      content_q[472] <= content_n_7__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[471] <= 1'b0;
    end else if(N4650) begin
      content_q[471] <= content_n_7__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[470] <= 1'b0;
    end else if(N4650) begin
      content_q[470] <= content_n_7__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[469] <= 1'b0;
    end else if(N4650) begin
      content_q[469] <= content_n_7__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[468] <= 1'b0;
    end else if(N4650) begin
      content_q[468] <= content_n_7__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[467] <= 1'b0;
    end else if(N4650) begin
      content_q[467] <= content_n_7__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[466] <= 1'b0;
    end else if(N4650) begin
      content_q[466] <= content_n_7__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[465] <= 1'b0;
    end else if(N4650) begin
      content_q[465] <= content_n_7__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[464] <= 1'b0;
    end else if(N4650) begin
      content_q[464] <= content_n_7__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[463] <= 1'b0;
    end else if(N4650) begin
      content_q[463] <= content_n_7__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[462] <= 1'b0;
    end else if(N4650) begin
      content_q[462] <= content_n_7__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[461] <= 1'b0;
    end else if(N4650) begin
      content_q[461] <= content_n_7__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[460] <= 1'b0;
    end else if(N4650) begin
      content_q[460] <= content_n_7__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[459] <= 1'b0;
    end else if(N4650) begin
      content_q[459] <= content_n_7__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[458] <= 1'b0;
    end else if(N4650) begin
      content_q[458] <= content_n_7__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[457] <= 1'b0;
    end else if(N4650) begin
      content_q[457] <= content_n_7__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[456] <= 1'b0;
    end else if(N4650) begin
      content_q[456] <= content_n_7__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[455] <= 1'b0;
    end else if(N4650) begin
      content_q[455] <= content_n_7__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[454] <= 1'b0;
    end else if(N4650) begin
      content_q[454] <= content_n_7__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[453] <= 1'b0;
    end else if(N4650) begin
      content_q[453] <= content_n_7__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[452] <= 1'b0;
    end else if(N4650) begin
      content_q[452] <= content_n_7__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[451] <= 1'b0;
    end else if(N4650) begin
      content_q[451] <= content_n_7__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[450] <= 1'b0;
    end else if(N4650) begin
      content_q[450] <= content_n_7__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[449] <= 1'b0;
    end else if(N4650) begin
      content_q[449] <= content_n_7__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[448] <= 1'b0;
    end else if(N4650) begin
      content_q[448] <= content_n_7__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[447] <= 1'b0;
    end else if(N4650) begin
      content_q[447] <= content_n_6__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[446] <= 1'b0;
    end else if(N4650) begin
      content_q[446] <= content_n_6__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[445] <= 1'b0;
    end else if(N4650) begin
      content_q[445] <= content_n_6__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[444] <= 1'b0;
    end else if(N4650) begin
      content_q[444] <= content_n_6__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[443] <= 1'b0;
    end else if(N4650) begin
      content_q[443] <= content_n_6__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[442] <= 1'b0;
    end else if(N4650) begin
      content_q[442] <= content_n_6__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[441] <= 1'b0;
    end else if(N4650) begin
      content_q[441] <= content_n_6__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[440] <= 1'b0;
    end else if(N4650) begin
      content_q[440] <= content_n_6__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[439] <= 1'b0;
    end else if(N4650) begin
      content_q[439] <= content_n_6__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[438] <= 1'b0;
    end else if(N4650) begin
      content_q[438] <= content_n_6__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[437] <= 1'b0;
    end else if(N4650) begin
      content_q[437] <= content_n_6__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[436] <= 1'b0;
    end else if(N4650) begin
      content_q[436] <= content_n_6__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[435] <= 1'b0;
    end else if(N4650) begin
      content_q[435] <= content_n_6__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[434] <= 1'b0;
    end else if(N4650) begin
      content_q[434] <= content_n_6__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[433] <= 1'b0;
    end else if(N4650) begin
      content_q[433] <= content_n_6__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[432] <= 1'b0;
    end else if(N4650) begin
      content_q[432] <= content_n_6__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[431] <= 1'b0;
    end else if(N4650) begin
      content_q[431] <= content_n_6__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[430] <= 1'b0;
    end else if(N4650) begin
      content_q[430] <= content_n_6__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[429] <= 1'b0;
    end else if(N4650) begin
      content_q[429] <= content_n_6__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[428] <= 1'b0;
    end else if(N4650) begin
      content_q[428] <= content_n_6__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[427] <= 1'b0;
    end else if(N4650) begin
      content_q[427] <= content_n_6__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[426] <= 1'b0;
    end else if(N4650) begin
      content_q[426] <= content_n_6__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[425] <= 1'b0;
    end else if(N4650) begin
      content_q[425] <= content_n_6__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[424] <= 1'b0;
    end else if(N4650) begin
      content_q[424] <= content_n_6__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[423] <= 1'b0;
    end else if(N4650) begin
      content_q[423] <= content_n_6__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[422] <= 1'b0;
    end else if(N4650) begin
      content_q[422] <= content_n_6__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[421] <= 1'b0;
    end else if(N4650) begin
      content_q[421] <= content_n_6__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[420] <= 1'b0;
    end else if(N4650) begin
      content_q[420] <= content_n_6__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[419] <= 1'b0;
    end else if(N4650) begin
      content_q[419] <= content_n_6__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[418] <= 1'b0;
    end else if(N4650) begin
      content_q[418] <= content_n_6__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[417] <= 1'b0;
    end else if(N4650) begin
      content_q[417] <= content_n_6__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[416] <= 1'b0;
    end else if(N4650) begin
      content_q[416] <= content_n_6__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[415] <= 1'b0;
    end else if(N4650) begin
      content_q[415] <= content_n_6__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[414] <= 1'b0;
    end else if(N4650) begin
      content_q[414] <= content_n_6__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[413] <= 1'b0;
    end else if(N4650) begin
      content_q[413] <= content_n_6__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[412] <= 1'b0;
    end else if(N4650) begin
      content_q[412] <= content_n_6__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[411] <= 1'b0;
    end else if(N4650) begin
      content_q[411] <= content_n_6__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[410] <= 1'b0;
    end else if(N4650) begin
      content_q[410] <= content_n_6__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[409] <= 1'b0;
    end else if(N4650) begin
      content_q[409] <= content_n_6__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[408] <= 1'b0;
    end else if(N4650) begin
      content_q[408] <= content_n_6__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[407] <= 1'b0;
    end else if(N4650) begin
      content_q[407] <= content_n_6__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[406] <= 1'b0;
    end else if(N4650) begin
      content_q[406] <= content_n_6__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[405] <= 1'b0;
    end else if(N4650) begin
      content_q[405] <= content_n_6__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[404] <= 1'b0;
    end else if(N4650) begin
      content_q[404] <= content_n_6__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[403] <= 1'b0;
    end else if(N4650) begin
      content_q[403] <= content_n_6__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[402] <= 1'b0;
    end else if(N4650) begin
      content_q[402] <= content_n_6__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[401] <= 1'b0;
    end else if(N4650) begin
      content_q[401] <= content_n_6__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[400] <= 1'b0;
    end else if(N4650) begin
      content_q[400] <= content_n_6__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[399] <= 1'b0;
    end else if(N4650) begin
      content_q[399] <= content_n_6__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[398] <= 1'b0;
    end else if(N4650) begin
      content_q[398] <= content_n_6__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[397] <= 1'b0;
    end else if(N4650) begin
      content_q[397] <= content_n_6__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[396] <= 1'b0;
    end else if(N4650) begin
      content_q[396] <= content_n_6__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[395] <= 1'b0;
    end else if(N4650) begin
      content_q[395] <= content_n_6__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[394] <= 1'b0;
    end else if(N4650) begin
      content_q[394] <= content_n_6__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[393] <= 1'b0;
    end else if(N4650) begin
      content_q[393] <= content_n_6__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[392] <= 1'b0;
    end else if(N4650) begin
      content_q[392] <= content_n_6__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[391] <= 1'b0;
    end else if(N4650) begin
      content_q[391] <= content_n_6__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[390] <= 1'b0;
    end else if(N4650) begin
      content_q[390] <= content_n_6__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[389] <= 1'b0;
    end else if(N4650) begin
      content_q[389] <= content_n_6__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[388] <= 1'b0;
    end else if(N4650) begin
      content_q[388] <= content_n_6__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[387] <= 1'b0;
    end else if(N4650) begin
      content_q[387] <= content_n_6__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[386] <= 1'b0;
    end else if(N4650) begin
      content_q[386] <= content_n_6__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[385] <= 1'b0;
    end else if(N4650) begin
      content_q[385] <= content_n_6__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[384] <= 1'b0;
    end else if(N4650) begin
      content_q[384] <= content_n_6__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[383] <= 1'b0;
    end else if(N4650) begin
      content_q[383] <= content_n_5__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[382] <= 1'b0;
    end else if(N4650) begin
      content_q[382] <= content_n_5__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[381] <= 1'b0;
    end else if(N4650) begin
      content_q[381] <= content_n_5__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[380] <= 1'b0;
    end else if(N4650) begin
      content_q[380] <= content_n_5__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[379] <= 1'b0;
    end else if(N4650) begin
      content_q[379] <= content_n_5__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[378] <= 1'b0;
    end else if(N4650) begin
      content_q[378] <= content_n_5__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[377] <= 1'b0;
    end else if(N4650) begin
      content_q[377] <= content_n_5__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[376] <= 1'b0;
    end else if(N4650) begin
      content_q[376] <= content_n_5__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[375] <= 1'b0;
    end else if(N4650) begin
      content_q[375] <= content_n_5__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[374] <= 1'b0;
    end else if(N4650) begin
      content_q[374] <= content_n_5__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[373] <= 1'b0;
    end else if(N4650) begin
      content_q[373] <= content_n_5__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[372] <= 1'b0;
    end else if(N4650) begin
      content_q[372] <= content_n_5__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[371] <= 1'b0;
    end else if(N4650) begin
      content_q[371] <= content_n_5__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[370] <= 1'b0;
    end else if(N4650) begin
      content_q[370] <= content_n_5__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[369] <= 1'b0;
    end else if(N4650) begin
      content_q[369] <= content_n_5__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[368] <= 1'b0;
    end else if(N4650) begin
      content_q[368] <= content_n_5__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[367] <= 1'b0;
    end else if(N4650) begin
      content_q[367] <= content_n_5__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[366] <= 1'b0;
    end else if(N4650) begin
      content_q[366] <= content_n_5__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[365] <= 1'b0;
    end else if(N4650) begin
      content_q[365] <= content_n_5__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[364] <= 1'b0;
    end else if(N4650) begin
      content_q[364] <= content_n_5__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[363] <= 1'b0;
    end else if(N4650) begin
      content_q[363] <= content_n_5__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[362] <= 1'b0;
    end else if(N4650) begin
      content_q[362] <= content_n_5__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[361] <= 1'b0;
    end else if(N4650) begin
      content_q[361] <= content_n_5__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[360] <= 1'b0;
    end else if(N4650) begin
      content_q[360] <= content_n_5__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[359] <= 1'b0;
    end else if(N4650) begin
      content_q[359] <= content_n_5__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[358] <= 1'b0;
    end else if(N4650) begin
      content_q[358] <= content_n_5__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[357] <= 1'b0;
    end else if(N4650) begin
      content_q[357] <= content_n_5__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[356] <= 1'b0;
    end else if(N4650) begin
      content_q[356] <= content_n_5__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[355] <= 1'b0;
    end else if(N4650) begin
      content_q[355] <= content_n_5__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[354] <= 1'b0;
    end else if(N4650) begin
      content_q[354] <= content_n_5__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[353] <= 1'b0;
    end else if(N4650) begin
      content_q[353] <= content_n_5__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[352] <= 1'b0;
    end else if(N4650) begin
      content_q[352] <= content_n_5__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[351] <= 1'b0;
    end else if(N4650) begin
      content_q[351] <= content_n_5__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[350] <= 1'b0;
    end else if(N4650) begin
      content_q[350] <= content_n_5__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[349] <= 1'b0;
    end else if(N4650) begin
      content_q[349] <= content_n_5__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[348] <= 1'b0;
    end else if(N4650) begin
      content_q[348] <= content_n_5__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[347] <= 1'b0;
    end else if(N4650) begin
      content_q[347] <= content_n_5__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[346] <= 1'b0;
    end else if(N4650) begin
      content_q[346] <= content_n_5__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[345] <= 1'b0;
    end else if(N4650) begin
      content_q[345] <= content_n_5__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[344] <= 1'b0;
    end else if(N4650) begin
      content_q[344] <= content_n_5__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[343] <= 1'b0;
    end else if(N4650) begin
      content_q[343] <= content_n_5__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[342] <= 1'b0;
    end else if(N4650) begin
      content_q[342] <= content_n_5__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[341] <= 1'b0;
    end else if(N4650) begin
      content_q[341] <= content_n_5__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[340] <= 1'b0;
    end else if(N4650) begin
      content_q[340] <= content_n_5__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[339] <= 1'b0;
    end else if(N4650) begin
      content_q[339] <= content_n_5__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[338] <= 1'b0;
    end else if(N4650) begin
      content_q[338] <= content_n_5__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[337] <= 1'b0;
    end else if(N4650) begin
      content_q[337] <= content_n_5__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[336] <= 1'b0;
    end else if(N4650) begin
      content_q[336] <= content_n_5__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[335] <= 1'b0;
    end else if(N4650) begin
      content_q[335] <= content_n_5__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[334] <= 1'b0;
    end else if(N4650) begin
      content_q[334] <= content_n_5__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[333] <= 1'b0;
    end else if(N4650) begin
      content_q[333] <= content_n_5__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[332] <= 1'b0;
    end else if(N4650) begin
      content_q[332] <= content_n_5__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[331] <= 1'b0;
    end else if(N4650) begin
      content_q[331] <= content_n_5__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[330] <= 1'b0;
    end else if(N4650) begin
      content_q[330] <= content_n_5__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[329] <= 1'b0;
    end else if(N4650) begin
      content_q[329] <= content_n_5__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[328] <= 1'b0;
    end else if(N4650) begin
      content_q[328] <= content_n_5__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[327] <= 1'b0;
    end else if(N4650) begin
      content_q[327] <= content_n_5__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[326] <= 1'b0;
    end else if(N4650) begin
      content_q[326] <= content_n_5__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[325] <= 1'b0;
    end else if(N4650) begin
      content_q[325] <= content_n_5__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[324] <= 1'b0;
    end else if(N4650) begin
      content_q[324] <= content_n_5__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[323] <= 1'b0;
    end else if(N4650) begin
      content_q[323] <= content_n_5__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[322] <= 1'b0;
    end else if(N4650) begin
      content_q[322] <= content_n_5__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[321] <= 1'b0;
    end else if(N4650) begin
      content_q[321] <= content_n_5__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[320] <= 1'b0;
    end else if(N4650) begin
      content_q[320] <= content_n_5__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[319] <= 1'b0;
    end else if(N4650) begin
      content_q[319] <= content_n_4__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[318] <= 1'b0;
    end else if(N4650) begin
      content_q[318] <= content_n_4__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[317] <= 1'b0;
    end else if(N4650) begin
      content_q[317] <= content_n_4__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[316] <= 1'b0;
    end else if(N4650) begin
      content_q[316] <= content_n_4__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[315] <= 1'b0;
    end else if(N4650) begin
      content_q[315] <= content_n_4__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[314] <= 1'b0;
    end else if(N4650) begin
      content_q[314] <= content_n_4__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[313] <= 1'b0;
    end else if(N4650) begin
      content_q[313] <= content_n_4__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[312] <= 1'b0;
    end else if(N4650) begin
      content_q[312] <= content_n_4__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[311] <= 1'b0;
    end else if(N4650) begin
      content_q[311] <= content_n_4__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[310] <= 1'b0;
    end else if(N4650) begin
      content_q[310] <= content_n_4__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[309] <= 1'b0;
    end else if(N4650) begin
      content_q[309] <= content_n_4__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[308] <= 1'b0;
    end else if(N4650) begin
      content_q[308] <= content_n_4__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[307] <= 1'b0;
    end else if(N4650) begin
      content_q[307] <= content_n_4__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[306] <= 1'b0;
    end else if(N4650) begin
      content_q[306] <= content_n_4__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[305] <= 1'b0;
    end else if(N4650) begin
      content_q[305] <= content_n_4__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[304] <= 1'b0;
    end else if(N4650) begin
      content_q[304] <= content_n_4__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[303] <= 1'b0;
    end else if(N4650) begin
      content_q[303] <= content_n_4__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[302] <= 1'b0;
    end else if(N4650) begin
      content_q[302] <= content_n_4__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[301] <= 1'b0;
    end else if(N4650) begin
      content_q[301] <= content_n_4__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[300] <= 1'b0;
    end else if(N4650) begin
      content_q[300] <= content_n_4__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[299] <= 1'b0;
    end else if(N4650) begin
      content_q[299] <= content_n_4__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[298] <= 1'b0;
    end else if(N4650) begin
      content_q[298] <= content_n_4__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[297] <= 1'b0;
    end else if(N4650) begin
      content_q[297] <= content_n_4__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[296] <= 1'b0;
    end else if(N4650) begin
      content_q[296] <= content_n_4__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[295] <= 1'b0;
    end else if(N4650) begin
      content_q[295] <= content_n_4__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[294] <= 1'b0;
    end else if(N4650) begin
      content_q[294] <= content_n_4__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[293] <= 1'b0;
    end else if(N4650) begin
      content_q[293] <= content_n_4__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[292] <= 1'b0;
    end else if(N4650) begin
      content_q[292] <= content_n_4__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[291] <= 1'b0;
    end else if(N4650) begin
      content_q[291] <= content_n_4__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[290] <= 1'b0;
    end else if(N4650) begin
      content_q[290] <= content_n_4__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[289] <= 1'b0;
    end else if(N4650) begin
      content_q[289] <= content_n_4__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[288] <= 1'b0;
    end else if(N4650) begin
      content_q[288] <= content_n_4__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[287] <= 1'b0;
    end else if(N4650) begin
      content_q[287] <= content_n_4__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[286] <= 1'b0;
    end else if(N4650) begin
      content_q[286] <= content_n_4__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[285] <= 1'b0;
    end else if(N4650) begin
      content_q[285] <= content_n_4__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[284] <= 1'b0;
    end else if(N4650) begin
      content_q[284] <= content_n_4__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[283] <= 1'b0;
    end else if(N4650) begin
      content_q[283] <= content_n_4__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[282] <= 1'b0;
    end else if(N4650) begin
      content_q[282] <= content_n_4__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[281] <= 1'b0;
    end else if(N4650) begin
      content_q[281] <= content_n_4__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[280] <= 1'b0;
    end else if(N4650) begin
      content_q[280] <= content_n_4__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[279] <= 1'b0;
    end else if(N4650) begin
      content_q[279] <= content_n_4__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[278] <= 1'b0;
    end else if(N4650) begin
      content_q[278] <= content_n_4__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[277] <= 1'b0;
    end else if(N4650) begin
      content_q[277] <= content_n_4__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[276] <= 1'b0;
    end else if(N4650) begin
      content_q[276] <= content_n_4__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[275] <= 1'b0;
    end else if(N4650) begin
      content_q[275] <= content_n_4__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[274] <= 1'b0;
    end else if(N4650) begin
      content_q[274] <= content_n_4__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[273] <= 1'b0;
    end else if(N4650) begin
      content_q[273] <= content_n_4__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[272] <= 1'b0;
    end else if(N4650) begin
      content_q[272] <= content_n_4__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[271] <= 1'b0;
    end else if(N4650) begin
      content_q[271] <= content_n_4__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[270] <= 1'b0;
    end else if(N4650) begin
      content_q[270] <= content_n_4__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[269] <= 1'b0;
    end else if(N4650) begin
      content_q[269] <= content_n_4__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[268] <= 1'b0;
    end else if(N4650) begin
      content_q[268] <= content_n_4__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[267] <= 1'b0;
    end else if(N4650) begin
      content_q[267] <= content_n_4__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[266] <= 1'b0;
    end else if(N4650) begin
      content_q[266] <= content_n_4__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[265] <= 1'b0;
    end else if(N4650) begin
      content_q[265] <= content_n_4__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[264] <= 1'b0;
    end else if(N4650) begin
      content_q[264] <= content_n_4__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[263] <= 1'b0;
    end else if(N4650) begin
      content_q[263] <= content_n_4__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[262] <= 1'b0;
    end else if(N4650) begin
      content_q[262] <= content_n_4__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[261] <= 1'b0;
    end else if(N4650) begin
      content_q[261] <= content_n_4__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[260] <= 1'b0;
    end else if(N4650) begin
      content_q[260] <= content_n_4__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[259] <= 1'b0;
    end else if(N4650) begin
      content_q[259] <= content_n_4__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[258] <= 1'b0;
    end else if(N4650) begin
      content_q[258] <= content_n_4__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[257] <= 1'b0;
    end else if(N4650) begin
      content_q[257] <= content_n_4__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[256] <= 1'b0;
    end else if(N4650) begin
      content_q[256] <= content_n_4__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[255] <= 1'b0;
    end else if(N4650) begin
      content_q[255] <= content_n_3__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[254] <= 1'b0;
    end else if(N4650) begin
      content_q[254] <= content_n_3__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[253] <= 1'b0;
    end else if(N4650) begin
      content_q[253] <= content_n_3__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[252] <= 1'b0;
    end else if(N4650) begin
      content_q[252] <= content_n_3__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[251] <= 1'b0;
    end else if(N4650) begin
      content_q[251] <= content_n_3__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[250] <= 1'b0;
    end else if(N4650) begin
      content_q[250] <= content_n_3__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[249] <= 1'b0;
    end else if(N4650) begin
      content_q[249] <= content_n_3__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[248] <= 1'b0;
    end else if(N4650) begin
      content_q[248] <= content_n_3__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[247] <= 1'b0;
    end else if(N4650) begin
      content_q[247] <= content_n_3__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[246] <= 1'b0;
    end else if(N4650) begin
      content_q[246] <= content_n_3__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[245] <= 1'b0;
    end else if(N4650) begin
      content_q[245] <= content_n_3__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[244] <= 1'b0;
    end else if(N4650) begin
      content_q[244] <= content_n_3__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[243] <= 1'b0;
    end else if(N4650) begin
      content_q[243] <= content_n_3__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[242] <= 1'b0;
    end else if(N4650) begin
      content_q[242] <= content_n_3__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[241] <= 1'b0;
    end else if(N4650) begin
      content_q[241] <= content_n_3__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[240] <= 1'b0;
    end else if(N4650) begin
      content_q[240] <= content_n_3__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[239] <= 1'b0;
    end else if(N4650) begin
      content_q[239] <= content_n_3__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[238] <= 1'b0;
    end else if(N4650) begin
      content_q[238] <= content_n_3__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[237] <= 1'b0;
    end else if(N4650) begin
      content_q[237] <= content_n_3__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[236] <= 1'b0;
    end else if(N4650) begin
      content_q[236] <= content_n_3__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[235] <= 1'b0;
    end else if(N4650) begin
      content_q[235] <= content_n_3__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[234] <= 1'b0;
    end else if(N4650) begin
      content_q[234] <= content_n_3__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[233] <= 1'b0;
    end else if(N4650) begin
      content_q[233] <= content_n_3__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[232] <= 1'b0;
    end else if(N4650) begin
      content_q[232] <= content_n_3__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[231] <= 1'b0;
    end else if(N4650) begin
      content_q[231] <= content_n_3__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[230] <= 1'b0;
    end else if(N4650) begin
      content_q[230] <= content_n_3__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[229] <= 1'b0;
    end else if(N4650) begin
      content_q[229] <= content_n_3__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[228] <= 1'b0;
    end else if(N4650) begin
      content_q[228] <= content_n_3__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[227] <= 1'b0;
    end else if(N4650) begin
      content_q[227] <= content_n_3__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[226] <= 1'b0;
    end else if(N4650) begin
      content_q[226] <= content_n_3__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[225] <= 1'b0;
    end else if(N4650) begin
      content_q[225] <= content_n_3__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[224] <= 1'b0;
    end else if(N4650) begin
      content_q[224] <= content_n_3__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[223] <= 1'b0;
    end else if(N4650) begin
      content_q[223] <= content_n_3__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[222] <= 1'b0;
    end else if(N4650) begin
      content_q[222] <= content_n_3__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[221] <= 1'b0;
    end else if(N4650) begin
      content_q[221] <= content_n_3__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[220] <= 1'b0;
    end else if(N4650) begin
      content_q[220] <= content_n_3__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[219] <= 1'b0;
    end else if(N4650) begin
      content_q[219] <= content_n_3__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[218] <= 1'b0;
    end else if(N4650) begin
      content_q[218] <= content_n_3__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[217] <= 1'b0;
    end else if(N4650) begin
      content_q[217] <= content_n_3__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[216] <= 1'b0;
    end else if(N4650) begin
      content_q[216] <= content_n_3__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[215] <= 1'b0;
    end else if(N4650) begin
      content_q[215] <= content_n_3__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[214] <= 1'b0;
    end else if(N4650) begin
      content_q[214] <= content_n_3__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[213] <= 1'b0;
    end else if(N4650) begin
      content_q[213] <= content_n_3__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[212] <= 1'b0;
    end else if(N4650) begin
      content_q[212] <= content_n_3__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[211] <= 1'b0;
    end else if(N4650) begin
      content_q[211] <= content_n_3__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[210] <= 1'b0;
    end else if(N4650) begin
      content_q[210] <= content_n_3__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[209] <= 1'b0;
    end else if(N4650) begin
      content_q[209] <= content_n_3__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[208] <= 1'b0;
    end else if(N4650) begin
      content_q[208] <= content_n_3__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[207] <= 1'b0;
    end else if(N4650) begin
      content_q[207] <= content_n_3__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[206] <= 1'b0;
    end else if(N4650) begin
      content_q[206] <= content_n_3__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[205] <= 1'b0;
    end else if(N4650) begin
      content_q[205] <= content_n_3__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[204] <= 1'b0;
    end else if(N4650) begin
      content_q[204] <= content_n_3__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[203] <= 1'b0;
    end else if(N4650) begin
      content_q[203] <= content_n_3__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[202] <= 1'b0;
    end else if(N4650) begin
      content_q[202] <= content_n_3__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[201] <= 1'b0;
    end else if(N4650) begin
      content_q[201] <= content_n_3__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[200] <= 1'b0;
    end else if(N4650) begin
      content_q[200] <= content_n_3__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[199] <= 1'b0;
    end else if(N4650) begin
      content_q[199] <= content_n_3__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[198] <= 1'b0;
    end else if(N4650) begin
      content_q[198] <= content_n_3__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[197] <= 1'b0;
    end else if(N4650) begin
      content_q[197] <= content_n_3__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[196] <= 1'b0;
    end else if(N4650) begin
      content_q[196] <= content_n_3__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[195] <= 1'b0;
    end else if(N4650) begin
      content_q[195] <= content_n_3__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[194] <= 1'b0;
    end else if(N4650) begin
      content_q[194] <= content_n_3__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[193] <= 1'b0;
    end else if(N4650) begin
      content_q[193] <= content_n_3__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[192] <= 1'b0;
    end else if(N4650) begin
      content_q[192] <= content_n_3__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[191] <= 1'b0;
    end else if(N4650) begin
      content_q[191] <= content_n_2__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[190] <= 1'b0;
    end else if(N4650) begin
      content_q[190] <= content_n_2__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[189] <= 1'b0;
    end else if(N4650) begin
      content_q[189] <= content_n_2__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[188] <= 1'b0;
    end else if(N4650) begin
      content_q[188] <= content_n_2__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[187] <= 1'b0;
    end else if(N4650) begin
      content_q[187] <= content_n_2__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[186] <= 1'b0;
    end else if(N4650) begin
      content_q[186] <= content_n_2__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[185] <= 1'b0;
    end else if(N4650) begin
      content_q[185] <= content_n_2__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[184] <= 1'b0;
    end else if(N4650) begin
      content_q[184] <= content_n_2__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[183] <= 1'b0;
    end else if(N4650) begin
      content_q[183] <= content_n_2__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[182] <= 1'b0;
    end else if(N4650) begin
      content_q[182] <= content_n_2__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[181] <= 1'b0;
    end else if(N4650) begin
      content_q[181] <= content_n_2__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[180] <= 1'b0;
    end else if(N4650) begin
      content_q[180] <= content_n_2__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[179] <= 1'b0;
    end else if(N4650) begin
      content_q[179] <= content_n_2__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[178] <= 1'b0;
    end else if(N4650) begin
      content_q[178] <= content_n_2__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[177] <= 1'b0;
    end else if(N4650) begin
      content_q[177] <= content_n_2__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[176] <= 1'b0;
    end else if(N4650) begin
      content_q[176] <= content_n_2__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[175] <= 1'b0;
    end else if(N4650) begin
      content_q[175] <= content_n_2__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[174] <= 1'b0;
    end else if(N4650) begin
      content_q[174] <= content_n_2__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[173] <= 1'b0;
    end else if(N4650) begin
      content_q[173] <= content_n_2__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[172] <= 1'b0;
    end else if(N4650) begin
      content_q[172] <= content_n_2__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[171] <= 1'b0;
    end else if(N4650) begin
      content_q[171] <= content_n_2__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[170] <= 1'b0;
    end else if(N4650) begin
      content_q[170] <= content_n_2__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[169] <= 1'b0;
    end else if(N4650) begin
      content_q[169] <= content_n_2__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[168] <= 1'b0;
    end else if(N4650) begin
      content_q[168] <= content_n_2__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[167] <= 1'b0;
    end else if(N4650) begin
      content_q[167] <= content_n_2__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[166] <= 1'b0;
    end else if(N4650) begin
      content_q[166] <= content_n_2__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[165] <= 1'b0;
    end else if(N4650) begin
      content_q[165] <= content_n_2__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[164] <= 1'b0;
    end else if(N4650) begin
      content_q[164] <= content_n_2__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[163] <= 1'b0;
    end else if(N4650) begin
      content_q[163] <= content_n_2__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[162] <= 1'b0;
    end else if(N4650) begin
      content_q[162] <= content_n_2__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[161] <= 1'b0;
    end else if(N4650) begin
      content_q[161] <= content_n_2__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[160] <= 1'b0;
    end else if(N4650) begin
      content_q[160] <= content_n_2__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[159] <= 1'b0;
    end else if(N4650) begin
      content_q[159] <= content_n_2__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[158] <= 1'b0;
    end else if(N4650) begin
      content_q[158] <= content_n_2__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[157] <= 1'b0;
    end else if(N4650) begin
      content_q[157] <= content_n_2__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[156] <= 1'b0;
    end else if(N4650) begin
      content_q[156] <= content_n_2__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[155] <= 1'b0;
    end else if(N4650) begin
      content_q[155] <= content_n_2__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[154] <= 1'b0;
    end else if(N4650) begin
      content_q[154] <= content_n_2__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[153] <= 1'b0;
    end else if(N4650) begin
      content_q[153] <= content_n_2__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[152] <= 1'b0;
    end else if(N4650) begin
      content_q[152] <= content_n_2__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[151] <= 1'b0;
    end else if(N4650) begin
      content_q[151] <= content_n_2__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[150] <= 1'b0;
    end else if(N4650) begin
      content_q[150] <= content_n_2__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[149] <= 1'b0;
    end else if(N4650) begin
      content_q[149] <= content_n_2__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[148] <= 1'b0;
    end else if(N4650) begin
      content_q[148] <= content_n_2__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[147] <= 1'b0;
    end else if(N4650) begin
      content_q[147] <= content_n_2__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[146] <= 1'b0;
    end else if(N4650) begin
      content_q[146] <= content_n_2__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[145] <= 1'b0;
    end else if(N4650) begin
      content_q[145] <= content_n_2__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[144] <= 1'b0;
    end else if(N4650) begin
      content_q[144] <= content_n_2__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[143] <= 1'b0;
    end else if(N4650) begin
      content_q[143] <= content_n_2__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[142] <= 1'b0;
    end else if(N4650) begin
      content_q[142] <= content_n_2__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[141] <= 1'b0;
    end else if(N4650) begin
      content_q[141] <= content_n_2__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[140] <= 1'b0;
    end else if(N4650) begin
      content_q[140] <= content_n_2__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[139] <= 1'b0;
    end else if(N4650) begin
      content_q[139] <= content_n_2__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[138] <= 1'b0;
    end else if(N4650) begin
      content_q[138] <= content_n_2__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[137] <= 1'b0;
    end else if(N4650) begin
      content_q[137] <= content_n_2__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[136] <= 1'b0;
    end else if(N4650) begin
      content_q[136] <= content_n_2__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[135] <= 1'b0;
    end else if(N4650) begin
      content_q[135] <= content_n_2__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[134] <= 1'b0;
    end else if(N4650) begin
      content_q[134] <= content_n_2__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[133] <= 1'b0;
    end else if(N4650) begin
      content_q[133] <= content_n_2__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[132] <= 1'b0;
    end else if(N4650) begin
      content_q[132] <= content_n_2__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[131] <= 1'b0;
    end else if(N4650) begin
      content_q[131] <= content_n_2__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[130] <= 1'b0;
    end else if(N4650) begin
      content_q[130] <= content_n_2__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[129] <= 1'b0;
    end else if(N4650) begin
      content_q[129] <= content_n_2__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[128] <= 1'b0;
    end else if(N4650) begin
      content_q[128] <= content_n_2__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[127] <= 1'b0;
    end else if(N4650) begin
      content_q[127] <= content_n_1__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[126] <= 1'b0;
    end else if(N4650) begin
      content_q[126] <= content_n_1__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[125] <= 1'b0;
    end else if(N4650) begin
      content_q[125] <= content_n_1__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[124] <= 1'b0;
    end else if(N4650) begin
      content_q[124] <= content_n_1__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[123] <= 1'b0;
    end else if(N4650) begin
      content_q[123] <= content_n_1__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[122] <= 1'b0;
    end else if(N4650) begin
      content_q[122] <= content_n_1__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[121] <= 1'b0;
    end else if(N4650) begin
      content_q[121] <= content_n_1__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[120] <= 1'b0;
    end else if(N4650) begin
      content_q[120] <= content_n_1__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[119] <= 1'b0;
    end else if(N4650) begin
      content_q[119] <= content_n_1__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[118] <= 1'b0;
    end else if(N4650) begin
      content_q[118] <= content_n_1__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[117] <= 1'b0;
    end else if(N4650) begin
      content_q[117] <= content_n_1__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[116] <= 1'b0;
    end else if(N4650) begin
      content_q[116] <= content_n_1__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[115] <= 1'b0;
    end else if(N4650) begin
      content_q[115] <= content_n_1__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[114] <= 1'b0;
    end else if(N4650) begin
      content_q[114] <= content_n_1__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[113] <= 1'b0;
    end else if(N4650) begin
      content_q[113] <= content_n_1__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[112] <= 1'b0;
    end else if(N4650) begin
      content_q[112] <= content_n_1__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[111] <= 1'b0;
    end else if(N4650) begin
      content_q[111] <= content_n_1__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[110] <= 1'b0;
    end else if(N4650) begin
      content_q[110] <= content_n_1__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[109] <= 1'b0;
    end else if(N4650) begin
      content_q[109] <= content_n_1__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[108] <= 1'b0;
    end else if(N4650) begin
      content_q[108] <= content_n_1__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[107] <= 1'b0;
    end else if(N4650) begin
      content_q[107] <= content_n_1__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[106] <= 1'b0;
    end else if(N4650) begin
      content_q[106] <= content_n_1__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[105] <= 1'b0;
    end else if(N4650) begin
      content_q[105] <= content_n_1__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[104] <= 1'b0;
    end else if(N4650) begin
      content_q[104] <= content_n_1__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[103] <= 1'b0;
    end else if(N4650) begin
      content_q[103] <= content_n_1__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[102] <= 1'b0;
    end else if(N4650) begin
      content_q[102] <= content_n_1__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[101] <= 1'b0;
    end else if(N4650) begin
      content_q[101] <= content_n_1__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[100] <= 1'b0;
    end else if(N4650) begin
      content_q[100] <= content_n_1__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[99] <= 1'b0;
    end else if(N4650) begin
      content_q[99] <= content_n_1__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[98] <= 1'b0;
    end else if(N4650) begin
      content_q[98] <= content_n_1__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[97] <= 1'b0;
    end else if(N4650) begin
      content_q[97] <= content_n_1__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[96] <= 1'b0;
    end else if(N4650) begin
      content_q[96] <= content_n_1__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[95] <= 1'b0;
    end else if(N4650) begin
      content_q[95] <= content_n_1__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[94] <= 1'b0;
    end else if(N4650) begin
      content_q[94] <= content_n_1__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[93] <= 1'b0;
    end else if(N4650) begin
      content_q[93] <= content_n_1__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[92] <= 1'b0;
    end else if(N4650) begin
      content_q[92] <= content_n_1__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[91] <= 1'b0;
    end else if(N4650) begin
      content_q[91] <= content_n_1__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[90] <= 1'b0;
    end else if(N4650) begin
      content_q[90] <= content_n_1__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[89] <= 1'b0;
    end else if(N4650) begin
      content_q[89] <= content_n_1__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[88] <= 1'b0;
    end else if(N4650) begin
      content_q[88] <= content_n_1__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[87] <= 1'b0;
    end else if(N4650) begin
      content_q[87] <= content_n_1__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[86] <= 1'b0;
    end else if(N4650) begin
      content_q[86] <= content_n_1__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[85] <= 1'b0;
    end else if(N4650) begin
      content_q[85] <= content_n_1__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[84] <= 1'b0;
    end else if(N4650) begin
      content_q[84] <= content_n_1__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[83] <= 1'b0;
    end else if(N4650) begin
      content_q[83] <= content_n_1__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[82] <= 1'b0;
    end else if(N4650) begin
      content_q[82] <= content_n_1__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[81] <= 1'b0;
    end else if(N4650) begin
      content_q[81] <= content_n_1__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[80] <= 1'b0;
    end else if(N4650) begin
      content_q[80] <= content_n_1__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[79] <= 1'b0;
    end else if(N4650) begin
      content_q[79] <= content_n_1__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[78] <= 1'b0;
    end else if(N4650) begin
      content_q[78] <= content_n_1__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[77] <= 1'b0;
    end else if(N4650) begin
      content_q[77] <= content_n_1__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[76] <= 1'b0;
    end else if(N4650) begin
      content_q[76] <= content_n_1__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[75] <= 1'b0;
    end else if(N4650) begin
      content_q[75] <= content_n_1__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[74] <= 1'b0;
    end else if(N4650) begin
      content_q[74] <= content_n_1__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[73] <= 1'b0;
    end else if(N4650) begin
      content_q[73] <= content_n_1__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[72] <= 1'b0;
    end else if(N4650) begin
      content_q[72] <= content_n_1__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[71] <= 1'b0;
    end else if(N4650) begin
      content_q[71] <= content_n_1__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[70] <= 1'b0;
    end else if(N4650) begin
      content_q[70] <= content_n_1__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[69] <= 1'b0;
    end else if(N4650) begin
      content_q[69] <= content_n_1__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[68] <= 1'b0;
    end else if(N4650) begin
      content_q[68] <= content_n_1__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[67] <= 1'b0;
    end else if(N4650) begin
      content_q[67] <= content_n_1__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[66] <= 1'b0;
    end else if(N4650) begin
      content_q[66] <= content_n_1__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[65] <= 1'b0;
    end else if(N4650) begin
      content_q[65] <= content_n_1__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[64] <= 1'b0;
    end else if(N4650) begin
      content_q[64] <= content_n_1__v_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[63] <= 1'b0;
    end else if(N4650) begin
      content_q[63] <= content_n_0__reserved__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[62] <= 1'b0;
    end else if(N4650) begin
      content_q[62] <= content_n_0__reserved__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[61] <= 1'b0;
    end else if(N4650) begin
      content_q[61] <= content_n_0__reserved__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[60] <= 1'b0;
    end else if(N4650) begin
      content_q[60] <= content_n_0__reserved__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[59] <= 1'b0;
    end else if(N4650) begin
      content_q[59] <= content_n_0__reserved__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[58] <= 1'b0;
    end else if(N4650) begin
      content_q[58] <= content_n_0__reserved__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[57] <= 1'b0;
    end else if(N4650) begin
      content_q[57] <= content_n_0__reserved__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[56] <= 1'b0;
    end else if(N4650) begin
      content_q[56] <= content_n_0__reserved__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[55] <= 1'b0;
    end else if(N4650) begin
      content_q[55] <= content_n_0__reserved__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[54] <= 1'b0;
    end else if(N4650) begin
      content_q[54] <= content_n_0__reserved__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[53] <= 1'b0;
    end else if(N4650) begin
      content_q[53] <= content_n_0__ppn__43_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[52] <= 1'b0;
    end else if(N4650) begin
      content_q[52] <= content_n_0__ppn__42_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[51] <= 1'b0;
    end else if(N4650) begin
      content_q[51] <= content_n_0__ppn__41_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[50] <= 1'b0;
    end else if(N4650) begin
      content_q[50] <= content_n_0__ppn__40_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[49] <= 1'b0;
    end else if(N4650) begin
      content_q[49] <= content_n_0__ppn__39_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[48] <= 1'b0;
    end else if(N4650) begin
      content_q[48] <= content_n_0__ppn__38_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[47] <= 1'b0;
    end else if(N4650) begin
      content_q[47] <= content_n_0__ppn__37_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[46] <= 1'b0;
    end else if(N4650) begin
      content_q[46] <= content_n_0__ppn__36_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[45] <= 1'b0;
    end else if(N4650) begin
      content_q[45] <= content_n_0__ppn__35_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[44] <= 1'b0;
    end else if(N4650) begin
      content_q[44] <= content_n_0__ppn__34_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[43] <= 1'b0;
    end else if(N4650) begin
      content_q[43] <= content_n_0__ppn__33_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[42] <= 1'b0;
    end else if(N4650) begin
      content_q[42] <= content_n_0__ppn__32_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[41] <= 1'b0;
    end else if(N4650) begin
      content_q[41] <= content_n_0__ppn__31_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[40] <= 1'b0;
    end else if(N4650) begin
      content_q[40] <= content_n_0__ppn__30_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[39] <= 1'b0;
    end else if(N4650) begin
      content_q[39] <= content_n_0__ppn__29_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[38] <= 1'b0;
    end else if(N4650) begin
      content_q[38] <= content_n_0__ppn__28_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[37] <= 1'b0;
    end else if(N4650) begin
      content_q[37] <= content_n_0__ppn__27_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[36] <= 1'b0;
    end else if(N4650) begin
      content_q[36] <= content_n_0__ppn__26_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[35] <= 1'b0;
    end else if(N4650) begin
      content_q[35] <= content_n_0__ppn__25_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[34] <= 1'b0;
    end else if(N4650) begin
      content_q[34] <= content_n_0__ppn__24_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[33] <= 1'b0;
    end else if(N4650) begin
      content_q[33] <= content_n_0__ppn__23_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[32] <= 1'b0;
    end else if(N4650) begin
      content_q[32] <= content_n_0__ppn__22_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[31] <= 1'b0;
    end else if(N4650) begin
      content_q[31] <= content_n_0__ppn__21_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[30] <= 1'b0;
    end else if(N4650) begin
      content_q[30] <= content_n_0__ppn__20_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[29] <= 1'b0;
    end else if(N4650) begin
      content_q[29] <= content_n_0__ppn__19_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[28] <= 1'b0;
    end else if(N4650) begin
      content_q[28] <= content_n_0__ppn__18_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[27] <= 1'b0;
    end else if(N4650) begin
      content_q[27] <= content_n_0__ppn__17_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[26] <= 1'b0;
    end else if(N4650) begin
      content_q[26] <= content_n_0__ppn__16_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[25] <= 1'b0;
    end else if(N4650) begin
      content_q[25] <= content_n_0__ppn__15_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[24] <= 1'b0;
    end else if(N4650) begin
      content_q[24] <= content_n_0__ppn__14_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[23] <= 1'b0;
    end else if(N4650) begin
      content_q[23] <= content_n_0__ppn__13_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[22] <= 1'b0;
    end else if(N4650) begin
      content_q[22] <= content_n_0__ppn__12_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[21] <= 1'b0;
    end else if(N4650) begin
      content_q[21] <= content_n_0__ppn__11_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[20] <= 1'b0;
    end else if(N4650) begin
      content_q[20] <= content_n_0__ppn__10_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[19] <= 1'b0;
    end else if(N4650) begin
      content_q[19] <= content_n_0__ppn__9_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[18] <= 1'b0;
    end else if(N4650) begin
      content_q[18] <= content_n_0__ppn__8_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[17] <= 1'b0;
    end else if(N4650) begin
      content_q[17] <= content_n_0__ppn__7_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[16] <= 1'b0;
    end else if(N4650) begin
      content_q[16] <= content_n_0__ppn__6_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[15] <= 1'b0;
    end else if(N4650) begin
      content_q[15] <= content_n_0__ppn__5_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[14] <= 1'b0;
    end else if(N4650) begin
      content_q[14] <= content_n_0__ppn__4_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[13] <= 1'b0;
    end else if(N4650) begin
      content_q[13] <= content_n_0__ppn__3_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[12] <= 1'b0;
    end else if(N4650) begin
      content_q[12] <= content_n_0__ppn__2_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[11] <= 1'b0;
    end else if(N4650) begin
      content_q[11] <= content_n_0__ppn__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[10] <= 1'b0;
    end else if(N4650) begin
      content_q[10] <= content_n_0__ppn__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[9] <= 1'b0;
    end else if(N4650) begin
      content_q[9] <= content_n_0__rsw__1_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[8] <= 1'b0;
    end else if(N4650) begin
      content_q[8] <= content_n_0__rsw__0_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[7] <= 1'b0;
    end else if(N4650) begin
      content_q[7] <= content_n_0__d_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[6] <= 1'b0;
    end else if(N4650) begin
      content_q[6] <= content_n_0__a_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[5] <= 1'b0;
    end else if(N4650) begin
      content_q[5] <= content_n_0__g_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[4] <= 1'b0;
    end else if(N4650) begin
      content_q[4] <= content_n_0__u_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[3] <= 1'b0;
    end else if(N4650) begin
      content_q[3] <= content_n_0__x_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[2] <= 1'b0;
    end else if(N4650) begin
      content_q[2] <= content_n_0__w_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[1] <= 1'b0;
    end else if(N4650) begin
      content_q[1] <= content_n_0__r_;
    end 
  end


  always @(posedge clk_i or posedge N4781) begin
    if(N4781) begin
      content_q[0] <= 1'b0;
    end else if(N4650) begin
      content_q[0] <= content_n_0__v_;
    end 
  end

  assign N4838 = ~lu_asid_i[0];
  assign N157 = (N32)? tags_q[2] : 
                (N156)? 1'b0 : 1'b0;
  assign N32 = N155;
  assign { N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158 } = (N32)? content_q[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N156)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N222 = (N33)? N157 : 
                (N34)? 1'b0 : 1'b0;
  assign N33 = N152;
  assign N34 = N153;
  assign { N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223 } = (N33)? { N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N287 = (N33)? N155 : 
                (N34)? 1'b0 : 1'b0;
  assign { N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288 } = (N35)? content_q[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N36)? { N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223 } : 1'b0;
  assign N35 = tags_q[1];
  assign N36 = N150;
  assign N352 = (N35)? 1'b1 : 
                (N36)? N287 : 1'b0;
  assign N353 = (N35)? 1'b0 : 
                (N36)? N222 : 1'b0;
  assign N354 = (N37)? N353 : 
                (N148)? 1'b0 : 1'b0;
  assign N37 = N147;
  assign N355 = (N37)? tags_q[1] : 
                (N148)? 1'b0 : 1'b0;
  assign { N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356 } = (N37)? { N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N148)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N420 = (N37)? N352 : 
                (N148)? 1'b0 : 1'b0;
  assign lu_hit[0] = (N37)? N352 : 
                     (N148)? 1'b0 : 1'b0;
  assign N433 = (N38)? tags_q[33] : 
                (N432)? N354 : 1'b0;
  assign N38 = N431;
  assign { N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434 } = (N38)? content_q[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N432)? { N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356 } : 1'b0;
  assign N498 = (N38)? 1'b1 : 
                (N432)? N420 : 1'b0;
  assign N499 = (N39)? N431 : 
                (N40)? 1'b0 : 1'b0;
  assign N39 = N428;
  assign N40 = N429;
  assign N500 = (N39)? N433 : 
                (N40)? N354 : 1'b0;
  assign { N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501 } = (N39)? { N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N40)? { N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356 } : 1'b0;
  assign N565 = (N39)? N498 : 
                (N40)? N420 : 1'b0;
  assign N566 = (N41)? 1'b1 : 
                (N42)? N355 : 1'b0;
  assign N41 = tags_q[32];
  assign N42 = N426;
  assign { N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567 } = (N41)? content_q[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N42)? { N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501 } : 1'b0;
  assign N631 = (N41)? 1'b1 : 
                (N42)? N565 : 1'b0;
  assign N632 = (N41)? 1'b1 : 
                (N42)? N499 : 1'b0;
  assign N633 = (N41)? N354 : 
                (N42)? N500 : 1'b0;
  assign N634 = (N43)? N633 : 
                (N424)? N354 : 1'b0;
  assign N43 = N423;
  assign N635 = (N43)? N566 : 
                (N424)? N355 : 1'b0;
  assign { N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636 } = (N43)? { N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N424)? { N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356 } : 1'b0;
  assign N700 = (N43)? N631 : 
                (N424)? N420 : 1'b0;
  assign lu_hit[1] = (N43)? N632 : 
                     (N424)? 1'b0 : 1'b0;
  assign N713 = (N44)? tags_q[64] : 
                (N712)? N634 : 1'b0;
  assign N44 = N711;
  assign { N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714 } = (N44)? content_q[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N712)? { N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636 } : 1'b0;
  assign N778 = (N44)? 1'b1 : 
                (N712)? N700 : 1'b0;
  assign N779 = (N45)? N711 : 
                (N46)? 1'b0 : 1'b0;
  assign N45 = N708;
  assign N46 = N709;
  assign N780 = (N45)? N713 : 
                (N46)? N634 : 1'b0;
  assign { N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781 } = (N45)? { N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N46)? { N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636 } : 1'b0;
  assign N845 = (N45)? N778 : 
                (N46)? N700 : 1'b0;
  assign N846 = (N47)? 1'b1 : 
                (N48)? N635 : 1'b0;
  assign N47 = tags_q[63];
  assign N48 = N706;
  assign { N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847 } = (N47)? content_q[191:128] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N48)? { N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781 } : 1'b0;
  assign N911 = (N47)? 1'b1 : 
                (N48)? N845 : 1'b0;
  assign N912 = (N47)? 1'b1 : 
                (N48)? N779 : 1'b0;
  assign N913 = (N47)? N634 : 
                (N48)? N780 : 1'b0;
  assign N914 = (N49)? N913 : 
                (N704)? N634 : 1'b0;
  assign N49 = N703;
  assign N915 = (N49)? N846 : 
                (N704)? N635 : 1'b0;
  assign { N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916 } = (N49)? { N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N704)? { N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636 } : 1'b0;
  assign N980 = (N49)? N911 : 
                (N704)? N700 : 1'b0;
  assign lu_hit[2] = (N49)? N912 : 
                     (N704)? 1'b0 : 1'b0;
  assign N993 = (N50)? tags_q[95] : 
                (N992)? N914 : 1'b0;
  assign N50 = N991;
  assign { N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994 } = (N50)? content_q[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N992)? { N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916 } : 1'b0;
  assign N1058 = (N50)? 1'b1 : 
                 (N992)? N980 : 1'b0;
  assign N1059 = (N51)? N991 : 
                 (N52)? 1'b0 : 1'b0;
  assign N51 = N988;
  assign N52 = N989;
  assign N1060 = (N51)? N993 : 
                 (N52)? N914 : 1'b0;
  assign { N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061 } = (N51)? { N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N52)? { N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916 } : 1'b0;
  assign N1125 = (N51)? N1058 : 
                 (N52)? N980 : 1'b0;
  assign N1126 = (N53)? 1'b1 : 
                 (N54)? N915 : 1'b0;
  assign N53 = tags_q[94];
  assign N54 = N986;
  assign { N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127 } = (N53)? content_q[255:192] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N54)? { N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061 } : 1'b0;
  assign N1191 = (N53)? 1'b1 : 
                 (N54)? N1125 : 1'b0;
  assign N1192 = (N53)? 1'b1 : 
                 (N54)? N1059 : 1'b0;
  assign N1193 = (N53)? N914 : 
                 (N54)? N1060 : 1'b0;
  assign N1194 = (N55)? N1193 : 
                 (N984)? N914 : 1'b0;
  assign N55 = N983;
  assign N1195 = (N55)? N1126 : 
                 (N984)? N915 : 1'b0;
  assign { N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196 } = (N55)? { N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N984)? { N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916 } : 1'b0;
  assign N1260 = (N55)? N1191 : 
                 (N984)? N980 : 1'b0;
  assign lu_hit[3] = (N55)? N1192 : 
                     (N984)? 1'b0 : 1'b0;
  assign N1273 = (N56)? tags_q[126] : 
                 (N1272)? N1194 : 1'b0;
  assign N56 = N1271;
  assign { N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274 } = (N56)? content_q[319:256] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1272)? { N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196 } : 1'b0;
  assign N1338 = (N56)? 1'b1 : 
                 (N1272)? N1260 : 1'b0;
  assign N1339 = (N57)? N1271 : 
                 (N58)? 1'b0 : 1'b0;
  assign N57 = N1268;
  assign N58 = N1269;
  assign N1340 = (N57)? N1273 : 
                 (N58)? N1194 : 1'b0;
  assign { N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341 } = (N57)? { N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N58)? { N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196 } : 1'b0;
  assign N1405 = (N57)? N1338 : 
                 (N58)? N1260 : 1'b0;
  assign N1406 = (N59)? 1'b1 : 
                 (N60)? N1195 : 1'b0;
  assign N59 = tags_q[125];
  assign N60 = N1266;
  assign { N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407 } = (N59)? content_q[319:256] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N60)? { N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341 } : 1'b0;
  assign N1471 = (N59)? 1'b1 : 
                 (N60)? N1405 : 1'b0;
  assign N1472 = (N59)? 1'b1 : 
                 (N60)? N1339 : 1'b0;
  assign N1473 = (N59)? N1194 : 
                 (N60)? N1340 : 1'b0;
  assign N1474 = (N61)? N1473 : 
                 (N1264)? N1194 : 1'b0;
  assign N61 = N1263;
  assign N1475 = (N61)? N1406 : 
                 (N1264)? N1195 : 1'b0;
  assign { N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476 } = (N61)? { N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1264)? { N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196 } : 1'b0;
  assign N1540 = (N61)? N1471 : 
                 (N1264)? N1260 : 1'b0;
  assign lu_hit[4] = (N61)? N1472 : 
                     (N1264)? 1'b0 : 1'b0;
  assign N1553 = (N62)? tags_q[157] : 
                 (N1552)? N1474 : 1'b0;
  assign N62 = N1551;
  assign { N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554 } = (N62)? content_q[383:320] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1552)? { N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476 } : 1'b0;
  assign N1618 = (N62)? 1'b1 : 
                 (N1552)? N1540 : 1'b0;
  assign N1619 = (N63)? N1551 : 
                 (N64)? 1'b0 : 1'b0;
  assign N63 = N1548;
  assign N64 = N1549;
  assign N1620 = (N63)? N1553 : 
                 (N64)? N1474 : 1'b0;
  assign { N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621 } = (N63)? { N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N64)? { N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476 } : 1'b0;
  assign N1685 = (N63)? N1618 : 
                 (N64)? N1540 : 1'b0;
  assign N1686 = (N65)? 1'b1 : 
                 (N66)? N1475 : 1'b0;
  assign N65 = tags_q[156];
  assign N66 = N1546;
  assign { N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687 } = (N65)? content_q[383:320] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N66)? { N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621 } : 1'b0;
  assign N1751 = (N65)? 1'b1 : 
                 (N66)? N1685 : 1'b0;
  assign N1752 = (N65)? 1'b1 : 
                 (N66)? N1619 : 1'b0;
  assign N1753 = (N65)? N1474 : 
                 (N66)? N1620 : 1'b0;
  assign N1754 = (N67)? N1753 : 
                 (N1544)? N1474 : 1'b0;
  assign N67 = N1543;
  assign N1755 = (N67)? N1686 : 
                 (N1544)? N1475 : 1'b0;
  assign { N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756 } = (N67)? { N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1544)? { N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476 } : 1'b0;
  assign N1820 = (N67)? N1751 : 
                 (N1544)? N1540 : 1'b0;
  assign lu_hit[5] = (N67)? N1752 : 
                     (N1544)? 1'b0 : 1'b0;
  assign N1833 = (N68)? tags_q[188] : 
                 (N1832)? N1754 : 1'b0;
  assign N68 = N1831;
  assign { N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834 } = (N68)? content_q[447:384] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1832)? { N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756 } : 1'b0;
  assign N1898 = (N68)? 1'b1 : 
                 (N1832)? N1820 : 1'b0;
  assign N1899 = (N69)? N1831 : 
                 (N70)? 1'b0 : 1'b0;
  assign N69 = N1828;
  assign N70 = N1829;
  assign N1900 = (N69)? N1833 : 
                 (N70)? N1754 : 1'b0;
  assign { N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901 } = (N69)? { N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N70)? { N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756 } : 1'b0;
  assign N1965 = (N69)? N1898 : 
                 (N70)? N1820 : 1'b0;
  assign N1966 = (N71)? 1'b1 : 
                 (N72)? N1755 : 1'b0;
  assign N71 = tags_q[187];
  assign N72 = N1826;
  assign { N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967 } = (N71)? content_q[447:384] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N72)? { N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901 } : 1'b0;
  assign N2031 = (N71)? 1'b1 : 
                 (N72)? N1965 : 1'b0;
  assign N2032 = (N71)? 1'b1 : 
                 (N72)? N1899 : 1'b0;
  assign N2033 = (N71)? N1754 : 
                 (N72)? N1900 : 1'b0;
  assign N2034 = (N73)? N2033 : 
                 (N1824)? N1754 : 1'b0;
  assign N73 = N1823;
  assign N2035 = (N73)? N1966 : 
                 (N1824)? N1755 : 1'b0;
  assign { N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036 } = (N73)? { N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1824)? { N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756 } : 1'b0;
  assign N2100 = (N73)? N2031 : 
                 (N1824)? N1820 : 1'b0;
  assign lu_hit[6] = (N73)? N2032 : 
                     (N1824)? 1'b0 : 1'b0;
  assign N2113 = (N74)? tags_q[219] : 
                 (N2112)? N2034 : 1'b0;
  assign N74 = N2111;
  assign { N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114 } = (N74)? content_q[511:448] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2112)? { N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036 } : 1'b0;
  assign N2178 = (N74)? 1'b1 : 
                 (N2112)? N2100 : 1'b0;
  assign N2179 = (N75)? N2111 : 
                 (N76)? 1'b0 : 1'b0;
  assign N75 = N2108;
  assign N76 = N2109;
  assign N2180 = (N75)? N2113 : 
                 (N76)? N2034 : 1'b0;
  assign { N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181 } = (N75)? { N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N76)? { N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036 } : 1'b0;
  assign N2245 = (N75)? N2178 : 
                 (N76)? N2100 : 1'b0;
  assign N2246 = (N77)? 1'b1 : 
                 (N78)? N2035 : 1'b0;
  assign N77 = tags_q[218];
  assign N78 = N2106;
  assign { N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247 } = (N77)? content_q[511:448] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N78)? { N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181 } : 1'b0;
  assign N2311 = (N77)? 1'b1 : 
                 (N78)? N2245 : 1'b0;
  assign N2312 = (N77)? 1'b1 : 
                 (N78)? N2179 : 1'b0;
  assign N2313 = (N77)? N2034 : 
                 (N78)? N2180 : 1'b0;
  assign N2314 = (N79)? N2313 : 
                 (N2104)? N2034 : 1'b0;
  assign N79 = N2103;
  assign N2315 = (N79)? N2246 : 
                 (N2104)? N2035 : 1'b0;
  assign { N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316 } = (N79)? { N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2104)? { N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036 } : 1'b0;
  assign N2380 = (N79)? N2311 : 
                 (N2104)? N2100 : 1'b0;
  assign lu_hit[7] = (N79)? N2312 : 
                     (N2104)? 1'b0 : 1'b0;
  assign N2393 = (N80)? tags_q[250] : 
                 (N2392)? N2314 : 1'b0;
  assign N80 = N2391;
  assign { N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394 } = (N80)? content_q[575:512] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2392)? { N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316 } : 1'b0;
  assign N2458 = (N80)? 1'b1 : 
                 (N2392)? N2380 : 1'b0;
  assign N2459 = (N81)? N2391 : 
                 (N82)? 1'b0 : 1'b0;
  assign N81 = N2388;
  assign N82 = N2389;
  assign N2460 = (N81)? N2393 : 
                 (N82)? N2314 : 1'b0;
  assign { N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461 } = (N81)? { N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N82)? { N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316 } : 1'b0;
  assign N2525 = (N81)? N2458 : 
                 (N82)? N2380 : 1'b0;
  assign N2526 = (N83)? 1'b1 : 
                 (N84)? N2315 : 1'b0;
  assign N83 = tags_q[249];
  assign N84 = N2386;
  assign { N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527 } = (N83)? content_q[575:512] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N84)? { N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461 } : 1'b0;
  assign N2591 = (N83)? 1'b1 : 
                 (N84)? N2525 : 1'b0;
  assign N2592 = (N83)? 1'b1 : 
                 (N84)? N2459 : 1'b0;
  assign N2593 = (N83)? N2314 : 
                 (N84)? N2460 : 1'b0;
  assign N2594 = (N85)? N2593 : 
                 (N2384)? N2314 : 1'b0;
  assign N85 = N2383;
  assign N2595 = (N85)? N2526 : 
                 (N2384)? N2315 : 1'b0;
  assign { N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596 } = (N85)? { N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2384)? { N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316 } : 1'b0;
  assign N2660 = (N85)? N2591 : 
                 (N2384)? N2380 : 1'b0;
  assign lu_hit[8] = (N85)? N2592 : 
                     (N2384)? 1'b0 : 1'b0;
  assign N2673 = (N86)? tags_q[281] : 
                 (N2672)? N2594 : 1'b0;
  assign N86 = N2671;
  assign { N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674 } = (N86)? content_q[639:576] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2672)? { N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596 } : 1'b0;
  assign N2738 = (N86)? 1'b1 : 
                 (N2672)? N2660 : 1'b0;
  assign N2739 = (N87)? N2671 : 
                 (N88)? 1'b0 : 1'b0;
  assign N87 = N2668;
  assign N88 = N2669;
  assign N2740 = (N87)? N2673 : 
                 (N88)? N2594 : 1'b0;
  assign { N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741 } = (N87)? { N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N88)? { N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596 } : 1'b0;
  assign N2805 = (N87)? N2738 : 
                 (N88)? N2660 : 1'b0;
  assign N2806 = (N89)? 1'b1 : 
                 (N90)? N2595 : 1'b0;
  assign N89 = tags_q[280];
  assign N90 = N2666;
  assign { N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807 } = (N89)? content_q[639:576] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N90)? { N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741 } : 1'b0;
  assign N2871 = (N89)? 1'b1 : 
                 (N90)? N2805 : 1'b0;
  assign N2872 = (N89)? 1'b1 : 
                 (N90)? N2739 : 1'b0;
  assign N2873 = (N89)? N2594 : 
                 (N90)? N2740 : 1'b0;
  assign N2874 = (N91)? N2873 : 
                 (N2664)? N2594 : 1'b0;
  assign N91 = N2663;
  assign N2875 = (N91)? N2806 : 
                 (N2664)? N2595 : 1'b0;
  assign { N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876 } = (N91)? { N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2664)? { N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596 } : 1'b0;
  assign N2940 = (N91)? N2871 : 
                 (N2664)? N2660 : 1'b0;
  assign lu_hit[9] = (N91)? N2872 : 
                     (N2664)? 1'b0 : 1'b0;
  assign N2953 = (N92)? tags_q[312] : 
                 (N2952)? N2874 : 1'b0;
  assign N92 = N2951;
  assign { N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954 } = (N92)? content_q[703:640] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2952)? { N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876 } : 1'b0;
  assign N3018 = (N92)? 1'b1 : 
                 (N2952)? N2940 : 1'b0;
  assign N3019 = (N93)? N2951 : 
                 (N94)? 1'b0 : 1'b0;
  assign N93 = N2948;
  assign N94 = N2949;
  assign N3020 = (N93)? N2953 : 
                 (N94)? N2874 : 1'b0;
  assign { N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021 } = (N93)? { N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N94)? { N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876 } : 1'b0;
  assign N3085 = (N93)? N3018 : 
                 (N94)? N2940 : 1'b0;
  assign N3086 = (N95)? 1'b1 : 
                 (N96)? N2875 : 1'b0;
  assign N95 = tags_q[311];
  assign N96 = N2946;
  assign { N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087 } = (N95)? content_q[703:640] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N96)? { N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021 } : 1'b0;
  assign N3151 = (N95)? 1'b1 : 
                 (N96)? N3085 : 1'b0;
  assign N3152 = (N95)? 1'b1 : 
                 (N96)? N3019 : 1'b0;
  assign N3153 = (N95)? N2874 : 
                 (N96)? N3020 : 1'b0;
  assign N3154 = (N97)? N3153 : 
                 (N2944)? N2874 : 1'b0;
  assign N97 = N2943;
  assign N3155 = (N97)? N3086 : 
                 (N2944)? N2875 : 1'b0;
  assign { N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156 } = (N97)? { N3150, N3149, N3148, N3147, N3146, N3145, N3144, N3143, N3142, N3141, N3140, N3139, N3138, N3137, N3136, N3135, N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2944)? { N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876 } : 1'b0;
  assign N3220 = (N97)? N3151 : 
                 (N2944)? N2940 : 1'b0;
  assign lu_hit[10] = (N97)? N3152 : 
                      (N2944)? 1'b0 : 1'b0;
  assign N3233 = (N98)? tags_q[343] : 
                 (N3232)? N3154 : 1'b0;
  assign N98 = N3231;
  assign { N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234 } = (N98)? content_q[767:704] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3232)? { N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156 } : 1'b0;
  assign N3298 = (N98)? 1'b1 : 
                 (N3232)? N3220 : 1'b0;
  assign N3299 = (N99)? N3231 : 
                 (N100)? 1'b0 : 1'b0;
  assign N99 = N3228;
  assign N100 = N3229;
  assign N3300 = (N99)? N3233 : 
                 (N100)? N3154 : 1'b0;
  assign { N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301 } = (N99)? { N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276, N3275, N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N100)? { N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156 } : 1'b0;
  assign N3365 = (N99)? N3298 : 
                 (N100)? N3220 : 1'b0;
  assign N3366 = (N101)? 1'b1 : 
                 (N102)? N3155 : 1'b0;
  assign N101 = tags_q[342];
  assign N102 = N3226;
  assign { N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367 } = (N101)? content_q[767:704] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N102)? { N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301 } : 1'b0;
  assign N3431 = (N101)? 1'b1 : 
                 (N102)? N3365 : 1'b0;
  assign N3432 = (N101)? 1'b1 : 
                 (N102)? N3299 : 1'b0;
  assign N3433 = (N101)? N3154 : 
                 (N102)? N3300 : 1'b0;
  assign N3434 = (N103)? N3433 : 
                 (N3224)? N3154 : 1'b0;
  assign N103 = N3223;
  assign N3435 = (N103)? N3366 : 
                 (N3224)? N3155 : 1'b0;
  assign { N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436 } = (N103)? { N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406, N3405, N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3224)? { N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156 } : 1'b0;
  assign N3500 = (N103)? N3431 : 
                 (N3224)? N3220 : 1'b0;
  assign lu_hit[11] = (N103)? N3432 : 
                      (N3224)? 1'b0 : 1'b0;
  assign N3513 = (N104)? tags_q[374] : 
                 (N3512)? N3434 : 1'b0;
  assign N104 = N3511;
  assign { N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514 } = (N104)? content_q[831:768] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3512)? { N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436 } : 1'b0;
  assign N3578 = (N104)? 1'b1 : 
                 (N3512)? N3500 : 1'b0;
  assign N3579 = (N105)? N3511 : 
                 (N106)? 1'b0 : 1'b0;
  assign N105 = N3508;
  assign N106 = N3509;
  assign N3580 = (N105)? N3513 : 
                 (N106)? N3434 : 1'b0;
  assign { N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581 } = (N105)? { N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N106)? { N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436 } : 1'b0;
  assign N3645 = (N105)? N3578 : 
                 (N106)? N3500 : 1'b0;
  assign N3646 = (N107)? 1'b1 : 
                 (N108)? N3435 : 1'b0;
  assign N107 = tags_q[373];
  assign N108 = N3506;
  assign { N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647 } = (N107)? content_q[831:768] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N108)? { N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581 } : 1'b0;
  assign N3711 = (N107)? 1'b1 : 
                 (N108)? N3645 : 1'b0;
  assign N3712 = (N107)? 1'b1 : 
                 (N108)? N3579 : 1'b0;
  assign N3713 = (N107)? N3434 : 
                 (N108)? N3580 : 1'b0;
  assign N3714 = (N109)? N3713 : 
                 (N3504)? N3434 : 1'b0;
  assign N109 = N3503;
  assign N3715 = (N109)? N3646 : 
                 (N3504)? N3435 : 1'b0;
  assign { N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716 } = (N109)? { N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666, N3665, N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3504)? { N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436 } : 1'b0;
  assign N3780 = (N109)? N3711 : 
                 (N3504)? N3500 : 1'b0;
  assign lu_hit[12] = (N109)? N3712 : 
                      (N3504)? 1'b0 : 1'b0;
  assign N3793 = (N110)? tags_q[405] : 
                 (N3792)? N3714 : 1'b0;
  assign N110 = N3791;
  assign { N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794 } = (N110)? content_q[895:832] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3792)? { N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716 } : 1'b0;
  assign N3858 = (N110)? 1'b1 : 
                 (N3792)? N3780 : 1'b0;
  assign N3859 = (N111)? N3791 : 
                 (N112)? 1'b0 : 1'b0;
  assign N111 = N3788;
  assign N112 = N3789;
  assign N3860 = (N111)? N3793 : 
                 (N112)? N3714 : 1'b0;
  assign { N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861 } = (N111)? { N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796, N3795, N3794 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N112)? { N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716 } : 1'b0;
  assign N3925 = (N111)? N3858 : 
                 (N112)? N3780 : 1'b0;
  assign N3926 = (N113)? 1'b1 : 
                 (N114)? N3715 : 1'b0;
  assign N113 = tags_q[404];
  assign N114 = N3786;
  assign { N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927 } = (N113)? content_q[895:832] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N114)? { N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861 } : 1'b0;
  assign N3991 = (N113)? 1'b1 : 
                 (N114)? N3925 : 1'b0;
  assign N3992 = (N113)? 1'b1 : 
                 (N114)? N3859 : 1'b0;
  assign N3993 = (N113)? N3714 : 
                 (N114)? N3860 : 1'b0;
  assign N3994 = (N115)? N3993 : 
                 (N3784)? N3714 : 1'b0;
  assign N115 = N3783;
  assign N3995 = (N115)? N3926 : 
                 (N3784)? N3715 : 1'b0;
  assign { N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996 } = (N115)? { N3990, N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3784)? { N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731, N3730, N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716 } : 1'b0;
  assign N4060 = (N115)? N3991 : 
                 (N3784)? N3780 : 1'b0;
  assign lu_hit[13] = (N115)? N3992 : 
                      (N3784)? 1'b0 : 1'b0;
  assign N4073 = (N116)? tags_q[436] : 
                 (N4072)? N3994 : 1'b0;
  assign N116 = N4071;
  assign { N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074 } = (N116)? content_q[959:896] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4072)? { N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996 } : 1'b0;
  assign N4138 = (N116)? 1'b1 : 
                 (N4072)? N4060 : 1'b0;
  assign N4139 = (N117)? N4071 : 
                 (N118)? 1'b0 : 1'b0;
  assign N117 = N4068;
  assign N118 = N4069;
  assign N4140 = (N117)? N4073 : 
                 (N118)? N3994 : 1'b0;
  assign { N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141 } = (N117)? { N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, N4128, N4127, N4126, N4125, N4124, N4123, N4122, N4121, N4120, N4119, N4118, N4117, N4116, N4115, N4114, N4113, N4112, N4111, N4110, N4109, N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095, N4094, N4093, N4092, N4091, N4090, N4089, N4088, N4087, N4086, N4085, N4084, N4083, N4082, N4081, N4080, N4079, N4078, N4077, N4076, N4075, N4074 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N118)? { N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996 } : 1'b0;
  assign N4205 = (N117)? N4138 : 
                 (N118)? N4060 : 1'b0;
  assign N4206 = (N119)? 1'b1 : 
                 (N120)? N3995 : 1'b0;
  assign N119 = tags_q[435];
  assign N120 = N4066;
  assign { N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207 } = (N119)? content_q[959:896] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N120)? { N4204, N4203, N4202, N4201, N4200, N4199, N4198, N4197, N4196, N4195, N4194, N4193, N4192, N4191, N4190, N4189, N4188, N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174, N4173, N4172, N4171, N4170, N4169, N4168, N4167, N4166, N4165, N4164, N4163, N4162, N4161, N4160, N4159, N4158, N4157, N4156, N4155, N4154, N4153, N4152, N4151, N4150, N4149, N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141 } : 1'b0;
  assign N4271 = (N119)? 1'b1 : 
                 (N120)? N4205 : 1'b0;
  assign N4272 = (N119)? 1'b1 : 
                 (N120)? N4139 : 1'b0;
  assign N4273 = (N119)? N3994 : 
                 (N120)? N4140 : 1'b0;
  assign N4274 = (N121)? N4273 : 
                 (N4064)? N3994 : 1'b0;
  assign N121 = N4063;
  assign N4275 = (N121)? N4206 : 
                 (N4064)? N3995 : 1'b0;
  assign { N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276 } = (N121)? { N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263, N4262, N4261, N4260, N4259, N4258, N4257, N4256, N4255, N4254, N4253, N4252, N4251, N4250, N4249, N4248, N4247, N4246, N4245, N4244, N4243, N4242, N4241, N4240, N4239, N4238, N4237, N4236, N4235, N4234, N4233, N4232, N4231, N4230, N4229, N4228, N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, N4207 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4064)? { N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996 } : 1'b0;
  assign N4340 = (N121)? N4271 : 
                 (N4064)? N4060 : 1'b0;
  assign lu_hit[14] = (N121)? N4272 : 
                      (N4064)? 1'b0 : 1'b0;
  assign N4353 = (N122)? tags_q[467] : 
                 (N4352)? N4274 : 1'b0;
  assign N122 = N4351;
  assign { N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354 } = (N122)? content_q[1023:960] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N4352)? { N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276 } : 1'b0;
  assign N4418 = (N122)? 1'b1 : 
                 (N4352)? N4340 : 1'b0;
  assign N4419 = (N123)? N4351 : 
                 (N124)? 1'b0 : 1'b0;
  assign N123 = N4348;
  assign N124 = N4349;
  assign N4420 = (N123)? N4353 : 
                 (N124)? N4274 : 1'b0;
  assign { N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421 } = (N123)? { N4417, N4416, N4415, N4414, N4413, N4412, N4411, N4410, N4409, N4408, N4407, N4406, N4405, N4404, N4403, N4402, N4401, N4400, N4399, N4398, N4397, N4396, N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, N4375, N4374, N4373, N4372, N4371, N4370, N4369, N4368, N4367, N4366, N4365, N4364, N4363, N4362, N4361, N4360, N4359, N4358, N4357, N4356, N4355, N4354 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N124)? { N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276 } : 1'b0;
  assign N4485 = (N123)? N4418 : 
                 (N124)? N4340 : 1'b0;
  assign N4486 = (N125)? 1'b1 : 
                 (N126)? N4275 : 1'b0;
  assign N125 = tags_q[466];
  assign N126 = N4346;
  assign { N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487 } = (N125)? content_q[1023:960] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N126)? { N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, N4465, N4464, N4463, N4462, N4461, N4460, N4459, N4458, N4457, N4456, N4455, N4454, N4453, N4452, N4451, N4450, N4449, N4448, N4447, N4446, N4445, N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431, N4430, N4429, N4428, N4427, N4426, N4425, N4424, N4423, N4422, N4421 } : 1'b0;
  assign N4551 = (N125)? 1'b1 : 
                 (N126)? N4485 : 1'b0;
  assign N4552 = (N125)? 1'b1 : 
                 (N126)? N4419 : 1'b0;
  assign N4553 = (N125)? N4274 : 
                 (N126)? N4420 : 1'b0;
  assign lu_is_2M_o = (N127)? N4553 : 
                      (N4344)? N4274 : 1'b0;
  assign N127 = N4343;
  assign lu_is_1G_o = (N127)? N4486 : 
                      (N4344)? N4275 : 1'b0;
  assign lu_content_o = (N127)? { N4550, N4549, N4548, N4547, N4546, N4545, N4544, N4543, N4542, N4541, N4540, N4539, N4538, N4537, N4536, N4535, N4534, N4533, N4532, N4531, N4530, N4529, N4528, N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513, N4512, N4511, N4510, N4509, N4508, N4507, N4506, N4505, N4504, N4503, N4502, N4501, N4500, N4499, N4498, N4497, N4496, N4495, N4494, N4493, N4492, N4491, N4490, N4489, N4488, N4487 } : 
                        (N4344)? { N4339, N4338, N4337, N4336, N4335, N4334, N4333, N4332, N4331, N4330, N4329, N4328, N4327, N4326, N4325, N4324, N4323, N4322, N4321, N4320, N4319, N4318, N4317, N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, N4296, N4295, N4294, N4293, N4292, N4291, N4290, N4289, N4288, N4287, N4286, N4285, N4284, N4283, N4282, N4281, N4280, N4279, N4278, N4277, N4276 } : 1'b0;
  assign lu_hit_o = (N127)? N4551 : 
                    (N4344)? N4340 : 1'b0;
  assign lu_hit[15] = (N127)? N4552 : 
                      (N4344)? 1'b0 : 1'b0;
  assign tags_n_0__valid_ = (N128)? 1'b0 : 
                            (N4651)? 1'b1 : 
                            (N4556)? tags_q[0] : 1'b0;
  assign N128 = flush_i;
  assign { tags_n_0__asid__0_, tags_n_0__vpn2__8_, tags_n_0__vpn2__7_, tags_n_0__vpn2__6_, tags_n_0__vpn2__5_, tags_n_0__vpn2__4_, tags_n_0__vpn2__3_, tags_n_0__vpn2__2_, tags_n_0__vpn2__1_, tags_n_0__vpn2__0_, tags_n_0__vpn1__8_, tags_n_0__vpn1__7_, tags_n_0__vpn1__6_, tags_n_0__vpn1__5_, tags_n_0__vpn1__4_, tags_n_0__vpn1__3_, tags_n_0__vpn1__2_, tags_n_0__vpn1__1_, tags_n_0__vpn1__0_, tags_n_0__vpn0__8_, tags_n_0__vpn0__7_, tags_n_0__vpn0__6_, tags_n_0__vpn0__5_, tags_n_0__vpn0__4_, tags_n_0__vpn0__3_, tags_n_0__vpn0__2_, tags_n_0__vpn0__1_, tags_n_0__vpn0__0_, tags_n_0__is_2M_, tags_n_0__is_1G_ } = (N4651)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4556)? tags_q[30:1] : 1'b0;
  assign { content_n_0__reserved__9_, content_n_0__reserved__8_, content_n_0__reserved__7_, content_n_0__reserved__6_, content_n_0__reserved__5_, content_n_0__reserved__4_, content_n_0__reserved__3_, content_n_0__reserved__2_, content_n_0__reserved__1_, content_n_0__reserved__0_, content_n_0__ppn__43_, content_n_0__ppn__42_, content_n_0__ppn__41_, content_n_0__ppn__40_, content_n_0__ppn__39_, content_n_0__ppn__38_, content_n_0__ppn__37_, content_n_0__ppn__36_, content_n_0__ppn__35_, content_n_0__ppn__34_, content_n_0__ppn__33_, content_n_0__ppn__32_, content_n_0__ppn__31_, content_n_0__ppn__30_, content_n_0__ppn__29_, content_n_0__ppn__28_, content_n_0__ppn__27_, content_n_0__ppn__26_, content_n_0__ppn__25_, content_n_0__ppn__24_, content_n_0__ppn__23_, content_n_0__ppn__22_, content_n_0__ppn__21_, content_n_0__ppn__20_, content_n_0__ppn__19_, content_n_0__ppn__18_, content_n_0__ppn__17_, content_n_0__ppn__16_, content_n_0__ppn__15_, content_n_0__ppn__14_, content_n_0__ppn__13_, content_n_0__ppn__12_, content_n_0__ppn__11_, content_n_0__ppn__10_, content_n_0__ppn__9_, content_n_0__ppn__8_, content_n_0__ppn__7_, content_n_0__ppn__6_, content_n_0__ppn__5_, content_n_0__ppn__4_, content_n_0__ppn__3_, content_n_0__ppn__2_, content_n_0__ppn__1_, content_n_0__ppn__0_, content_n_0__rsw__1_, content_n_0__rsw__0_, content_n_0__d_, content_n_0__a_, content_n_0__g_, content_n_0__u_, content_n_0__x_, content_n_0__w_, content_n_0__r_, content_n_0__v_ } = (N4651)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4556)? content_q[63:0] : 1'b0;
  assign tags_n_1__valid_ = (N128)? 1'b0 : 
                            (N4652)? 1'b1 : 
                            (N4562)? tags_q[31] : 1'b0;
  assign { tags_n_1__asid__0_, tags_n_1__vpn2__8_, tags_n_1__vpn2__7_, tags_n_1__vpn2__6_, tags_n_1__vpn2__5_, tags_n_1__vpn2__4_, tags_n_1__vpn2__3_, tags_n_1__vpn2__2_, tags_n_1__vpn2__1_, tags_n_1__vpn2__0_, tags_n_1__vpn1__8_, tags_n_1__vpn1__7_, tags_n_1__vpn1__6_, tags_n_1__vpn1__5_, tags_n_1__vpn1__4_, tags_n_1__vpn1__3_, tags_n_1__vpn1__2_, tags_n_1__vpn1__1_, tags_n_1__vpn1__0_, tags_n_1__vpn0__8_, tags_n_1__vpn0__7_, tags_n_1__vpn0__6_, tags_n_1__vpn0__5_, tags_n_1__vpn0__4_, tags_n_1__vpn0__3_, tags_n_1__vpn0__2_, tags_n_1__vpn0__1_, tags_n_1__vpn0__0_, tags_n_1__is_2M_, tags_n_1__is_1G_ } = (N4652)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4562)? tags_q[61:32] : 1'b0;
  assign { content_n_1__reserved__9_, content_n_1__reserved__8_, content_n_1__reserved__7_, content_n_1__reserved__6_, content_n_1__reserved__5_, content_n_1__reserved__4_, content_n_1__reserved__3_, content_n_1__reserved__2_, content_n_1__reserved__1_, content_n_1__reserved__0_, content_n_1__ppn__43_, content_n_1__ppn__42_, content_n_1__ppn__41_, content_n_1__ppn__40_, content_n_1__ppn__39_, content_n_1__ppn__38_, content_n_1__ppn__37_, content_n_1__ppn__36_, content_n_1__ppn__35_, content_n_1__ppn__34_, content_n_1__ppn__33_, content_n_1__ppn__32_, content_n_1__ppn__31_, content_n_1__ppn__30_, content_n_1__ppn__29_, content_n_1__ppn__28_, content_n_1__ppn__27_, content_n_1__ppn__26_, content_n_1__ppn__25_, content_n_1__ppn__24_, content_n_1__ppn__23_, content_n_1__ppn__22_, content_n_1__ppn__21_, content_n_1__ppn__20_, content_n_1__ppn__19_, content_n_1__ppn__18_, content_n_1__ppn__17_, content_n_1__ppn__16_, content_n_1__ppn__15_, content_n_1__ppn__14_, content_n_1__ppn__13_, content_n_1__ppn__12_, content_n_1__ppn__11_, content_n_1__ppn__10_, content_n_1__ppn__9_, content_n_1__ppn__8_, content_n_1__ppn__7_, content_n_1__ppn__6_, content_n_1__ppn__5_, content_n_1__ppn__4_, content_n_1__ppn__3_, content_n_1__ppn__2_, content_n_1__ppn__1_, content_n_1__ppn__0_, content_n_1__rsw__1_, content_n_1__rsw__0_, content_n_1__d_, content_n_1__a_, content_n_1__g_, content_n_1__u_, content_n_1__x_, content_n_1__w_, content_n_1__r_, content_n_1__v_ } = (N4652)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4562)? content_q[127:64] : 1'b0;
  assign tags_n_2__valid_ = (N128)? 1'b0 : 
                            (N4653)? 1'b1 : 
                            (N4568)? tags_q[62] : 1'b0;
  assign { tags_n_2__asid__0_, tags_n_2__vpn2__8_, tags_n_2__vpn2__7_, tags_n_2__vpn2__6_, tags_n_2__vpn2__5_, tags_n_2__vpn2__4_, tags_n_2__vpn2__3_, tags_n_2__vpn2__2_, tags_n_2__vpn2__1_, tags_n_2__vpn2__0_, tags_n_2__vpn1__8_, tags_n_2__vpn1__7_, tags_n_2__vpn1__6_, tags_n_2__vpn1__5_, tags_n_2__vpn1__4_, tags_n_2__vpn1__3_, tags_n_2__vpn1__2_, tags_n_2__vpn1__1_, tags_n_2__vpn1__0_, tags_n_2__vpn0__8_, tags_n_2__vpn0__7_, tags_n_2__vpn0__6_, tags_n_2__vpn0__5_, tags_n_2__vpn0__4_, tags_n_2__vpn0__3_, tags_n_2__vpn0__2_, tags_n_2__vpn0__1_, tags_n_2__vpn0__0_, tags_n_2__is_2M_, tags_n_2__is_1G_ } = (N4653)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4568)? tags_q[92:63] : 1'b0;
  assign { content_n_2__reserved__9_, content_n_2__reserved__8_, content_n_2__reserved__7_, content_n_2__reserved__6_, content_n_2__reserved__5_, content_n_2__reserved__4_, content_n_2__reserved__3_, content_n_2__reserved__2_, content_n_2__reserved__1_, content_n_2__reserved__0_, content_n_2__ppn__43_, content_n_2__ppn__42_, content_n_2__ppn__41_, content_n_2__ppn__40_, content_n_2__ppn__39_, content_n_2__ppn__38_, content_n_2__ppn__37_, content_n_2__ppn__36_, content_n_2__ppn__35_, content_n_2__ppn__34_, content_n_2__ppn__33_, content_n_2__ppn__32_, content_n_2__ppn__31_, content_n_2__ppn__30_, content_n_2__ppn__29_, content_n_2__ppn__28_, content_n_2__ppn__27_, content_n_2__ppn__26_, content_n_2__ppn__25_, content_n_2__ppn__24_, content_n_2__ppn__23_, content_n_2__ppn__22_, content_n_2__ppn__21_, content_n_2__ppn__20_, content_n_2__ppn__19_, content_n_2__ppn__18_, content_n_2__ppn__17_, content_n_2__ppn__16_, content_n_2__ppn__15_, content_n_2__ppn__14_, content_n_2__ppn__13_, content_n_2__ppn__12_, content_n_2__ppn__11_, content_n_2__ppn__10_, content_n_2__ppn__9_, content_n_2__ppn__8_, content_n_2__ppn__7_, content_n_2__ppn__6_, content_n_2__ppn__5_, content_n_2__ppn__4_, content_n_2__ppn__3_, content_n_2__ppn__2_, content_n_2__ppn__1_, content_n_2__ppn__0_, content_n_2__rsw__1_, content_n_2__rsw__0_, content_n_2__d_, content_n_2__a_, content_n_2__g_, content_n_2__u_, content_n_2__x_, content_n_2__w_, content_n_2__r_, content_n_2__v_ } = (N4653)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4568)? content_q[191:128] : 1'b0;
  assign tags_n_3__valid_ = (N128)? 1'b0 : 
                            (N4654)? 1'b1 : 
                            (N4574)? tags_q[93] : 1'b0;
  assign { tags_n_3__asid__0_, tags_n_3__vpn2__8_, tags_n_3__vpn2__7_, tags_n_3__vpn2__6_, tags_n_3__vpn2__5_, tags_n_3__vpn2__4_, tags_n_3__vpn2__3_, tags_n_3__vpn2__2_, tags_n_3__vpn2__1_, tags_n_3__vpn2__0_, tags_n_3__vpn1__8_, tags_n_3__vpn1__7_, tags_n_3__vpn1__6_, tags_n_3__vpn1__5_, tags_n_3__vpn1__4_, tags_n_3__vpn1__3_, tags_n_3__vpn1__2_, tags_n_3__vpn1__1_, tags_n_3__vpn1__0_, tags_n_3__vpn0__8_, tags_n_3__vpn0__7_, tags_n_3__vpn0__6_, tags_n_3__vpn0__5_, tags_n_3__vpn0__4_, tags_n_3__vpn0__3_, tags_n_3__vpn0__2_, tags_n_3__vpn0__1_, tags_n_3__vpn0__0_, tags_n_3__is_2M_, tags_n_3__is_1G_ } = (N4654)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4574)? tags_q[123:94] : 1'b0;
  assign { content_n_3__reserved__9_, content_n_3__reserved__8_, content_n_3__reserved__7_, content_n_3__reserved__6_, content_n_3__reserved__5_, content_n_3__reserved__4_, content_n_3__reserved__3_, content_n_3__reserved__2_, content_n_3__reserved__1_, content_n_3__reserved__0_, content_n_3__ppn__43_, content_n_3__ppn__42_, content_n_3__ppn__41_, content_n_3__ppn__40_, content_n_3__ppn__39_, content_n_3__ppn__38_, content_n_3__ppn__37_, content_n_3__ppn__36_, content_n_3__ppn__35_, content_n_3__ppn__34_, content_n_3__ppn__33_, content_n_3__ppn__32_, content_n_3__ppn__31_, content_n_3__ppn__30_, content_n_3__ppn__29_, content_n_3__ppn__28_, content_n_3__ppn__27_, content_n_3__ppn__26_, content_n_3__ppn__25_, content_n_3__ppn__24_, content_n_3__ppn__23_, content_n_3__ppn__22_, content_n_3__ppn__21_, content_n_3__ppn__20_, content_n_3__ppn__19_, content_n_3__ppn__18_, content_n_3__ppn__17_, content_n_3__ppn__16_, content_n_3__ppn__15_, content_n_3__ppn__14_, content_n_3__ppn__13_, content_n_3__ppn__12_, content_n_3__ppn__11_, content_n_3__ppn__10_, content_n_3__ppn__9_, content_n_3__ppn__8_, content_n_3__ppn__7_, content_n_3__ppn__6_, content_n_3__ppn__5_, content_n_3__ppn__4_, content_n_3__ppn__3_, content_n_3__ppn__2_, content_n_3__ppn__1_, content_n_3__ppn__0_, content_n_3__rsw__1_, content_n_3__rsw__0_, content_n_3__d_, content_n_3__a_, content_n_3__g_, content_n_3__u_, content_n_3__x_, content_n_3__w_, content_n_3__r_, content_n_3__v_ } = (N4654)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4574)? content_q[255:192] : 1'b0;
  assign tags_n_4__valid_ = (N128)? 1'b0 : 
                            (N4655)? 1'b1 : 
                            (N4580)? tags_q[124] : 1'b0;
  assign { tags_n_4__asid__0_, tags_n_4__vpn2__8_, tags_n_4__vpn2__7_, tags_n_4__vpn2__6_, tags_n_4__vpn2__5_, tags_n_4__vpn2__4_, tags_n_4__vpn2__3_, tags_n_4__vpn2__2_, tags_n_4__vpn2__1_, tags_n_4__vpn2__0_, tags_n_4__vpn1__8_, tags_n_4__vpn1__7_, tags_n_4__vpn1__6_, tags_n_4__vpn1__5_, tags_n_4__vpn1__4_, tags_n_4__vpn1__3_, tags_n_4__vpn1__2_, tags_n_4__vpn1__1_, tags_n_4__vpn1__0_, tags_n_4__vpn0__8_, tags_n_4__vpn0__7_, tags_n_4__vpn0__6_, tags_n_4__vpn0__5_, tags_n_4__vpn0__4_, tags_n_4__vpn0__3_, tags_n_4__vpn0__2_, tags_n_4__vpn0__1_, tags_n_4__vpn0__0_, tags_n_4__is_2M_, tags_n_4__is_1G_ } = (N4655)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4580)? tags_q[154:125] : 1'b0;
  assign { content_n_4__reserved__9_, content_n_4__reserved__8_, content_n_4__reserved__7_, content_n_4__reserved__6_, content_n_4__reserved__5_, content_n_4__reserved__4_, content_n_4__reserved__3_, content_n_4__reserved__2_, content_n_4__reserved__1_, content_n_4__reserved__0_, content_n_4__ppn__43_, content_n_4__ppn__42_, content_n_4__ppn__41_, content_n_4__ppn__40_, content_n_4__ppn__39_, content_n_4__ppn__38_, content_n_4__ppn__37_, content_n_4__ppn__36_, content_n_4__ppn__35_, content_n_4__ppn__34_, content_n_4__ppn__33_, content_n_4__ppn__32_, content_n_4__ppn__31_, content_n_4__ppn__30_, content_n_4__ppn__29_, content_n_4__ppn__28_, content_n_4__ppn__27_, content_n_4__ppn__26_, content_n_4__ppn__25_, content_n_4__ppn__24_, content_n_4__ppn__23_, content_n_4__ppn__22_, content_n_4__ppn__21_, content_n_4__ppn__20_, content_n_4__ppn__19_, content_n_4__ppn__18_, content_n_4__ppn__17_, content_n_4__ppn__16_, content_n_4__ppn__15_, content_n_4__ppn__14_, content_n_4__ppn__13_, content_n_4__ppn__12_, content_n_4__ppn__11_, content_n_4__ppn__10_, content_n_4__ppn__9_, content_n_4__ppn__8_, content_n_4__ppn__7_, content_n_4__ppn__6_, content_n_4__ppn__5_, content_n_4__ppn__4_, content_n_4__ppn__3_, content_n_4__ppn__2_, content_n_4__ppn__1_, content_n_4__ppn__0_, content_n_4__rsw__1_, content_n_4__rsw__0_, content_n_4__d_, content_n_4__a_, content_n_4__g_, content_n_4__u_, content_n_4__x_, content_n_4__w_, content_n_4__r_, content_n_4__v_ } = (N4655)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4580)? content_q[319:256] : 1'b0;
  assign tags_n_5__valid_ = (N128)? 1'b0 : 
                            (N4656)? 1'b1 : 
                            (N4586)? tags_q[155] : 1'b0;
  assign { tags_n_5__asid__0_, tags_n_5__vpn2__8_, tags_n_5__vpn2__7_, tags_n_5__vpn2__6_, tags_n_5__vpn2__5_, tags_n_5__vpn2__4_, tags_n_5__vpn2__3_, tags_n_5__vpn2__2_, tags_n_5__vpn2__1_, tags_n_5__vpn2__0_, tags_n_5__vpn1__8_, tags_n_5__vpn1__7_, tags_n_5__vpn1__6_, tags_n_5__vpn1__5_, tags_n_5__vpn1__4_, tags_n_5__vpn1__3_, tags_n_5__vpn1__2_, tags_n_5__vpn1__1_, tags_n_5__vpn1__0_, tags_n_5__vpn0__8_, tags_n_5__vpn0__7_, tags_n_5__vpn0__6_, tags_n_5__vpn0__5_, tags_n_5__vpn0__4_, tags_n_5__vpn0__3_, tags_n_5__vpn0__2_, tags_n_5__vpn0__1_, tags_n_5__vpn0__0_, tags_n_5__is_2M_, tags_n_5__is_1G_ } = (N4656)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4586)? tags_q[185:156] : 1'b0;
  assign { content_n_5__reserved__9_, content_n_5__reserved__8_, content_n_5__reserved__7_, content_n_5__reserved__6_, content_n_5__reserved__5_, content_n_5__reserved__4_, content_n_5__reserved__3_, content_n_5__reserved__2_, content_n_5__reserved__1_, content_n_5__reserved__0_, content_n_5__ppn__43_, content_n_5__ppn__42_, content_n_5__ppn__41_, content_n_5__ppn__40_, content_n_5__ppn__39_, content_n_5__ppn__38_, content_n_5__ppn__37_, content_n_5__ppn__36_, content_n_5__ppn__35_, content_n_5__ppn__34_, content_n_5__ppn__33_, content_n_5__ppn__32_, content_n_5__ppn__31_, content_n_5__ppn__30_, content_n_5__ppn__29_, content_n_5__ppn__28_, content_n_5__ppn__27_, content_n_5__ppn__26_, content_n_5__ppn__25_, content_n_5__ppn__24_, content_n_5__ppn__23_, content_n_5__ppn__22_, content_n_5__ppn__21_, content_n_5__ppn__20_, content_n_5__ppn__19_, content_n_5__ppn__18_, content_n_5__ppn__17_, content_n_5__ppn__16_, content_n_5__ppn__15_, content_n_5__ppn__14_, content_n_5__ppn__13_, content_n_5__ppn__12_, content_n_5__ppn__11_, content_n_5__ppn__10_, content_n_5__ppn__9_, content_n_5__ppn__8_, content_n_5__ppn__7_, content_n_5__ppn__6_, content_n_5__ppn__5_, content_n_5__ppn__4_, content_n_5__ppn__3_, content_n_5__ppn__2_, content_n_5__ppn__1_, content_n_5__ppn__0_, content_n_5__rsw__1_, content_n_5__rsw__0_, content_n_5__d_, content_n_5__a_, content_n_5__g_, content_n_5__u_, content_n_5__x_, content_n_5__w_, content_n_5__r_, content_n_5__v_ } = (N4656)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4586)? content_q[383:320] : 1'b0;
  assign tags_n_6__valid_ = (N128)? 1'b0 : 
                            (N4657)? 1'b1 : 
                            (N4592)? tags_q[186] : 1'b0;
  assign { tags_n_6__asid__0_, tags_n_6__vpn2__8_, tags_n_6__vpn2__7_, tags_n_6__vpn2__6_, tags_n_6__vpn2__5_, tags_n_6__vpn2__4_, tags_n_6__vpn2__3_, tags_n_6__vpn2__2_, tags_n_6__vpn2__1_, tags_n_6__vpn2__0_, tags_n_6__vpn1__8_, tags_n_6__vpn1__7_, tags_n_6__vpn1__6_, tags_n_6__vpn1__5_, tags_n_6__vpn1__4_, tags_n_6__vpn1__3_, tags_n_6__vpn1__2_, tags_n_6__vpn1__1_, tags_n_6__vpn1__0_, tags_n_6__vpn0__8_, tags_n_6__vpn0__7_, tags_n_6__vpn0__6_, tags_n_6__vpn0__5_, tags_n_6__vpn0__4_, tags_n_6__vpn0__3_, tags_n_6__vpn0__2_, tags_n_6__vpn0__1_, tags_n_6__vpn0__0_, tags_n_6__is_2M_, tags_n_6__is_1G_ } = (N4657)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4592)? tags_q[216:187] : 1'b0;
  assign { content_n_6__reserved__9_, content_n_6__reserved__8_, content_n_6__reserved__7_, content_n_6__reserved__6_, content_n_6__reserved__5_, content_n_6__reserved__4_, content_n_6__reserved__3_, content_n_6__reserved__2_, content_n_6__reserved__1_, content_n_6__reserved__0_, content_n_6__ppn__43_, content_n_6__ppn__42_, content_n_6__ppn__41_, content_n_6__ppn__40_, content_n_6__ppn__39_, content_n_6__ppn__38_, content_n_6__ppn__37_, content_n_6__ppn__36_, content_n_6__ppn__35_, content_n_6__ppn__34_, content_n_6__ppn__33_, content_n_6__ppn__32_, content_n_6__ppn__31_, content_n_6__ppn__30_, content_n_6__ppn__29_, content_n_6__ppn__28_, content_n_6__ppn__27_, content_n_6__ppn__26_, content_n_6__ppn__25_, content_n_6__ppn__24_, content_n_6__ppn__23_, content_n_6__ppn__22_, content_n_6__ppn__21_, content_n_6__ppn__20_, content_n_6__ppn__19_, content_n_6__ppn__18_, content_n_6__ppn__17_, content_n_6__ppn__16_, content_n_6__ppn__15_, content_n_6__ppn__14_, content_n_6__ppn__13_, content_n_6__ppn__12_, content_n_6__ppn__11_, content_n_6__ppn__10_, content_n_6__ppn__9_, content_n_6__ppn__8_, content_n_6__ppn__7_, content_n_6__ppn__6_, content_n_6__ppn__5_, content_n_6__ppn__4_, content_n_6__ppn__3_, content_n_6__ppn__2_, content_n_6__ppn__1_, content_n_6__ppn__0_, content_n_6__rsw__1_, content_n_6__rsw__0_, content_n_6__d_, content_n_6__a_, content_n_6__g_, content_n_6__u_, content_n_6__x_, content_n_6__w_, content_n_6__r_, content_n_6__v_ } = (N4657)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4592)? content_q[447:384] : 1'b0;
  assign tags_n_7__valid_ = (N128)? 1'b0 : 
                            (N4658)? 1'b1 : 
                            (N4598)? tags_q[217] : 1'b0;
  assign { tags_n_7__asid__0_, tags_n_7__vpn2__8_, tags_n_7__vpn2__7_, tags_n_7__vpn2__6_, tags_n_7__vpn2__5_, tags_n_7__vpn2__4_, tags_n_7__vpn2__3_, tags_n_7__vpn2__2_, tags_n_7__vpn2__1_, tags_n_7__vpn2__0_, tags_n_7__vpn1__8_, tags_n_7__vpn1__7_, tags_n_7__vpn1__6_, tags_n_7__vpn1__5_, tags_n_7__vpn1__4_, tags_n_7__vpn1__3_, tags_n_7__vpn1__2_, tags_n_7__vpn1__1_, tags_n_7__vpn1__0_, tags_n_7__vpn0__8_, tags_n_7__vpn0__7_, tags_n_7__vpn0__6_, tags_n_7__vpn0__5_, tags_n_7__vpn0__4_, tags_n_7__vpn0__3_, tags_n_7__vpn0__2_, tags_n_7__vpn0__1_, tags_n_7__vpn0__0_, tags_n_7__is_2M_, tags_n_7__is_1G_ } = (N4658)? { update_i[64:64], update_i[91:65], update_i[93:92] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  (N4598)? tags_q[247:218] : 1'b0;
  assign { content_n_7__reserved__9_, content_n_7__reserved__8_, content_n_7__reserved__7_, content_n_7__reserved__6_, content_n_7__reserved__5_, content_n_7__reserved__4_, content_n_7__reserved__3_, content_n_7__reserved__2_, content_n_7__reserved__1_, content_n_7__reserved__0_, content_n_7__ppn__43_, content_n_7__ppn__42_, content_n_7__ppn__41_, content_n_7__ppn__40_, content_n_7__ppn__39_, content_n_7__ppn__38_, content_n_7__ppn__37_, content_n_7__ppn__36_, content_n_7__ppn__35_, content_n_7__ppn__34_, content_n_7__ppn__33_, content_n_7__ppn__32_, content_n_7__ppn__31_, content_n_7__ppn__30_, content_n_7__ppn__29_, content_n_7__ppn__28_, content_n_7__ppn__27_, content_n_7__ppn__26_, content_n_7__ppn__25_, content_n_7__ppn__24_, content_n_7__ppn__23_, content_n_7__ppn__22_, content_n_7__ppn__21_, content_n_7__ppn__20_, content_n_7__ppn__19_, content_n_7__ppn__18_, content_n_7__ppn__17_, content_n_7__ppn__16_, content_n_7__ppn__15_, content_n_7__ppn__14_, content_n_7__ppn__13_, content_n_7__ppn__12_, content_n_7__ppn__11_, content_n_7__ppn__10_, content_n_7__ppn__9_, content_n_7__ppn__8_, content_n_7__ppn__7_, content_n_7__ppn__6_, content_n_7__ppn__5_, content_n_7__ppn__4_, content_n_7__ppn__3_, content_n_7__ppn__2_, content_n_7__ppn__1_, content_n_7__ppn__0_, content_n_7__rsw__1_, content_n_7__rsw__0_, content_n_7__d_, content_n_7__a_, content_n_7__g_, content_n_7__u_, content_n_7__x_, content_n_7__w_, content_n_7__r_, content_n_7__v_ } = (N4658)? update_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N4598)? content_q[511:448] : 1'b0;
  assign tags_n_8__valid_ = (N128)? 1'b0 : 
                            (N4659)? 1'b1 : 1'b0;
  assign tags_n_9__valid_ = (N128)? 1'b0 : 
                            (N4660)? 1'b1 : 1'b0;
  assign tags_n_10__valid_ = (N128)? 1'b0 : 
                             (N4661)? 1'b1 : 1'b0;
  assign tags_n_11__valid_ = (N128)? 1'b0 : 
                             (N4662)? 1'b1 : 1'b0;
  assign tags_n_12__valid_ = (N128)? 1'b0 : 
                             (N4663)? 1'b1 : 1'b0;
  assign tags_n_13__valid_ = (N128)? 1'b0 : 
                             (N4664)? 1'b1 : 1'b0;
  assign tags_n_14__valid_ = (N128)? 1'b0 : 
                             (N4665)? 1'b1 : 1'b0;
  assign tags_n_15__valid_ = (N128)? 1'b0 : 
                             (N4666)? 1'b1 : 1'b0;
  assign { N4672, N4671, N4670, N4669 } = (N129)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                          (N4668)? { plru_tree_q[7:7], plru_tree_q[3:3], plru_tree_q[1:0] } : 1'b0;
  assign N129 = N4667;
  assign { plru_tree_n[7:7], N4677, N4676, N4675 } = (N130)? { 1'b0, 1'b1, 1'b1, 1'b1 } : 
                                                     (N4674)? { N4672, N4671, N4670, N4669 } : 1'b0;
  assign N130 = N4673;
  assign { N4683, N4682, N4681, N4680 } = (N131)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                                          (N4679)? { plru_tree_q[8:8], N4677, N4676, N4675 } : 1'b0;
  assign N131 = N4678;
  assign { plru_tree_n[8:8], plru_tree_n[3:3], N4687, N4686 } = (N132)? { 1'b0, 1'b0, 1'b1, 1'b1 } : 
                                                                (N4685)? { N4683, N4682, N4681, N4680 } : 1'b0;
  assign N132 = N4684;
  assign { N4693, N4692, N4691, N4690 } = (N133)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                                          (N4689)? { plru_tree_q[9:9], plru_tree_q[4:4], N4687, N4686 } : 1'b0;
  assign N133 = N4688;
  assign { plru_tree_n[9:9], N4698, N4697, N4696 } = (N134)? { 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                     (N4695)? { N4693, N4692, N4691, N4690 } : 1'b0;
  assign N134 = N4694;
  assign { N4704, N4703, N4702, N4701 } = (N135)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                                          (N4700)? { plru_tree_q[10:10], N4698, N4697, N4696 } : 1'b0;
  assign N135 = N4699;
  assign { plru_tree_n[10:10], plru_tree_n[4:4], plru_tree_n[1:1], N4707 } = (N136)? { 1'b0, 1'b0, 1'b0, 1'b1 } : 
                                                                             (N4706)? { N4704, N4703, N4702, N4701 } : 1'b0;
  assign N136 = N4705;
  assign { N4713, N4712, N4711, N4710 } = (N137)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                                          (N4709)? { plru_tree_q[11:11], plru_tree_q[5:5], plru_tree_q[2:2], N4707 } : 1'b0;
  assign N137 = N4708;
  assign { plru_tree_n[11:11], N4718, N4717, N4716 } = (N138)? { 1'b0, 1'b1, 1'b1, 1'b0 } : 
                                                       (N4715)? { N4713, N4712, N4711, N4710 } : 1'b0;
  assign N138 = N4714;
  assign { N4724, N4723, N4722, N4721 } = (N139)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                          (N4720)? { plru_tree_q[12:12], N4718, N4717, N4716 } : 1'b0;
  assign N139 = N4719;
  assign { plru_tree_n[12:12], plru_tree_n[5:5], N4728, N4727 } = (N140)? { 1'b0, 1'b0, 1'b1, 1'b0 } : 
                                                                  (N4726)? { N4724, N4723, N4722, N4721 } : 1'b0;
  assign N140 = N4725;
  assign { N4734, N4733, N4732, N4731 } = (N141)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                                          (N4730)? { plru_tree_q[13:13], plru_tree_q[6:6], N4728, N4727 } : 1'b0;
  assign N141 = N4729;
  assign { plru_tree_n[13:13], N4739, N4738, N4737 } = (N142)? { 1'b0, 1'b1, 1'b0, 1'b0 } : 
                                                       (N4736)? { N4734, N4733, N4732, N4731 } : 1'b0;
  assign N142 = N4735;
  assign { N4745, N4744, N4743, N4742 } = (N143)? { 1'b1, 1'b0, 1'b0, 1'b0 } : 
                                          (N4741)? { plru_tree_q[14:14], N4739, N4738, N4737 } : 1'b0;
  assign N143 = N4740;
  assign { plru_tree_n[14:14], plru_tree_n[6:6], plru_tree_n[2:2], plru_tree_n[0:0] } = (N144)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                        (N4747)? { N4745, N4744, N4743, N4742 } : 1'b0;
  assign N144 = N4746;
  assign N147 = N4839 & N146;
  assign N4839 = tags_q[0] & N145;
  assign N148 = ~N147;
  assign N149 = N147;
  assign N150 = ~tags_q[1];
  assign N151 = N149 & N150;
  assign N153 = ~N152;
  assign N155 = tags_q[2] | N154;
  assign N156 = ~N155;
  assign N423 = N4840 & N422;
  assign N4840 = tags_q[31] & N421;
  assign N424 = ~N423;
  assign N425 = N423;
  assign N426 = ~tags_q[32];
  assign N427 = N425 & N426;
  assign N429 = ~N428;
  assign N431 = tags_q[33] | N430;
  assign N432 = ~N431;
  assign N703 = N4841 & N702;
  assign N4841 = tags_q[62] & N701;
  assign N704 = ~N703;
  assign N705 = N703;
  assign N706 = ~tags_q[63];
  assign N707 = N705 & N706;
  assign N709 = ~N708;
  assign N711 = tags_q[64] | N710;
  assign N712 = ~N711;
  assign N983 = N4842 & N982;
  assign N4842 = tags_q[93] & N981;
  assign N984 = ~N983;
  assign N985 = N983;
  assign N986 = ~tags_q[94];
  assign N987 = N985 & N986;
  assign N989 = ~N988;
  assign N991 = tags_q[95] | N990;
  assign N992 = ~N991;
  assign N1263 = N4843 & N1262;
  assign N4843 = tags_q[124] & N1261;
  assign N1264 = ~N1263;
  assign N1265 = N1263;
  assign N1266 = ~tags_q[125];
  assign N1267 = N1265 & N1266;
  assign N1269 = ~N1268;
  assign N1271 = tags_q[126] | N1270;
  assign N1272 = ~N1271;
  assign N1543 = N4844 & N1542;
  assign N4844 = tags_q[155] & N1541;
  assign N1544 = ~N1543;
  assign N1545 = N1543;
  assign N1546 = ~tags_q[156];
  assign N1547 = N1545 & N1546;
  assign N1549 = ~N1548;
  assign N1551 = tags_q[157] | N1550;
  assign N1552 = ~N1551;
  assign N1823 = N4845 & N1822;
  assign N4845 = tags_q[186] & N1821;
  assign N1824 = ~N1823;
  assign N1825 = N1823;
  assign N1826 = ~tags_q[187];
  assign N1827 = N1825 & N1826;
  assign N1829 = ~N1828;
  assign N1831 = tags_q[188] | N1830;
  assign N1832 = ~N1831;
  assign N2103 = N4846 & N2102;
  assign N4846 = tags_q[217] & N2101;
  assign N2104 = ~N2103;
  assign N2105 = N2103;
  assign N2106 = ~tags_q[218];
  assign N2107 = N2105 & N2106;
  assign N2109 = ~N2108;
  assign N2111 = tags_q[219] | N2110;
  assign N2112 = ~N2111;
  assign N2383 = N4847 & N2382;
  assign N4847 = tags_q[248] & N2381;
  assign N2384 = ~N2383;
  assign N2385 = N2383;
  assign N2386 = ~tags_q[249];
  assign N2387 = N2385 & N2386;
  assign N2389 = ~N2388;
  assign N2391 = tags_q[250] | N2390;
  assign N2392 = ~N2391;
  assign N2663 = N4848 & N2662;
  assign N4848 = tags_q[279] & N2661;
  assign N2664 = ~N2663;
  assign N2665 = N2663;
  assign N2666 = ~tags_q[280];
  assign N2667 = N2665 & N2666;
  assign N2669 = ~N2668;
  assign N2671 = tags_q[281] | N2670;
  assign N2672 = ~N2671;
  assign N2943 = N4849 & N2942;
  assign N4849 = tags_q[310] & N2941;
  assign N2944 = ~N2943;
  assign N2945 = N2943;
  assign N2946 = ~tags_q[311];
  assign N2947 = N2945 & N2946;
  assign N2949 = ~N2948;
  assign N2951 = tags_q[312] | N2950;
  assign N2952 = ~N2951;
  assign N3223 = N4850 & N3222;
  assign N4850 = tags_q[341] & N3221;
  assign N3224 = ~N3223;
  assign N3225 = N3223;
  assign N3226 = ~tags_q[342];
  assign N3227 = N3225 & N3226;
  assign N3229 = ~N3228;
  assign N3231 = tags_q[343] | N3230;
  assign N3232 = ~N3231;
  assign N3503 = N4851 & N3502;
  assign N4851 = tags_q[372] & N3501;
  assign N3504 = ~N3503;
  assign N3505 = N3503;
  assign N3506 = ~tags_q[373];
  assign N3507 = N3505 & N3506;
  assign N3509 = ~N3508;
  assign N3511 = tags_q[374] | N3510;
  assign N3512 = ~N3511;
  assign N3783 = N4852 & N3782;
  assign N4852 = tags_q[403] & N3781;
  assign N3784 = ~N3783;
  assign N3785 = N3783;
  assign N3786 = ~tags_q[404];
  assign N3787 = N3785 & N3786;
  assign N3789 = ~N3788;
  assign N3791 = tags_q[405] | N3790;
  assign N3792 = ~N3791;
  assign N4063 = N4853 & N4062;
  assign N4853 = tags_q[434] & N4061;
  assign N4064 = ~N4063;
  assign N4065 = N4063;
  assign N4066 = ~tags_q[435];
  assign N4067 = N4065 & N4066;
  assign N4069 = ~N4068;
  assign N4071 = tags_q[436] | N4070;
  assign N4072 = ~N4071;
  assign N4343 = N4854 & N4342;
  assign N4854 = tags_q[465] & N4341;
  assign N4344 = ~N4343;
  assign N4345 = N4343;
  assign N4346 = ~tags_q[466];
  assign N4347 = N4345 & N4346;
  assign N4349 = ~N4348;
  assign N4351 = tags_q[467] | N4350;
  assign N4352 = ~N4351;
  assign N4554 = update_i[94] & replace_en[0];
  assign N4555 = N4554 | flush_i;
  assign N4556 = ~N4555;
  assign N4558 = N4557 | N4838;
  assign N4559 = ~N4558;
  assign N4560 = update_i[94] & replace_en[1];
  assign N4561 = N4560 | flush_i;
  assign N4562 = ~N4561;
  assign N4564 = N4563 | N4838;
  assign N4565 = ~N4564;
  assign N4566 = update_i[94] & replace_en[2];
  assign N4567 = N4566 | flush_i;
  assign N4568 = ~N4567;
  assign N4570 = N4569 | N4838;
  assign N4571 = ~N4570;
  assign N4572 = update_i[94] & replace_en[3];
  assign N4573 = N4572 | flush_i;
  assign N4574 = ~N4573;
  assign N4576 = N4575 | N4838;
  assign N4577 = ~N4576;
  assign N4578 = update_i[94] & replace_en[4];
  assign N4579 = N4578 | flush_i;
  assign N4580 = ~N4579;
  assign N4582 = N4581 | N4838;
  assign N4583 = ~N4582;
  assign N4584 = update_i[94] & replace_en[5];
  assign N4585 = N4584 | flush_i;
  assign N4586 = ~N4585;
  assign N4588 = N4587 | N4838;
  assign N4589 = ~N4588;
  assign N4590 = update_i[94] & replace_en[6];
  assign N4591 = N4590 | flush_i;
  assign N4592 = ~N4591;
  assign N4594 = N4593 | N4838;
  assign N4595 = ~N4594;
  assign N4596 = update_i[94] & replace_en[7];
  assign N4597 = N4596 | flush_i;
  assign N4598 = ~N4597;
  assign N4600 = N4599 | N4838;
  assign N4601 = ~N4600;
  assign N4602 = update_i[94] & replace_en[8];
  assign N4603 = N4602 | flush_i;
  assign N4604 = ~N4603;
  assign N4606 = N4605 | N4838;
  assign N4607 = ~N4606;
  assign N4608 = update_i[94] & replace_en[9];
  assign N4609 = N4608 | flush_i;
  assign N4610 = ~N4609;
  assign N4612 = N4611 | N4838;
  assign N4613 = ~N4612;
  assign N4614 = update_i[94] & replace_en[10];
  assign N4615 = N4614 | flush_i;
  assign N4616 = ~N4615;
  assign N4618 = N4617 | N4838;
  assign N4619 = ~N4618;
  assign N4620 = update_i[94] & replace_en[11];
  assign N4621 = N4620 | flush_i;
  assign N4622 = ~N4621;
  assign N4624 = N4623 | N4838;
  assign N4625 = ~N4624;
  assign N4626 = update_i[94] & replace_en[12];
  assign N4627 = N4626 | flush_i;
  assign N4628 = ~N4627;
  assign N4630 = N4629 | N4838;
  assign N4631 = ~N4630;
  assign N4632 = update_i[94] & replace_en[13];
  assign N4633 = N4632 | flush_i;
  assign N4634 = ~N4633;
  assign N4636 = N4635 | N4838;
  assign N4637 = ~N4636;
  assign N4638 = update_i[94] & replace_en[14];
  assign N4639 = N4638 | flush_i;
  assign N4640 = ~N4639;
  assign N4642 = N4641 | N4838;
  assign N4643 = ~N4642;
  assign N4644 = update_i[94] & replace_en[15];
  assign N4645 = N4644 | flush_i;
  assign N4646 = ~N4645;
  assign N4648 = N4647 | N4838;
  assign N4649 = ~N4648;
  assign N4650 = ~flush_i;
  assign N4651 = N4554 & N4650;
  assign N4652 = N4560 & N4650;
  assign N4653 = N4566 & N4650;
  assign N4654 = N4572 & N4650;
  assign N4655 = N4578 & N4650;
  assign N4656 = N4584 & N4650;
  assign N4657 = N4590 & N4650;
  assign N4658 = N4596 & N4650;
  assign N4659 = N4602 & N4650;
  assign N4660 = N4608 & N4650;
  assign N4661 = N4614 & N4650;
  assign N4662 = N4620 & N4650;
  assign N4663 = N4626 & N4650;
  assign N4664 = N4632 & N4650;
  assign N4665 = N4638 & N4650;
  assign N4666 = N4644 & N4650;
  assign N4667 = lu_hit[0] & lu_access_i;
  assign N4668 = ~N4667;
  assign N4673 = lu_hit[1] & lu_access_i;
  assign N4674 = ~N4673;
  assign N4678 = lu_hit[2] & lu_access_i;
  assign N4679 = ~N4678;
  assign N4684 = lu_hit[3] & lu_access_i;
  assign N4685 = ~N4684;
  assign N4688 = lu_hit[4] & lu_access_i;
  assign N4689 = ~N4688;
  assign N4694 = lu_hit[5] & lu_access_i;
  assign N4695 = ~N4694;
  assign N4699 = lu_hit[6] & lu_access_i;
  assign N4700 = ~N4699;
  assign N4705 = lu_hit[7] & lu_access_i;
  assign N4706 = ~N4705;
  assign N4708 = lu_hit[8] & lu_access_i;
  assign N4709 = ~N4708;
  assign N4714 = lu_hit[9] & lu_access_i;
  assign N4715 = ~N4714;
  assign N4719 = lu_hit[10] & lu_access_i;
  assign N4720 = ~N4719;
  assign N4725 = lu_hit[11] & lu_access_i;
  assign N4726 = ~N4725;
  assign N4729 = lu_hit[12] & lu_access_i;
  assign N4730 = ~N4729;
  assign N4735 = lu_hit[13] & lu_access_i;
  assign N4736 = ~N4735;
  assign N4740 = lu_hit[14] & lu_access_i;
  assign N4741 = ~N4740;
  assign N4746 = lu_hit[15] & lu_access_i;
  assign N4747 = ~N4746;
  assign N4748 = ~plru_tree_q[0];
  assign N4749 = N4748 & N4855;
  assign N4855 = ~plru_tree_q[1];
  assign N4750 = N4749 & N4856;
  assign N4856 = ~plru_tree_q[3];
  assign replace_en[0] = N4750 & N4857;
  assign N4857 = ~plru_tree_q[7];
  assign N4751 = N4748 & N4855;
  assign N4752 = N4751 & N4856;
  assign replace_en[1] = N4752 & plru_tree_q[7];
  assign N4753 = N4748 & N4855;
  assign N4754 = N4753 & plru_tree_q[3];
  assign replace_en[2] = N4754 & N4858;
  assign N4858 = ~plru_tree_q[8];
  assign N4755 = N4748 & N4855;
  assign N4756 = N4755 & plru_tree_q[3];
  assign replace_en[3] = N4756 & plru_tree_q[8];
  assign N4757 = N4748 & plru_tree_q[1];
  assign N4758 = N4757 & N4859;
  assign N4859 = ~plru_tree_q[4];
  assign replace_en[4] = N4758 & N4860;
  assign N4860 = ~plru_tree_q[9];
  assign N4759 = N4748 & plru_tree_q[1];
  assign N4760 = N4759 & N4859;
  assign replace_en[5] = N4760 & plru_tree_q[9];
  assign N4761 = N4748 & plru_tree_q[1];
  assign N4762 = N4761 & plru_tree_q[4];
  assign replace_en[6] = N4762 & N4861;
  assign N4861 = ~plru_tree_q[10];
  assign N4763 = N4748 & plru_tree_q[1];
  assign N4764 = N4763 & plru_tree_q[4];
  assign replace_en[7] = N4764 & plru_tree_q[10];
  assign N4765 = plru_tree_q[0] & N4862;
  assign N4862 = ~plru_tree_q[2];
  assign N4766 = N4765 & N4863;
  assign N4863 = ~plru_tree_q[5];
  assign replace_en[8] = N4766 & N4864;
  assign N4864 = ~plru_tree_q[11];
  assign N4767 = plru_tree_q[0] & N4862;
  assign N4768 = N4767 & N4863;
  assign replace_en[9] = N4768 & plru_tree_q[11];
  assign N4769 = plru_tree_q[0] & N4862;
  assign N4770 = N4769 & plru_tree_q[5];
  assign replace_en[10] = N4770 & N4865;
  assign N4865 = ~plru_tree_q[12];
  assign N4771 = plru_tree_q[0] & N4862;
  assign N4772 = N4771 & plru_tree_q[5];
  assign replace_en[11] = N4772 & plru_tree_q[12];
  assign N4773 = plru_tree_q[0] & plru_tree_q[2];
  assign N4774 = N4773 & N4866;
  assign N4866 = ~plru_tree_q[6];
  assign replace_en[12] = N4774 & N4867;
  assign N4867 = ~plru_tree_q[13];
  assign N4775 = plru_tree_q[0] & plru_tree_q[2];
  assign N4776 = N4775 & N4866;
  assign replace_en[13] = N4776 & plru_tree_q[13];
  assign N4777 = plru_tree_q[0] & plru_tree_q[2];
  assign N4778 = N4777 & plru_tree_q[6];
  assign replace_en[14] = N4778 & N4868;
  assign N4868 = ~plru_tree_q[14];
  assign N4779 = plru_tree_q[0] & plru_tree_q[2];
  assign N4780 = N4779 & plru_tree_q[6];
  assign replace_en[15] = N4780 & plru_tree_q[14];
  assign N4781 = ~rst_ni;
  assign N4782 = flush_i | N4646;
  assign N4783 = ~N4782;
  assign N4784 = N4649 & flush_i;
  assign N4785 = N4784 | N4646;
  assign N4786 = ~N4785;
  assign N4787 = flush_i | N4640;
  assign N4788 = ~N4787;
  assign N4789 = N4643 & flush_i;
  assign N4790 = N4789 | N4640;
  assign N4791 = ~N4790;
  assign N4792 = flush_i | N4634;
  assign N4793 = ~N4792;
  assign N4794 = N4637 & flush_i;
  assign N4795 = N4794 | N4634;
  assign N4796 = ~N4795;
  assign N4797 = flush_i | N4628;
  assign N4798 = ~N4797;
  assign N4799 = N4631 & flush_i;
  assign N4800 = N4799 | N4628;
  assign N4801 = ~N4800;
  assign N4802 = flush_i | N4622;
  assign N4803 = ~N4802;
  assign N4804 = N4625 & flush_i;
  assign N4805 = N4804 | N4622;
  assign N4806 = ~N4805;
  assign N4807 = flush_i | N4616;
  assign N4808 = ~N4807;
  assign N4809 = N4619 & flush_i;
  assign N4810 = N4809 | N4616;
  assign N4811 = ~N4810;
  assign N4812 = flush_i | N4610;
  assign N4813 = ~N4812;
  assign N4814 = N4613 & flush_i;
  assign N4815 = N4814 | N4610;
  assign N4816 = ~N4815;
  assign N4817 = flush_i | N4604;
  assign N4818 = ~N4817;
  assign N4819 = N4607 & flush_i;
  assign N4820 = N4819 | N4604;
  assign N4821 = ~N4820;
  assign N4822 = N4601 & flush_i;
  assign N4823 = ~N4822;
  assign N4824 = N4595 & flush_i;
  assign N4825 = ~N4824;
  assign N4826 = N4589 & flush_i;
  assign N4827 = ~N4826;
  assign N4828 = N4583 & flush_i;
  assign N4829 = ~N4828;
  assign N4830 = N4577 & flush_i;
  assign N4831 = ~N4830;
  assign N4832 = N4571 & flush_i;
  assign N4833 = ~N4832;
  assign N4834 = N4565 & flush_i;
  assign N4835 = ~N4834;
  assign N4836 = N4559 & flush_i;
  assign N4837 = ~N4836;

endmodule