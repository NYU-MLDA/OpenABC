module bsg_buf_ctrl_width_p33
(
  i,
  o
);

  output [32:0] o;
  input i;
  wire [32:0] o;
  wire i;
  assign o[0] = i;
  assign o[1] = i;
  assign o[2] = i;
  assign o[3] = i;
  assign o[4] = i;
  assign o[5] = i;
  assign o[6] = i;
  assign o[7] = i;
  assign o[8] = i;
  assign o[9] = i;
  assign o[10] = i;
  assign o[11] = i;
  assign o[12] = i;
  assign o[13] = i;
  assign o[14] = i;
  assign o[15] = i;
  assign o[16] = i;
  assign o[17] = i;
  assign o[18] = i;
  assign o[19] = i;
  assign o[20] = i;
  assign o[21] = i;
  assign o[22] = i;
  assign o[23] = i;
  assign o[24] = i;
  assign o[25] = i;
  assign o[26] = i;
  assign o[27] = i;
  assign o[28] = i;
  assign o[29] = i;
  assign o[30] = i;
  assign o[31] = i;
  assign o[32] = i;

endmodule