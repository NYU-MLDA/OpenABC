module fifo_v3_0_00000020_00000008
(
  clk_i,
  rst_ni,
  flush_i,
  testmode_i,
  full_o,
  empty_o,
  usage_o,
  data_i,
  push_i,
  data_o,
  pop_i
);

  output [2:0] usage_o;
  input [166:0] data_i;
  output [166:0] data_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input testmode_i;
  input push_i;
  input pop_i;
  output full_o;
  output empty_o;
  wire [166:0] data_o;
  wire full_o,empty_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,
  N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,
  N38,gate_clock,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,
  N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,
  N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,
  N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,
  N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,
  N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,
  N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,
  N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,
  N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,
  N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,
  N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,
  N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
  N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,
  N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,
  N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,
  N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,
  N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,
  N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,
  N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,
  N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,
  N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,
  N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,
  N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,
  N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,
  N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,
  N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,
  N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,
  N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,
  N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,
  N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,
  N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,
  N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,
  N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,
  N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
  N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,
  N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,
  N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,
  N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,
  N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,
  N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,
  N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,
  N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,
  N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,
  N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,
  N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,
  N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,
  N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,
  N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,
  N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,
  N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,
  N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,
  N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,
  N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,
  N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,
  N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,
  N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,
  N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,
  N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,
  N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,
  N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,
  N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,
  N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,
  N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,
  N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,
  N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,
  N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,
  N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,
  N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,
  N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,
  N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,
  N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,
  N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,
  N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,
  N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,
  N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,
  N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,
  N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,
  N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,
  N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,
  N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,
  N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1442,N1443,N1444,N1445,N1447,N1448,
  N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456;
  wire [1335:0] mem_n;
  reg [3:3] status_cnt_q;
  reg [2:0] usage_o,read_pointer_q,write_pointer_q;
  reg [1335:0] mem_q;
  assign data_o[166] = (N31)? mem_q[166] : 
                       (N33)? mem_q[333] : 
                       (N35)? mem_q[500] : 
                       (N37)? mem_q[667] : 
                       (N32)? mem_q[834] : 
                       (N34)? mem_q[1001] : 
                       (N36)? mem_q[1168] : 
                       (N38)? mem_q[1335] : 1'b0;
  assign data_o[165] = (N31)? mem_q[165] : 
                       (N33)? mem_q[332] : 
                       (N35)? mem_q[499] : 
                       (N37)? mem_q[666] : 
                       (N32)? mem_q[833] : 
                       (N34)? mem_q[1000] : 
                       (N36)? mem_q[1167] : 
                       (N38)? mem_q[1334] : 1'b0;
  assign data_o[164] = (N31)? mem_q[164] : 
                       (N33)? mem_q[331] : 
                       (N35)? mem_q[498] : 
                       (N37)? mem_q[665] : 
                       (N32)? mem_q[832] : 
                       (N34)? mem_q[999] : 
                       (N36)? mem_q[1166] : 
                       (N38)? mem_q[1333] : 1'b0;
  assign data_o[163] = (N31)? mem_q[163] : 
                       (N33)? mem_q[330] : 
                       (N35)? mem_q[497] : 
                       (N37)? mem_q[664] : 
                       (N32)? mem_q[831] : 
                       (N34)? mem_q[998] : 
                       (N36)? mem_q[1165] : 
                       (N38)? mem_q[1332] : 1'b0;
  assign data_o[162] = (N31)? mem_q[162] : 
                       (N33)? mem_q[329] : 
                       (N35)? mem_q[496] : 
                       (N37)? mem_q[663] : 
                       (N32)? mem_q[830] : 
                       (N34)? mem_q[997] : 
                       (N36)? mem_q[1164] : 
                       (N38)? mem_q[1331] : 1'b0;
  assign data_o[161] = (N31)? mem_q[161] : 
                       (N33)? mem_q[328] : 
                       (N35)? mem_q[495] : 
                       (N37)? mem_q[662] : 
                       (N32)? mem_q[829] : 
                       (N34)? mem_q[996] : 
                       (N36)? mem_q[1163] : 
                       (N38)? mem_q[1330] : 1'b0;
  assign data_o[160] = (N31)? mem_q[160] : 
                       (N33)? mem_q[327] : 
                       (N35)? mem_q[494] : 
                       (N37)? mem_q[661] : 
                       (N32)? mem_q[828] : 
                       (N34)? mem_q[995] : 
                       (N36)? mem_q[1162] : 
                       (N38)? mem_q[1329] : 1'b0;
  assign data_o[159] = (N31)? mem_q[159] : 
                       (N33)? mem_q[326] : 
                       (N35)? mem_q[493] : 
                       (N37)? mem_q[660] : 
                       (N32)? mem_q[827] : 
                       (N34)? mem_q[994] : 
                       (N36)? mem_q[1161] : 
                       (N38)? mem_q[1328] : 1'b0;
  assign data_o[158] = (N31)? mem_q[158] : 
                       (N33)? mem_q[325] : 
                       (N35)? mem_q[492] : 
                       (N37)? mem_q[659] : 
                       (N32)? mem_q[826] : 
                       (N34)? mem_q[993] : 
                       (N36)? mem_q[1160] : 
                       (N38)? mem_q[1327] : 1'b0;
  assign data_o[157] = (N31)? mem_q[157] : 
                       (N33)? mem_q[324] : 
                       (N35)? mem_q[491] : 
                       (N37)? mem_q[658] : 
                       (N32)? mem_q[825] : 
                       (N34)? mem_q[992] : 
                       (N36)? mem_q[1159] : 
                       (N38)? mem_q[1326] : 1'b0;
  assign data_o[156] = (N31)? mem_q[156] : 
                       (N33)? mem_q[323] : 
                       (N35)? mem_q[490] : 
                       (N37)? mem_q[657] : 
                       (N32)? mem_q[824] : 
                       (N34)? mem_q[991] : 
                       (N36)? mem_q[1158] : 
                       (N38)? mem_q[1325] : 1'b0;
  assign data_o[155] = (N31)? mem_q[155] : 
                       (N33)? mem_q[322] : 
                       (N35)? mem_q[489] : 
                       (N37)? mem_q[656] : 
                       (N32)? mem_q[823] : 
                       (N34)? mem_q[990] : 
                       (N36)? mem_q[1157] : 
                       (N38)? mem_q[1324] : 1'b0;
  assign data_o[154] = (N31)? mem_q[154] : 
                       (N33)? mem_q[321] : 
                       (N35)? mem_q[488] : 
                       (N37)? mem_q[655] : 
                       (N32)? mem_q[822] : 
                       (N34)? mem_q[989] : 
                       (N36)? mem_q[1156] : 
                       (N38)? mem_q[1323] : 1'b0;
  assign data_o[153] = (N31)? mem_q[153] : 
                       (N33)? mem_q[320] : 
                       (N35)? mem_q[487] : 
                       (N37)? mem_q[654] : 
                       (N32)? mem_q[821] : 
                       (N34)? mem_q[988] : 
                       (N36)? mem_q[1155] : 
                       (N38)? mem_q[1322] : 1'b0;
  assign data_o[152] = (N31)? mem_q[152] : 
                       (N33)? mem_q[319] : 
                       (N35)? mem_q[486] : 
                       (N37)? mem_q[653] : 
                       (N32)? mem_q[820] : 
                       (N34)? mem_q[987] : 
                       (N36)? mem_q[1154] : 
                       (N38)? mem_q[1321] : 1'b0;
  assign data_o[151] = (N31)? mem_q[151] : 
                       (N33)? mem_q[318] : 
                       (N35)? mem_q[485] : 
                       (N37)? mem_q[652] : 
                       (N32)? mem_q[819] : 
                       (N34)? mem_q[986] : 
                       (N36)? mem_q[1153] : 
                       (N38)? mem_q[1320] : 1'b0;
  assign data_o[150] = (N31)? mem_q[150] : 
                       (N33)? mem_q[317] : 
                       (N35)? mem_q[484] : 
                       (N37)? mem_q[651] : 
                       (N32)? mem_q[818] : 
                       (N34)? mem_q[985] : 
                       (N36)? mem_q[1152] : 
                       (N38)? mem_q[1319] : 1'b0;
  assign data_o[149] = (N31)? mem_q[149] : 
                       (N33)? mem_q[316] : 
                       (N35)? mem_q[483] : 
                       (N37)? mem_q[650] : 
                       (N32)? mem_q[817] : 
                       (N34)? mem_q[984] : 
                       (N36)? mem_q[1151] : 
                       (N38)? mem_q[1318] : 1'b0;
  assign data_o[148] = (N31)? mem_q[148] : 
                       (N33)? mem_q[315] : 
                       (N35)? mem_q[482] : 
                       (N37)? mem_q[649] : 
                       (N32)? mem_q[816] : 
                       (N34)? mem_q[983] : 
                       (N36)? mem_q[1150] : 
                       (N38)? mem_q[1317] : 1'b0;
  assign data_o[147] = (N31)? mem_q[147] : 
                       (N33)? mem_q[314] : 
                       (N35)? mem_q[481] : 
                       (N37)? mem_q[648] : 
                       (N32)? mem_q[815] : 
                       (N34)? mem_q[982] : 
                       (N36)? mem_q[1149] : 
                       (N38)? mem_q[1316] : 1'b0;
  assign data_o[146] = (N31)? mem_q[146] : 
                       (N33)? mem_q[313] : 
                       (N35)? mem_q[480] : 
                       (N37)? mem_q[647] : 
                       (N32)? mem_q[814] : 
                       (N34)? mem_q[981] : 
                       (N36)? mem_q[1148] : 
                       (N38)? mem_q[1315] : 1'b0;
  assign data_o[145] = (N31)? mem_q[145] : 
                       (N33)? mem_q[312] : 
                       (N35)? mem_q[479] : 
                       (N37)? mem_q[646] : 
                       (N32)? mem_q[813] : 
                       (N34)? mem_q[980] : 
                       (N36)? mem_q[1147] : 
                       (N38)? mem_q[1314] : 1'b0;
  assign data_o[144] = (N31)? mem_q[144] : 
                       (N33)? mem_q[311] : 
                       (N35)? mem_q[478] : 
                       (N37)? mem_q[645] : 
                       (N32)? mem_q[812] : 
                       (N34)? mem_q[979] : 
                       (N36)? mem_q[1146] : 
                       (N38)? mem_q[1313] : 1'b0;
  assign data_o[143] = (N31)? mem_q[143] : 
                       (N33)? mem_q[310] : 
                       (N35)? mem_q[477] : 
                       (N37)? mem_q[644] : 
                       (N32)? mem_q[811] : 
                       (N34)? mem_q[978] : 
                       (N36)? mem_q[1145] : 
                       (N38)? mem_q[1312] : 1'b0;
  assign data_o[142] = (N31)? mem_q[142] : 
                       (N33)? mem_q[309] : 
                       (N35)? mem_q[476] : 
                       (N37)? mem_q[643] : 
                       (N32)? mem_q[810] : 
                       (N34)? mem_q[977] : 
                       (N36)? mem_q[1144] : 
                       (N38)? mem_q[1311] : 1'b0;
  assign data_o[141] = (N31)? mem_q[141] : 
                       (N33)? mem_q[308] : 
                       (N35)? mem_q[475] : 
                       (N37)? mem_q[642] : 
                       (N32)? mem_q[809] : 
                       (N34)? mem_q[976] : 
                       (N36)? mem_q[1143] : 
                       (N38)? mem_q[1310] : 1'b0;
  assign data_o[140] = (N31)? mem_q[140] : 
                       (N33)? mem_q[307] : 
                       (N35)? mem_q[474] : 
                       (N37)? mem_q[641] : 
                       (N32)? mem_q[808] : 
                       (N34)? mem_q[975] : 
                       (N36)? mem_q[1142] : 
                       (N38)? mem_q[1309] : 1'b0;
  assign data_o[139] = (N31)? mem_q[139] : 
                       (N33)? mem_q[306] : 
                       (N35)? mem_q[473] : 
                       (N37)? mem_q[640] : 
                       (N32)? mem_q[807] : 
                       (N34)? mem_q[974] : 
                       (N36)? mem_q[1141] : 
                       (N38)? mem_q[1308] : 1'b0;
  assign data_o[138] = (N31)? mem_q[138] : 
                       (N33)? mem_q[305] : 
                       (N35)? mem_q[472] : 
                       (N37)? mem_q[639] : 
                       (N32)? mem_q[806] : 
                       (N34)? mem_q[973] : 
                       (N36)? mem_q[1140] : 
                       (N38)? mem_q[1307] : 1'b0;
  assign data_o[137] = (N31)? mem_q[137] : 
                       (N33)? mem_q[304] : 
                       (N35)? mem_q[471] : 
                       (N37)? mem_q[638] : 
                       (N32)? mem_q[805] : 
                       (N34)? mem_q[972] : 
                       (N36)? mem_q[1139] : 
                       (N38)? mem_q[1306] : 1'b0;
  assign data_o[136] = (N31)? mem_q[136] : 
                       (N33)? mem_q[303] : 
                       (N35)? mem_q[470] : 
                       (N37)? mem_q[637] : 
                       (N32)? mem_q[804] : 
                       (N34)? mem_q[971] : 
                       (N36)? mem_q[1138] : 
                       (N38)? mem_q[1305] : 1'b0;
  assign data_o[135] = (N31)? mem_q[135] : 
                       (N33)? mem_q[302] : 
                       (N35)? mem_q[469] : 
                       (N37)? mem_q[636] : 
                       (N32)? mem_q[803] : 
                       (N34)? mem_q[970] : 
                       (N36)? mem_q[1137] : 
                       (N38)? mem_q[1304] : 1'b0;
  assign data_o[134] = (N31)? mem_q[134] : 
                       (N33)? mem_q[301] : 
                       (N35)? mem_q[468] : 
                       (N37)? mem_q[635] : 
                       (N32)? mem_q[802] : 
                       (N34)? mem_q[969] : 
                       (N36)? mem_q[1136] : 
                       (N38)? mem_q[1303] : 1'b0;
  assign data_o[133] = (N31)? mem_q[133] : 
                       (N33)? mem_q[300] : 
                       (N35)? mem_q[467] : 
                       (N37)? mem_q[634] : 
                       (N32)? mem_q[801] : 
                       (N34)? mem_q[968] : 
                       (N36)? mem_q[1135] : 
                       (N38)? mem_q[1302] : 1'b0;
  assign data_o[132] = (N31)? mem_q[132] : 
                       (N33)? mem_q[299] : 
                       (N35)? mem_q[466] : 
                       (N37)? mem_q[633] : 
                       (N32)? mem_q[800] : 
                       (N34)? mem_q[967] : 
                       (N36)? mem_q[1134] : 
                       (N38)? mem_q[1301] : 1'b0;
  assign data_o[131] = (N31)? mem_q[131] : 
                       (N33)? mem_q[298] : 
                       (N35)? mem_q[465] : 
                       (N37)? mem_q[632] : 
                       (N32)? mem_q[799] : 
                       (N34)? mem_q[966] : 
                       (N36)? mem_q[1133] : 
                       (N38)? mem_q[1300] : 1'b0;
  assign data_o[130] = (N31)? mem_q[130] : 
                       (N33)? mem_q[297] : 
                       (N35)? mem_q[464] : 
                       (N37)? mem_q[631] : 
                       (N32)? mem_q[798] : 
                       (N34)? mem_q[965] : 
                       (N36)? mem_q[1132] : 
                       (N38)? mem_q[1299] : 1'b0;
  assign data_o[129] = (N31)? mem_q[129] : 
                       (N33)? mem_q[296] : 
                       (N35)? mem_q[463] : 
                       (N37)? mem_q[630] : 
                       (N32)? mem_q[797] : 
                       (N34)? mem_q[964] : 
                       (N36)? mem_q[1131] : 
                       (N38)? mem_q[1298] : 1'b0;
  assign data_o[128] = (N31)? mem_q[128] : 
                       (N33)? mem_q[295] : 
                       (N35)? mem_q[462] : 
                       (N37)? mem_q[629] : 
                       (N32)? mem_q[796] : 
                       (N34)? mem_q[963] : 
                       (N36)? mem_q[1130] : 
                       (N38)? mem_q[1297] : 1'b0;
  assign data_o[127] = (N31)? mem_q[127] : 
                       (N33)? mem_q[294] : 
                       (N35)? mem_q[461] : 
                       (N37)? mem_q[628] : 
                       (N32)? mem_q[795] : 
                       (N34)? mem_q[962] : 
                       (N36)? mem_q[1129] : 
                       (N38)? mem_q[1296] : 1'b0;
  assign data_o[126] = (N31)? mem_q[126] : 
                       (N33)? mem_q[293] : 
                       (N35)? mem_q[460] : 
                       (N37)? mem_q[627] : 
                       (N32)? mem_q[794] : 
                       (N34)? mem_q[961] : 
                       (N36)? mem_q[1128] : 
                       (N38)? mem_q[1295] : 1'b0;
  assign data_o[125] = (N31)? mem_q[125] : 
                       (N33)? mem_q[292] : 
                       (N35)? mem_q[459] : 
                       (N37)? mem_q[626] : 
                       (N32)? mem_q[793] : 
                       (N34)? mem_q[960] : 
                       (N36)? mem_q[1127] : 
                       (N38)? mem_q[1294] : 1'b0;
  assign data_o[124] = (N31)? mem_q[124] : 
                       (N33)? mem_q[291] : 
                       (N35)? mem_q[458] : 
                       (N37)? mem_q[625] : 
                       (N32)? mem_q[792] : 
                       (N34)? mem_q[959] : 
                       (N36)? mem_q[1126] : 
                       (N38)? mem_q[1293] : 1'b0;
  assign data_o[123] = (N31)? mem_q[123] : 
                       (N33)? mem_q[290] : 
                       (N35)? mem_q[457] : 
                       (N37)? mem_q[624] : 
                       (N32)? mem_q[791] : 
                       (N34)? mem_q[958] : 
                       (N36)? mem_q[1125] : 
                       (N38)? mem_q[1292] : 1'b0;
  assign data_o[122] = (N31)? mem_q[122] : 
                       (N33)? mem_q[289] : 
                       (N35)? mem_q[456] : 
                       (N37)? mem_q[623] : 
                       (N32)? mem_q[790] : 
                       (N34)? mem_q[957] : 
                       (N36)? mem_q[1124] : 
                       (N38)? mem_q[1291] : 1'b0;
  assign data_o[121] = (N31)? mem_q[121] : 
                       (N33)? mem_q[288] : 
                       (N35)? mem_q[455] : 
                       (N37)? mem_q[622] : 
                       (N32)? mem_q[789] : 
                       (N34)? mem_q[956] : 
                       (N36)? mem_q[1123] : 
                       (N38)? mem_q[1290] : 1'b0;
  assign data_o[120] = (N31)? mem_q[120] : 
                       (N33)? mem_q[287] : 
                       (N35)? mem_q[454] : 
                       (N37)? mem_q[621] : 
                       (N32)? mem_q[788] : 
                       (N34)? mem_q[955] : 
                       (N36)? mem_q[1122] : 
                       (N38)? mem_q[1289] : 1'b0;
  assign data_o[119] = (N31)? mem_q[119] : 
                       (N33)? mem_q[286] : 
                       (N35)? mem_q[453] : 
                       (N37)? mem_q[620] : 
                       (N32)? mem_q[787] : 
                       (N34)? mem_q[954] : 
                       (N36)? mem_q[1121] : 
                       (N38)? mem_q[1288] : 1'b0;
  assign data_o[118] = (N31)? mem_q[118] : 
                       (N33)? mem_q[285] : 
                       (N35)? mem_q[452] : 
                       (N37)? mem_q[619] : 
                       (N32)? mem_q[786] : 
                       (N34)? mem_q[953] : 
                       (N36)? mem_q[1120] : 
                       (N38)? mem_q[1287] : 1'b0;
  assign data_o[117] = (N31)? mem_q[117] : 
                       (N33)? mem_q[284] : 
                       (N35)? mem_q[451] : 
                       (N37)? mem_q[618] : 
                       (N32)? mem_q[785] : 
                       (N34)? mem_q[952] : 
                       (N36)? mem_q[1119] : 
                       (N38)? mem_q[1286] : 1'b0;
  assign data_o[116] = (N31)? mem_q[116] : 
                       (N33)? mem_q[283] : 
                       (N35)? mem_q[450] : 
                       (N37)? mem_q[617] : 
                       (N32)? mem_q[784] : 
                       (N34)? mem_q[951] : 
                       (N36)? mem_q[1118] : 
                       (N38)? mem_q[1285] : 1'b0;
  assign data_o[115] = (N31)? mem_q[115] : 
                       (N33)? mem_q[282] : 
                       (N35)? mem_q[449] : 
                       (N37)? mem_q[616] : 
                       (N32)? mem_q[783] : 
                       (N34)? mem_q[950] : 
                       (N36)? mem_q[1117] : 
                       (N38)? mem_q[1284] : 1'b0;
  assign data_o[114] = (N31)? mem_q[114] : 
                       (N33)? mem_q[281] : 
                       (N35)? mem_q[448] : 
                       (N37)? mem_q[615] : 
                       (N32)? mem_q[782] : 
                       (N34)? mem_q[949] : 
                       (N36)? mem_q[1116] : 
                       (N38)? mem_q[1283] : 1'b0;
  assign data_o[113] = (N31)? mem_q[113] : 
                       (N33)? mem_q[280] : 
                       (N35)? mem_q[447] : 
                       (N37)? mem_q[614] : 
                       (N32)? mem_q[781] : 
                       (N34)? mem_q[948] : 
                       (N36)? mem_q[1115] : 
                       (N38)? mem_q[1282] : 1'b0;
  assign data_o[112] = (N31)? mem_q[112] : 
                       (N33)? mem_q[279] : 
                       (N35)? mem_q[446] : 
                       (N37)? mem_q[613] : 
                       (N32)? mem_q[780] : 
                       (N34)? mem_q[947] : 
                       (N36)? mem_q[1114] : 
                       (N38)? mem_q[1281] : 1'b0;
  assign data_o[111] = (N31)? mem_q[111] : 
                       (N33)? mem_q[278] : 
                       (N35)? mem_q[445] : 
                       (N37)? mem_q[612] : 
                       (N32)? mem_q[779] : 
                       (N34)? mem_q[946] : 
                       (N36)? mem_q[1113] : 
                       (N38)? mem_q[1280] : 1'b0;
  assign data_o[110] = (N31)? mem_q[110] : 
                       (N33)? mem_q[277] : 
                       (N35)? mem_q[444] : 
                       (N37)? mem_q[611] : 
                       (N32)? mem_q[778] : 
                       (N34)? mem_q[945] : 
                       (N36)? mem_q[1112] : 
                       (N38)? mem_q[1279] : 1'b0;
  assign data_o[109] = (N31)? mem_q[109] : 
                       (N33)? mem_q[276] : 
                       (N35)? mem_q[443] : 
                       (N37)? mem_q[610] : 
                       (N32)? mem_q[777] : 
                       (N34)? mem_q[944] : 
                       (N36)? mem_q[1111] : 
                       (N38)? mem_q[1278] : 1'b0;
  assign data_o[108] = (N31)? mem_q[108] : 
                       (N33)? mem_q[275] : 
                       (N35)? mem_q[442] : 
                       (N37)? mem_q[609] : 
                       (N32)? mem_q[776] : 
                       (N34)? mem_q[943] : 
                       (N36)? mem_q[1110] : 
                       (N38)? mem_q[1277] : 1'b0;
  assign data_o[107] = (N31)? mem_q[107] : 
                       (N33)? mem_q[274] : 
                       (N35)? mem_q[441] : 
                       (N37)? mem_q[608] : 
                       (N32)? mem_q[775] : 
                       (N34)? mem_q[942] : 
                       (N36)? mem_q[1109] : 
                       (N38)? mem_q[1276] : 1'b0;
  assign data_o[106] = (N31)? mem_q[106] : 
                       (N33)? mem_q[273] : 
                       (N35)? mem_q[440] : 
                       (N37)? mem_q[607] : 
                       (N32)? mem_q[774] : 
                       (N34)? mem_q[941] : 
                       (N36)? mem_q[1108] : 
                       (N38)? mem_q[1275] : 1'b0;
  assign data_o[105] = (N31)? mem_q[105] : 
                       (N33)? mem_q[272] : 
                       (N35)? mem_q[439] : 
                       (N37)? mem_q[606] : 
                       (N32)? mem_q[773] : 
                       (N34)? mem_q[940] : 
                       (N36)? mem_q[1107] : 
                       (N38)? mem_q[1274] : 1'b0;
  assign data_o[104] = (N31)? mem_q[104] : 
                       (N33)? mem_q[271] : 
                       (N35)? mem_q[438] : 
                       (N37)? mem_q[605] : 
                       (N32)? mem_q[772] : 
                       (N34)? mem_q[939] : 
                       (N36)? mem_q[1106] : 
                       (N38)? mem_q[1273] : 1'b0;
  assign data_o[103] = (N31)? mem_q[103] : 
                       (N33)? mem_q[270] : 
                       (N35)? mem_q[437] : 
                       (N37)? mem_q[604] : 
                       (N32)? mem_q[771] : 
                       (N34)? mem_q[938] : 
                       (N36)? mem_q[1105] : 
                       (N38)? mem_q[1272] : 1'b0;
  assign data_o[102] = (N31)? mem_q[102] : 
                       (N33)? mem_q[269] : 
                       (N35)? mem_q[436] : 
                       (N37)? mem_q[603] : 
                       (N32)? mem_q[770] : 
                       (N34)? mem_q[937] : 
                       (N36)? mem_q[1104] : 
                       (N38)? mem_q[1271] : 1'b0;
  assign data_o[101] = (N31)? mem_q[101] : 
                       (N33)? mem_q[268] : 
                       (N35)? mem_q[435] : 
                       (N37)? mem_q[602] : 
                       (N32)? mem_q[769] : 
                       (N34)? mem_q[936] : 
                       (N36)? mem_q[1103] : 
                       (N38)? mem_q[1270] : 1'b0;
  assign data_o[100] = (N31)? mem_q[100] : 
                       (N33)? mem_q[267] : 
                       (N35)? mem_q[434] : 
                       (N37)? mem_q[601] : 
                       (N32)? mem_q[768] : 
                       (N34)? mem_q[935] : 
                       (N36)? mem_q[1102] : 
                       (N38)? mem_q[1269] : 1'b0;
  assign data_o[99] = (N31)? mem_q[99] : 
                      (N33)? mem_q[266] : 
                      (N35)? mem_q[433] : 
                      (N37)? mem_q[600] : 
                      (N32)? mem_q[767] : 
                      (N34)? mem_q[934] : 
                      (N36)? mem_q[1101] : 
                      (N38)? mem_q[1268] : 1'b0;
  assign data_o[98] = (N31)? mem_q[98] : 
                      (N33)? mem_q[265] : 
                      (N35)? mem_q[432] : 
                      (N37)? mem_q[599] : 
                      (N32)? mem_q[766] : 
                      (N34)? mem_q[933] : 
                      (N36)? mem_q[1100] : 
                      (N38)? mem_q[1267] : 1'b0;
  assign data_o[97] = (N31)? mem_q[97] : 
                      (N33)? mem_q[264] : 
                      (N35)? mem_q[431] : 
                      (N37)? mem_q[598] : 
                      (N32)? mem_q[765] : 
                      (N34)? mem_q[932] : 
                      (N36)? mem_q[1099] : 
                      (N38)? mem_q[1266] : 1'b0;
  assign data_o[96] = (N31)? mem_q[96] : 
                      (N33)? mem_q[263] : 
                      (N35)? mem_q[430] : 
                      (N37)? mem_q[597] : 
                      (N32)? mem_q[764] : 
                      (N34)? mem_q[931] : 
                      (N36)? mem_q[1098] : 
                      (N38)? mem_q[1265] : 1'b0;
  assign data_o[95] = (N31)? mem_q[95] : 
                      (N33)? mem_q[262] : 
                      (N35)? mem_q[429] : 
                      (N37)? mem_q[596] : 
                      (N32)? mem_q[763] : 
                      (N34)? mem_q[930] : 
                      (N36)? mem_q[1097] : 
                      (N38)? mem_q[1264] : 1'b0;
  assign data_o[94] = (N31)? mem_q[94] : 
                      (N33)? mem_q[261] : 
                      (N35)? mem_q[428] : 
                      (N37)? mem_q[595] : 
                      (N32)? mem_q[762] : 
                      (N34)? mem_q[929] : 
                      (N36)? mem_q[1096] : 
                      (N38)? mem_q[1263] : 1'b0;
  assign data_o[93] = (N31)? mem_q[93] : 
                      (N33)? mem_q[260] : 
                      (N35)? mem_q[427] : 
                      (N37)? mem_q[594] : 
                      (N32)? mem_q[761] : 
                      (N34)? mem_q[928] : 
                      (N36)? mem_q[1095] : 
                      (N38)? mem_q[1262] : 1'b0;
  assign data_o[92] = (N31)? mem_q[92] : 
                      (N33)? mem_q[259] : 
                      (N35)? mem_q[426] : 
                      (N37)? mem_q[593] : 
                      (N32)? mem_q[760] : 
                      (N34)? mem_q[927] : 
                      (N36)? mem_q[1094] : 
                      (N38)? mem_q[1261] : 1'b0;
  assign data_o[91] = (N31)? mem_q[91] : 
                      (N33)? mem_q[258] : 
                      (N35)? mem_q[425] : 
                      (N37)? mem_q[592] : 
                      (N32)? mem_q[759] : 
                      (N34)? mem_q[926] : 
                      (N36)? mem_q[1093] : 
                      (N38)? mem_q[1260] : 1'b0;
  assign data_o[90] = (N31)? mem_q[90] : 
                      (N33)? mem_q[257] : 
                      (N35)? mem_q[424] : 
                      (N37)? mem_q[591] : 
                      (N32)? mem_q[758] : 
                      (N34)? mem_q[925] : 
                      (N36)? mem_q[1092] : 
                      (N38)? mem_q[1259] : 1'b0;
  assign data_o[89] = (N31)? mem_q[89] : 
                      (N33)? mem_q[256] : 
                      (N35)? mem_q[423] : 
                      (N37)? mem_q[590] : 
                      (N32)? mem_q[757] : 
                      (N34)? mem_q[924] : 
                      (N36)? mem_q[1091] : 
                      (N38)? mem_q[1258] : 1'b0;
  assign data_o[88] = (N31)? mem_q[88] : 
                      (N33)? mem_q[255] : 
                      (N35)? mem_q[422] : 
                      (N37)? mem_q[589] : 
                      (N32)? mem_q[756] : 
                      (N34)? mem_q[923] : 
                      (N36)? mem_q[1090] : 
                      (N38)? mem_q[1257] : 1'b0;
  assign data_o[87] = (N31)? mem_q[87] : 
                      (N33)? mem_q[254] : 
                      (N35)? mem_q[421] : 
                      (N37)? mem_q[588] : 
                      (N32)? mem_q[755] : 
                      (N34)? mem_q[922] : 
                      (N36)? mem_q[1089] : 
                      (N38)? mem_q[1256] : 1'b0;
  assign data_o[86] = (N31)? mem_q[86] : 
                      (N33)? mem_q[253] : 
                      (N35)? mem_q[420] : 
                      (N37)? mem_q[587] : 
                      (N32)? mem_q[754] : 
                      (N34)? mem_q[921] : 
                      (N36)? mem_q[1088] : 
                      (N38)? mem_q[1255] : 1'b0;
  assign data_o[85] = (N31)? mem_q[85] : 
                      (N33)? mem_q[252] : 
                      (N35)? mem_q[419] : 
                      (N37)? mem_q[586] : 
                      (N32)? mem_q[753] : 
                      (N34)? mem_q[920] : 
                      (N36)? mem_q[1087] : 
                      (N38)? mem_q[1254] : 1'b0;
  assign data_o[84] = (N31)? mem_q[84] : 
                      (N33)? mem_q[251] : 
                      (N35)? mem_q[418] : 
                      (N37)? mem_q[585] : 
                      (N32)? mem_q[752] : 
                      (N34)? mem_q[919] : 
                      (N36)? mem_q[1086] : 
                      (N38)? mem_q[1253] : 1'b0;
  assign data_o[83] = (N31)? mem_q[83] : 
                      (N33)? mem_q[250] : 
                      (N35)? mem_q[417] : 
                      (N37)? mem_q[584] : 
                      (N32)? mem_q[751] : 
                      (N34)? mem_q[918] : 
                      (N36)? mem_q[1085] : 
                      (N38)? mem_q[1252] : 1'b0;
  assign data_o[82] = (N31)? mem_q[82] : 
                      (N33)? mem_q[249] : 
                      (N35)? mem_q[416] : 
                      (N37)? mem_q[583] : 
                      (N32)? mem_q[750] : 
                      (N34)? mem_q[917] : 
                      (N36)? mem_q[1084] : 
                      (N38)? mem_q[1251] : 1'b0;
  assign data_o[81] = (N31)? mem_q[81] : 
                      (N33)? mem_q[248] : 
                      (N35)? mem_q[415] : 
                      (N37)? mem_q[582] : 
                      (N32)? mem_q[749] : 
                      (N34)? mem_q[916] : 
                      (N36)? mem_q[1083] : 
                      (N38)? mem_q[1250] : 1'b0;
  assign data_o[80] = (N31)? mem_q[80] : 
                      (N33)? mem_q[247] : 
                      (N35)? mem_q[414] : 
                      (N37)? mem_q[581] : 
                      (N32)? mem_q[748] : 
                      (N34)? mem_q[915] : 
                      (N36)? mem_q[1082] : 
                      (N38)? mem_q[1249] : 1'b0;
  assign data_o[79] = (N31)? mem_q[79] : 
                      (N33)? mem_q[246] : 
                      (N35)? mem_q[413] : 
                      (N37)? mem_q[580] : 
                      (N32)? mem_q[747] : 
                      (N34)? mem_q[914] : 
                      (N36)? mem_q[1081] : 
                      (N38)? mem_q[1248] : 1'b0;
  assign data_o[78] = (N31)? mem_q[78] : 
                      (N33)? mem_q[245] : 
                      (N35)? mem_q[412] : 
                      (N37)? mem_q[579] : 
                      (N32)? mem_q[746] : 
                      (N34)? mem_q[913] : 
                      (N36)? mem_q[1080] : 
                      (N38)? mem_q[1247] : 1'b0;
  assign data_o[77] = (N31)? mem_q[77] : 
                      (N33)? mem_q[244] : 
                      (N35)? mem_q[411] : 
                      (N37)? mem_q[578] : 
                      (N32)? mem_q[745] : 
                      (N34)? mem_q[912] : 
                      (N36)? mem_q[1079] : 
                      (N38)? mem_q[1246] : 1'b0;
  assign data_o[76] = (N31)? mem_q[76] : 
                      (N33)? mem_q[243] : 
                      (N35)? mem_q[410] : 
                      (N37)? mem_q[577] : 
                      (N32)? mem_q[744] : 
                      (N34)? mem_q[911] : 
                      (N36)? mem_q[1078] : 
                      (N38)? mem_q[1245] : 1'b0;
  assign data_o[75] = (N31)? mem_q[75] : 
                      (N33)? mem_q[242] : 
                      (N35)? mem_q[409] : 
                      (N37)? mem_q[576] : 
                      (N32)? mem_q[743] : 
                      (N34)? mem_q[910] : 
                      (N36)? mem_q[1077] : 
                      (N38)? mem_q[1244] : 1'b0;
  assign data_o[74] = (N31)? mem_q[74] : 
                      (N33)? mem_q[241] : 
                      (N35)? mem_q[408] : 
                      (N37)? mem_q[575] : 
                      (N32)? mem_q[742] : 
                      (N34)? mem_q[909] : 
                      (N36)? mem_q[1076] : 
                      (N38)? mem_q[1243] : 1'b0;
  assign data_o[73] = (N31)? mem_q[73] : 
                      (N33)? mem_q[240] : 
                      (N35)? mem_q[407] : 
                      (N37)? mem_q[574] : 
                      (N32)? mem_q[741] : 
                      (N34)? mem_q[908] : 
                      (N36)? mem_q[1075] : 
                      (N38)? mem_q[1242] : 1'b0;
  assign data_o[72] = (N31)? mem_q[72] : 
                      (N33)? mem_q[239] : 
                      (N35)? mem_q[406] : 
                      (N37)? mem_q[573] : 
                      (N32)? mem_q[740] : 
                      (N34)? mem_q[907] : 
                      (N36)? mem_q[1074] : 
                      (N38)? mem_q[1241] : 1'b0;
  assign data_o[71] = (N31)? mem_q[71] : 
                      (N33)? mem_q[238] : 
                      (N35)? mem_q[405] : 
                      (N37)? mem_q[572] : 
                      (N32)? mem_q[739] : 
                      (N34)? mem_q[906] : 
                      (N36)? mem_q[1073] : 
                      (N38)? mem_q[1240] : 1'b0;
  assign data_o[70] = (N31)? mem_q[70] : 
                      (N33)? mem_q[237] : 
                      (N35)? mem_q[404] : 
                      (N37)? mem_q[571] : 
                      (N32)? mem_q[738] : 
                      (N34)? mem_q[905] : 
                      (N36)? mem_q[1072] : 
                      (N38)? mem_q[1239] : 1'b0;
  assign data_o[69] = (N31)? mem_q[69] : 
                      (N33)? mem_q[236] : 
                      (N35)? mem_q[403] : 
                      (N37)? mem_q[570] : 
                      (N32)? mem_q[737] : 
                      (N34)? mem_q[904] : 
                      (N36)? mem_q[1071] : 
                      (N38)? mem_q[1238] : 1'b0;
  assign data_o[68] = (N31)? mem_q[68] : 
                      (N33)? mem_q[235] : 
                      (N35)? mem_q[402] : 
                      (N37)? mem_q[569] : 
                      (N32)? mem_q[736] : 
                      (N34)? mem_q[903] : 
                      (N36)? mem_q[1070] : 
                      (N38)? mem_q[1237] : 1'b0;
  assign data_o[67] = (N31)? mem_q[67] : 
                      (N33)? mem_q[234] : 
                      (N35)? mem_q[401] : 
                      (N37)? mem_q[568] : 
                      (N32)? mem_q[735] : 
                      (N34)? mem_q[902] : 
                      (N36)? mem_q[1069] : 
                      (N38)? mem_q[1236] : 1'b0;
  assign data_o[66] = (N31)? mem_q[66] : 
                      (N33)? mem_q[233] : 
                      (N35)? mem_q[400] : 
                      (N37)? mem_q[567] : 
                      (N32)? mem_q[734] : 
                      (N34)? mem_q[901] : 
                      (N36)? mem_q[1068] : 
                      (N38)? mem_q[1235] : 1'b0;
  assign data_o[65] = (N31)? mem_q[65] : 
                      (N33)? mem_q[232] : 
                      (N35)? mem_q[399] : 
                      (N37)? mem_q[566] : 
                      (N32)? mem_q[733] : 
                      (N34)? mem_q[900] : 
                      (N36)? mem_q[1067] : 
                      (N38)? mem_q[1234] : 1'b0;
  assign data_o[64] = (N31)? mem_q[64] : 
                      (N33)? mem_q[231] : 
                      (N35)? mem_q[398] : 
                      (N37)? mem_q[565] : 
                      (N32)? mem_q[732] : 
                      (N34)? mem_q[899] : 
                      (N36)? mem_q[1066] : 
                      (N38)? mem_q[1233] : 1'b0;
  assign data_o[63] = (N31)? mem_q[63] : 
                      (N33)? mem_q[230] : 
                      (N35)? mem_q[397] : 
                      (N37)? mem_q[564] : 
                      (N32)? mem_q[731] : 
                      (N34)? mem_q[898] : 
                      (N36)? mem_q[1065] : 
                      (N38)? mem_q[1232] : 1'b0;
  assign data_o[62] = (N31)? mem_q[62] : 
                      (N33)? mem_q[229] : 
                      (N35)? mem_q[396] : 
                      (N37)? mem_q[563] : 
                      (N32)? mem_q[730] : 
                      (N34)? mem_q[897] : 
                      (N36)? mem_q[1064] : 
                      (N38)? mem_q[1231] : 1'b0;
  assign data_o[61] = (N31)? mem_q[61] : 
                      (N33)? mem_q[228] : 
                      (N35)? mem_q[395] : 
                      (N37)? mem_q[562] : 
                      (N32)? mem_q[729] : 
                      (N34)? mem_q[896] : 
                      (N36)? mem_q[1063] : 
                      (N38)? mem_q[1230] : 1'b0;
  assign data_o[60] = (N31)? mem_q[60] : 
                      (N33)? mem_q[227] : 
                      (N35)? mem_q[394] : 
                      (N37)? mem_q[561] : 
                      (N32)? mem_q[728] : 
                      (N34)? mem_q[895] : 
                      (N36)? mem_q[1062] : 
                      (N38)? mem_q[1229] : 1'b0;
  assign data_o[59] = (N31)? mem_q[59] : 
                      (N33)? mem_q[226] : 
                      (N35)? mem_q[393] : 
                      (N37)? mem_q[560] : 
                      (N32)? mem_q[727] : 
                      (N34)? mem_q[894] : 
                      (N36)? mem_q[1061] : 
                      (N38)? mem_q[1228] : 1'b0;
  assign data_o[58] = (N31)? mem_q[58] : 
                      (N33)? mem_q[225] : 
                      (N35)? mem_q[392] : 
                      (N37)? mem_q[559] : 
                      (N32)? mem_q[726] : 
                      (N34)? mem_q[893] : 
                      (N36)? mem_q[1060] : 
                      (N38)? mem_q[1227] : 1'b0;
  assign data_o[57] = (N31)? mem_q[57] : 
                      (N33)? mem_q[224] : 
                      (N35)? mem_q[391] : 
                      (N37)? mem_q[558] : 
                      (N32)? mem_q[725] : 
                      (N34)? mem_q[892] : 
                      (N36)? mem_q[1059] : 
                      (N38)? mem_q[1226] : 1'b0;
  assign data_o[56] = (N31)? mem_q[56] : 
                      (N33)? mem_q[223] : 
                      (N35)? mem_q[390] : 
                      (N37)? mem_q[557] : 
                      (N32)? mem_q[724] : 
                      (N34)? mem_q[891] : 
                      (N36)? mem_q[1058] : 
                      (N38)? mem_q[1225] : 1'b0;
  assign data_o[55] = (N31)? mem_q[55] : 
                      (N33)? mem_q[222] : 
                      (N35)? mem_q[389] : 
                      (N37)? mem_q[556] : 
                      (N32)? mem_q[723] : 
                      (N34)? mem_q[890] : 
                      (N36)? mem_q[1057] : 
                      (N38)? mem_q[1224] : 1'b0;
  assign data_o[54] = (N31)? mem_q[54] : 
                      (N33)? mem_q[221] : 
                      (N35)? mem_q[388] : 
                      (N37)? mem_q[555] : 
                      (N32)? mem_q[722] : 
                      (N34)? mem_q[889] : 
                      (N36)? mem_q[1056] : 
                      (N38)? mem_q[1223] : 1'b0;
  assign data_o[53] = (N31)? mem_q[53] : 
                      (N33)? mem_q[220] : 
                      (N35)? mem_q[387] : 
                      (N37)? mem_q[554] : 
                      (N32)? mem_q[721] : 
                      (N34)? mem_q[888] : 
                      (N36)? mem_q[1055] : 
                      (N38)? mem_q[1222] : 1'b0;
  assign data_o[52] = (N31)? mem_q[52] : 
                      (N33)? mem_q[219] : 
                      (N35)? mem_q[386] : 
                      (N37)? mem_q[553] : 
                      (N32)? mem_q[720] : 
                      (N34)? mem_q[887] : 
                      (N36)? mem_q[1054] : 
                      (N38)? mem_q[1221] : 1'b0;
  assign data_o[51] = (N31)? mem_q[51] : 
                      (N33)? mem_q[218] : 
                      (N35)? mem_q[385] : 
                      (N37)? mem_q[552] : 
                      (N32)? mem_q[719] : 
                      (N34)? mem_q[886] : 
                      (N36)? mem_q[1053] : 
                      (N38)? mem_q[1220] : 1'b0;
  assign data_o[50] = (N31)? mem_q[50] : 
                      (N33)? mem_q[217] : 
                      (N35)? mem_q[384] : 
                      (N37)? mem_q[551] : 
                      (N32)? mem_q[718] : 
                      (N34)? mem_q[885] : 
                      (N36)? mem_q[1052] : 
                      (N38)? mem_q[1219] : 1'b0;
  assign data_o[49] = (N31)? mem_q[49] : 
                      (N33)? mem_q[216] : 
                      (N35)? mem_q[383] : 
                      (N37)? mem_q[550] : 
                      (N32)? mem_q[717] : 
                      (N34)? mem_q[884] : 
                      (N36)? mem_q[1051] : 
                      (N38)? mem_q[1218] : 1'b0;
  assign data_o[48] = (N31)? mem_q[48] : 
                      (N33)? mem_q[215] : 
                      (N35)? mem_q[382] : 
                      (N37)? mem_q[549] : 
                      (N32)? mem_q[716] : 
                      (N34)? mem_q[883] : 
                      (N36)? mem_q[1050] : 
                      (N38)? mem_q[1217] : 1'b0;
  assign data_o[47] = (N31)? mem_q[47] : 
                      (N33)? mem_q[214] : 
                      (N35)? mem_q[381] : 
                      (N37)? mem_q[548] : 
                      (N32)? mem_q[715] : 
                      (N34)? mem_q[882] : 
                      (N36)? mem_q[1049] : 
                      (N38)? mem_q[1216] : 1'b0;
  assign data_o[46] = (N31)? mem_q[46] : 
                      (N33)? mem_q[213] : 
                      (N35)? mem_q[380] : 
                      (N37)? mem_q[547] : 
                      (N32)? mem_q[714] : 
                      (N34)? mem_q[881] : 
                      (N36)? mem_q[1048] : 
                      (N38)? mem_q[1215] : 1'b0;
  assign data_o[45] = (N31)? mem_q[45] : 
                      (N33)? mem_q[212] : 
                      (N35)? mem_q[379] : 
                      (N37)? mem_q[546] : 
                      (N32)? mem_q[713] : 
                      (N34)? mem_q[880] : 
                      (N36)? mem_q[1047] : 
                      (N38)? mem_q[1214] : 1'b0;
  assign data_o[44] = (N31)? mem_q[44] : 
                      (N33)? mem_q[211] : 
                      (N35)? mem_q[378] : 
                      (N37)? mem_q[545] : 
                      (N32)? mem_q[712] : 
                      (N34)? mem_q[879] : 
                      (N36)? mem_q[1046] : 
                      (N38)? mem_q[1213] : 1'b0;
  assign data_o[43] = (N31)? mem_q[43] : 
                      (N33)? mem_q[210] : 
                      (N35)? mem_q[377] : 
                      (N37)? mem_q[544] : 
                      (N32)? mem_q[711] : 
                      (N34)? mem_q[878] : 
                      (N36)? mem_q[1045] : 
                      (N38)? mem_q[1212] : 1'b0;
  assign data_o[42] = (N31)? mem_q[42] : 
                      (N33)? mem_q[209] : 
                      (N35)? mem_q[376] : 
                      (N37)? mem_q[543] : 
                      (N32)? mem_q[710] : 
                      (N34)? mem_q[877] : 
                      (N36)? mem_q[1044] : 
                      (N38)? mem_q[1211] : 1'b0;
  assign data_o[41] = (N31)? mem_q[41] : 
                      (N33)? mem_q[208] : 
                      (N35)? mem_q[375] : 
                      (N37)? mem_q[542] : 
                      (N32)? mem_q[709] : 
                      (N34)? mem_q[876] : 
                      (N36)? mem_q[1043] : 
                      (N38)? mem_q[1210] : 1'b0;
  assign data_o[40] = (N31)? mem_q[40] : 
                      (N33)? mem_q[207] : 
                      (N35)? mem_q[374] : 
                      (N37)? mem_q[541] : 
                      (N32)? mem_q[708] : 
                      (N34)? mem_q[875] : 
                      (N36)? mem_q[1042] : 
                      (N38)? mem_q[1209] : 1'b0;
  assign data_o[39] = (N31)? mem_q[39] : 
                      (N33)? mem_q[206] : 
                      (N35)? mem_q[373] : 
                      (N37)? mem_q[540] : 
                      (N32)? mem_q[707] : 
                      (N34)? mem_q[874] : 
                      (N36)? mem_q[1041] : 
                      (N38)? mem_q[1208] : 1'b0;
  assign data_o[38] = (N31)? mem_q[38] : 
                      (N33)? mem_q[205] : 
                      (N35)? mem_q[372] : 
                      (N37)? mem_q[539] : 
                      (N32)? mem_q[706] : 
                      (N34)? mem_q[873] : 
                      (N36)? mem_q[1040] : 
                      (N38)? mem_q[1207] : 1'b0;
  assign data_o[37] = (N31)? mem_q[37] : 
                      (N33)? mem_q[204] : 
                      (N35)? mem_q[371] : 
                      (N37)? mem_q[538] : 
                      (N32)? mem_q[705] : 
                      (N34)? mem_q[872] : 
                      (N36)? mem_q[1039] : 
                      (N38)? mem_q[1206] : 1'b0;
  assign data_o[36] = (N31)? mem_q[36] : 
                      (N33)? mem_q[203] : 
                      (N35)? mem_q[370] : 
                      (N37)? mem_q[537] : 
                      (N32)? mem_q[704] : 
                      (N34)? mem_q[871] : 
                      (N36)? mem_q[1038] : 
                      (N38)? mem_q[1205] : 1'b0;
  assign data_o[35] = (N31)? mem_q[35] : 
                      (N33)? mem_q[202] : 
                      (N35)? mem_q[369] : 
                      (N37)? mem_q[536] : 
                      (N32)? mem_q[703] : 
                      (N34)? mem_q[870] : 
                      (N36)? mem_q[1037] : 
                      (N38)? mem_q[1204] : 1'b0;
  assign data_o[34] = (N31)? mem_q[34] : 
                      (N33)? mem_q[201] : 
                      (N35)? mem_q[368] : 
                      (N37)? mem_q[535] : 
                      (N32)? mem_q[702] : 
                      (N34)? mem_q[869] : 
                      (N36)? mem_q[1036] : 
                      (N38)? mem_q[1203] : 1'b0;
  assign data_o[33] = (N31)? mem_q[33] : 
                      (N33)? mem_q[200] : 
                      (N35)? mem_q[367] : 
                      (N37)? mem_q[534] : 
                      (N32)? mem_q[701] : 
                      (N34)? mem_q[868] : 
                      (N36)? mem_q[1035] : 
                      (N38)? mem_q[1202] : 1'b0;
  assign data_o[32] = (N31)? mem_q[32] : 
                      (N33)? mem_q[199] : 
                      (N35)? mem_q[366] : 
                      (N37)? mem_q[533] : 
                      (N32)? mem_q[700] : 
                      (N34)? mem_q[867] : 
                      (N36)? mem_q[1034] : 
                      (N38)? mem_q[1201] : 1'b0;
  assign data_o[31] = (N31)? mem_q[31] : 
                      (N33)? mem_q[198] : 
                      (N35)? mem_q[365] : 
                      (N37)? mem_q[532] : 
                      (N32)? mem_q[699] : 
                      (N34)? mem_q[866] : 
                      (N36)? mem_q[1033] : 
                      (N38)? mem_q[1200] : 1'b0;
  assign data_o[30] = (N31)? mem_q[30] : 
                      (N33)? mem_q[197] : 
                      (N35)? mem_q[364] : 
                      (N37)? mem_q[531] : 
                      (N32)? mem_q[698] : 
                      (N34)? mem_q[865] : 
                      (N36)? mem_q[1032] : 
                      (N38)? mem_q[1199] : 1'b0;
  assign data_o[29] = (N31)? mem_q[29] : 
                      (N33)? mem_q[196] : 
                      (N35)? mem_q[363] : 
                      (N37)? mem_q[530] : 
                      (N32)? mem_q[697] : 
                      (N34)? mem_q[864] : 
                      (N36)? mem_q[1031] : 
                      (N38)? mem_q[1198] : 1'b0;
  assign data_o[28] = (N31)? mem_q[28] : 
                      (N33)? mem_q[195] : 
                      (N35)? mem_q[362] : 
                      (N37)? mem_q[529] : 
                      (N32)? mem_q[696] : 
                      (N34)? mem_q[863] : 
                      (N36)? mem_q[1030] : 
                      (N38)? mem_q[1197] : 1'b0;
  assign data_o[27] = (N31)? mem_q[27] : 
                      (N33)? mem_q[194] : 
                      (N35)? mem_q[361] : 
                      (N37)? mem_q[528] : 
                      (N32)? mem_q[695] : 
                      (N34)? mem_q[862] : 
                      (N36)? mem_q[1029] : 
                      (N38)? mem_q[1196] : 1'b0;
  assign data_o[26] = (N31)? mem_q[26] : 
                      (N33)? mem_q[193] : 
                      (N35)? mem_q[360] : 
                      (N37)? mem_q[527] : 
                      (N32)? mem_q[694] : 
                      (N34)? mem_q[861] : 
                      (N36)? mem_q[1028] : 
                      (N38)? mem_q[1195] : 1'b0;
  assign data_o[25] = (N31)? mem_q[25] : 
                      (N33)? mem_q[192] : 
                      (N35)? mem_q[359] : 
                      (N37)? mem_q[526] : 
                      (N32)? mem_q[693] : 
                      (N34)? mem_q[860] : 
                      (N36)? mem_q[1027] : 
                      (N38)? mem_q[1194] : 1'b0;
  assign data_o[24] = (N31)? mem_q[24] : 
                      (N33)? mem_q[191] : 
                      (N35)? mem_q[358] : 
                      (N37)? mem_q[525] : 
                      (N32)? mem_q[692] : 
                      (N34)? mem_q[859] : 
                      (N36)? mem_q[1026] : 
                      (N38)? mem_q[1193] : 1'b0;
  assign data_o[23] = (N31)? mem_q[23] : 
                      (N33)? mem_q[190] : 
                      (N35)? mem_q[357] : 
                      (N37)? mem_q[524] : 
                      (N32)? mem_q[691] : 
                      (N34)? mem_q[858] : 
                      (N36)? mem_q[1025] : 
                      (N38)? mem_q[1192] : 1'b0;
  assign data_o[22] = (N31)? mem_q[22] : 
                      (N33)? mem_q[189] : 
                      (N35)? mem_q[356] : 
                      (N37)? mem_q[523] : 
                      (N32)? mem_q[690] : 
                      (N34)? mem_q[857] : 
                      (N36)? mem_q[1024] : 
                      (N38)? mem_q[1191] : 1'b0;
  assign data_o[21] = (N31)? mem_q[21] : 
                      (N33)? mem_q[188] : 
                      (N35)? mem_q[355] : 
                      (N37)? mem_q[522] : 
                      (N32)? mem_q[689] : 
                      (N34)? mem_q[856] : 
                      (N36)? mem_q[1023] : 
                      (N38)? mem_q[1190] : 1'b0;
  assign data_o[20] = (N31)? mem_q[20] : 
                      (N33)? mem_q[187] : 
                      (N35)? mem_q[354] : 
                      (N37)? mem_q[521] : 
                      (N32)? mem_q[688] : 
                      (N34)? mem_q[855] : 
                      (N36)? mem_q[1022] : 
                      (N38)? mem_q[1189] : 1'b0;
  assign data_o[19] = (N31)? mem_q[19] : 
                      (N33)? mem_q[186] : 
                      (N35)? mem_q[353] : 
                      (N37)? mem_q[520] : 
                      (N32)? mem_q[687] : 
                      (N34)? mem_q[854] : 
                      (N36)? mem_q[1021] : 
                      (N38)? mem_q[1188] : 1'b0;
  assign data_o[18] = (N31)? mem_q[18] : 
                      (N33)? mem_q[185] : 
                      (N35)? mem_q[352] : 
                      (N37)? mem_q[519] : 
                      (N32)? mem_q[686] : 
                      (N34)? mem_q[853] : 
                      (N36)? mem_q[1020] : 
                      (N38)? mem_q[1187] : 1'b0;
  assign data_o[17] = (N31)? mem_q[17] : 
                      (N33)? mem_q[184] : 
                      (N35)? mem_q[351] : 
                      (N37)? mem_q[518] : 
                      (N32)? mem_q[685] : 
                      (N34)? mem_q[852] : 
                      (N36)? mem_q[1019] : 
                      (N38)? mem_q[1186] : 1'b0;
  assign data_o[16] = (N31)? mem_q[16] : 
                      (N33)? mem_q[183] : 
                      (N35)? mem_q[350] : 
                      (N37)? mem_q[517] : 
                      (N32)? mem_q[684] : 
                      (N34)? mem_q[851] : 
                      (N36)? mem_q[1018] : 
                      (N38)? mem_q[1185] : 1'b0;
  assign data_o[15] = (N31)? mem_q[15] : 
                      (N33)? mem_q[182] : 
                      (N35)? mem_q[349] : 
                      (N37)? mem_q[516] : 
                      (N32)? mem_q[683] : 
                      (N34)? mem_q[850] : 
                      (N36)? mem_q[1017] : 
                      (N38)? mem_q[1184] : 1'b0;
  assign data_o[14] = (N31)? mem_q[14] : 
                      (N33)? mem_q[181] : 
                      (N35)? mem_q[348] : 
                      (N37)? mem_q[515] : 
                      (N32)? mem_q[682] : 
                      (N34)? mem_q[849] : 
                      (N36)? mem_q[1016] : 
                      (N38)? mem_q[1183] : 1'b0;
  assign data_o[13] = (N31)? mem_q[13] : 
                      (N33)? mem_q[180] : 
                      (N35)? mem_q[347] : 
                      (N37)? mem_q[514] : 
                      (N32)? mem_q[681] : 
                      (N34)? mem_q[848] : 
                      (N36)? mem_q[1015] : 
                      (N38)? mem_q[1182] : 1'b0;
  assign data_o[12] = (N31)? mem_q[12] : 
                      (N33)? mem_q[179] : 
                      (N35)? mem_q[346] : 
                      (N37)? mem_q[513] : 
                      (N32)? mem_q[680] : 
                      (N34)? mem_q[847] : 
                      (N36)? mem_q[1014] : 
                      (N38)? mem_q[1181] : 1'b0;
  assign data_o[11] = (N31)? mem_q[11] : 
                      (N33)? mem_q[178] : 
                      (N35)? mem_q[345] : 
                      (N37)? mem_q[512] : 
                      (N32)? mem_q[679] : 
                      (N34)? mem_q[846] : 
                      (N36)? mem_q[1013] : 
                      (N38)? mem_q[1180] : 1'b0;
  assign data_o[10] = (N31)? mem_q[10] : 
                      (N33)? mem_q[177] : 
                      (N35)? mem_q[344] : 
                      (N37)? mem_q[511] : 
                      (N32)? mem_q[678] : 
                      (N34)? mem_q[845] : 
                      (N36)? mem_q[1012] : 
                      (N38)? mem_q[1179] : 1'b0;
  assign data_o[9] = (N31)? mem_q[9] : 
                     (N33)? mem_q[176] : 
                     (N35)? mem_q[343] : 
                     (N37)? mem_q[510] : 
                     (N32)? mem_q[677] : 
                     (N34)? mem_q[844] : 
                     (N36)? mem_q[1011] : 
                     (N38)? mem_q[1178] : 1'b0;
  assign data_o[8] = (N31)? mem_q[8] : 
                     (N33)? mem_q[175] : 
                     (N35)? mem_q[342] : 
                     (N37)? mem_q[509] : 
                     (N32)? mem_q[676] : 
                     (N34)? mem_q[843] : 
                     (N36)? mem_q[1010] : 
                     (N38)? mem_q[1177] : 1'b0;
  assign data_o[7] = (N31)? mem_q[7] : 
                     (N33)? mem_q[174] : 
                     (N35)? mem_q[341] : 
                     (N37)? mem_q[508] : 
                     (N32)? mem_q[675] : 
                     (N34)? mem_q[842] : 
                     (N36)? mem_q[1009] : 
                     (N38)? mem_q[1176] : 1'b0;
  assign data_o[6] = (N31)? mem_q[6] : 
                     (N33)? mem_q[173] : 
                     (N35)? mem_q[340] : 
                     (N37)? mem_q[507] : 
                     (N32)? mem_q[674] : 
                     (N34)? mem_q[841] : 
                     (N36)? mem_q[1008] : 
                     (N38)? mem_q[1175] : 1'b0;
  assign data_o[5] = (N31)? mem_q[5] : 
                     (N33)? mem_q[172] : 
                     (N35)? mem_q[339] : 
                     (N37)? mem_q[506] : 
                     (N32)? mem_q[673] : 
                     (N34)? mem_q[840] : 
                     (N36)? mem_q[1007] : 
                     (N38)? mem_q[1174] : 1'b0;
  assign data_o[4] = (N31)? mem_q[4] : 
                     (N33)? mem_q[171] : 
                     (N35)? mem_q[338] : 
                     (N37)? mem_q[505] : 
                     (N32)? mem_q[672] : 
                     (N34)? mem_q[839] : 
                     (N36)? mem_q[1006] : 
                     (N38)? mem_q[1173] : 1'b0;
  assign data_o[3] = (N31)? mem_q[3] : 
                     (N33)? mem_q[170] : 
                     (N35)? mem_q[337] : 
                     (N37)? mem_q[504] : 
                     (N32)? mem_q[671] : 
                     (N34)? mem_q[838] : 
                     (N36)? mem_q[1005] : 
                     (N38)? mem_q[1172] : 1'b0;
  assign data_o[2] = (N31)? mem_q[2] : 
                     (N33)? mem_q[169] : 
                     (N35)? mem_q[336] : 
                     (N37)? mem_q[503] : 
                     (N32)? mem_q[670] : 
                     (N34)? mem_q[837] : 
                     (N36)? mem_q[1004] : 
                     (N38)? mem_q[1171] : 1'b0;
  assign data_o[1] = (N31)? mem_q[1] : 
                     (N33)? mem_q[168] : 
                     (N35)? mem_q[335] : 
                     (N37)? mem_q[502] : 
                     (N32)? mem_q[669] : 
                     (N34)? mem_q[836] : 
                     (N36)? mem_q[1003] : 
                     (N38)? mem_q[1170] : 1'b0;
  assign data_o[0] = (N31)? mem_q[0] : 
                     (N33)? mem_q[167] : 
                     (N35)? mem_q[334] : 
                     (N37)? mem_q[501] : 
                     (N32)? mem_q[668] : 
                     (N34)? mem_q[835] : 
                     (N36)? mem_q[1002] : 
                     (N38)? mem_q[1169] : 1'b0;

  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      status_cnt_q[3] <= 1'b0;
    end else if(N1433) begin
      status_cnt_q[3] <= N1426;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      usage_o[2] <= 1'b0;
    end else if(N1433) begin
      usage_o[2] <= N1425;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      usage_o[1] <= 1'b0;
    end else if(N1433) begin
      usage_o[1] <= N1424;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      usage_o[0] <= 1'b0;
    end else if(N1433) begin
      usage_o[0] <= N1423;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      read_pointer_q[2] <= 1'b0;
    end else if(N1435) begin
      read_pointer_q[2] <= N1419;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      read_pointer_q[1] <= 1'b0;
    end else if(N1435) begin
      read_pointer_q[1] <= N1418;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      read_pointer_q[0] <= 1'b0;
    end else if(N1435) begin
      read_pointer_q[0] <= N1417;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      write_pointer_q[2] <= 1'b0;
    end else if(N1437) begin
      write_pointer_q[2] <= N1422;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      write_pointer_q[1] <= 1'b0;
    end else if(N1437) begin
      write_pointer_q[1] <= N1421;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      write_pointer_q[0] <= 1'b0;
    end else if(N1437) begin
      write_pointer_q[0] <= N1420;
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1335] <= 1'b0;
    end else if(N1427) begin
      mem_q[1335] <= mem_n[1335];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1334] <= 1'b0;
    end else if(N1427) begin
      mem_q[1334] <= mem_n[1334];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1333] <= 1'b0;
    end else if(N1427) begin
      mem_q[1333] <= mem_n[1333];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1332] <= 1'b0;
    end else if(N1427) begin
      mem_q[1332] <= mem_n[1332];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1331] <= 1'b0;
    end else if(N1427) begin
      mem_q[1331] <= mem_n[1331];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1330] <= 1'b0;
    end else if(N1427) begin
      mem_q[1330] <= mem_n[1330];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1329] <= 1'b0;
    end else if(N1427) begin
      mem_q[1329] <= mem_n[1329];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1328] <= 1'b0;
    end else if(N1427) begin
      mem_q[1328] <= mem_n[1328];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1327] <= 1'b0;
    end else if(N1427) begin
      mem_q[1327] <= mem_n[1327];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1326] <= 1'b0;
    end else if(N1427) begin
      mem_q[1326] <= mem_n[1326];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1325] <= 1'b0;
    end else if(N1427) begin
      mem_q[1325] <= mem_n[1325];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1324] <= 1'b0;
    end else if(N1427) begin
      mem_q[1324] <= mem_n[1324];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1323] <= 1'b0;
    end else if(N1427) begin
      mem_q[1323] <= mem_n[1323];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1322] <= 1'b0;
    end else if(N1427) begin
      mem_q[1322] <= mem_n[1322];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1321] <= 1'b0;
    end else if(N1427) begin
      mem_q[1321] <= mem_n[1321];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1320] <= 1'b0;
    end else if(N1427) begin
      mem_q[1320] <= mem_n[1320];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1319] <= 1'b0;
    end else if(N1427) begin
      mem_q[1319] <= mem_n[1319];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1318] <= 1'b0;
    end else if(N1427) begin
      mem_q[1318] <= mem_n[1318];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1317] <= 1'b0;
    end else if(N1427) begin
      mem_q[1317] <= mem_n[1317];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1316] <= 1'b0;
    end else if(N1427) begin
      mem_q[1316] <= mem_n[1316];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1315] <= 1'b0;
    end else if(N1427) begin
      mem_q[1315] <= mem_n[1315];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1314] <= 1'b0;
    end else if(N1427) begin
      mem_q[1314] <= mem_n[1314];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1313] <= 1'b0;
    end else if(N1427) begin
      mem_q[1313] <= mem_n[1313];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1312] <= 1'b0;
    end else if(N1427) begin
      mem_q[1312] <= mem_n[1312];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1311] <= 1'b0;
    end else if(N1427) begin
      mem_q[1311] <= mem_n[1311];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1310] <= 1'b0;
    end else if(N1427) begin
      mem_q[1310] <= mem_n[1310];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1309] <= 1'b0;
    end else if(N1427) begin
      mem_q[1309] <= mem_n[1309];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1308] <= 1'b0;
    end else if(N1427) begin
      mem_q[1308] <= mem_n[1308];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1307] <= 1'b0;
    end else if(N1427) begin
      mem_q[1307] <= mem_n[1307];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1306] <= 1'b0;
    end else if(N1427) begin
      mem_q[1306] <= mem_n[1306];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1305] <= 1'b0;
    end else if(N1427) begin
      mem_q[1305] <= mem_n[1305];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1304] <= 1'b0;
    end else if(N1427) begin
      mem_q[1304] <= mem_n[1304];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1303] <= 1'b0;
    end else if(N1427) begin
      mem_q[1303] <= mem_n[1303];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1302] <= 1'b0;
    end else if(N1427) begin
      mem_q[1302] <= mem_n[1302];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1301] <= 1'b0;
    end else if(N1427) begin
      mem_q[1301] <= mem_n[1301];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1300] <= 1'b0;
    end else if(N1427) begin
      mem_q[1300] <= mem_n[1300];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1299] <= 1'b0;
    end else if(N1427) begin
      mem_q[1299] <= mem_n[1299];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1298] <= 1'b0;
    end else if(N1427) begin
      mem_q[1298] <= mem_n[1298];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1297] <= 1'b0;
    end else if(N1427) begin
      mem_q[1297] <= mem_n[1297];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1296] <= 1'b0;
    end else if(N1427) begin
      mem_q[1296] <= mem_n[1296];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1295] <= 1'b0;
    end else if(N1427) begin
      mem_q[1295] <= mem_n[1295];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1294] <= 1'b0;
    end else if(N1427) begin
      mem_q[1294] <= mem_n[1294];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1293] <= 1'b0;
    end else if(N1427) begin
      mem_q[1293] <= mem_n[1293];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1292] <= 1'b0;
    end else if(N1427) begin
      mem_q[1292] <= mem_n[1292];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1291] <= 1'b0;
    end else if(N1427) begin
      mem_q[1291] <= mem_n[1291];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1290] <= 1'b0;
    end else if(N1427) begin
      mem_q[1290] <= mem_n[1290];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1289] <= 1'b0;
    end else if(N1427) begin
      mem_q[1289] <= mem_n[1289];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1288] <= 1'b0;
    end else if(N1427) begin
      mem_q[1288] <= mem_n[1288];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1287] <= 1'b0;
    end else if(N1427) begin
      mem_q[1287] <= mem_n[1287];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1286] <= 1'b0;
    end else if(N1427) begin
      mem_q[1286] <= mem_n[1286];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1285] <= 1'b0;
    end else if(N1427) begin
      mem_q[1285] <= mem_n[1285];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1284] <= 1'b0;
    end else if(N1427) begin
      mem_q[1284] <= mem_n[1284];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1283] <= 1'b0;
    end else if(N1427) begin
      mem_q[1283] <= mem_n[1283];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1282] <= 1'b0;
    end else if(N1427) begin
      mem_q[1282] <= mem_n[1282];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1281] <= 1'b0;
    end else if(N1427) begin
      mem_q[1281] <= mem_n[1281];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1280] <= 1'b0;
    end else if(N1427) begin
      mem_q[1280] <= mem_n[1280];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1279] <= 1'b0;
    end else if(N1427) begin
      mem_q[1279] <= mem_n[1279];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1278] <= 1'b0;
    end else if(N1427) begin
      mem_q[1278] <= mem_n[1278];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1277] <= 1'b0;
    end else if(N1427) begin
      mem_q[1277] <= mem_n[1277];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1276] <= 1'b0;
    end else if(N1427) begin
      mem_q[1276] <= mem_n[1276];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1275] <= 1'b0;
    end else if(N1427) begin
      mem_q[1275] <= mem_n[1275];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1274] <= 1'b0;
    end else if(N1427) begin
      mem_q[1274] <= mem_n[1274];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1273] <= 1'b0;
    end else if(N1427) begin
      mem_q[1273] <= mem_n[1273];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1272] <= 1'b0;
    end else if(N1427) begin
      mem_q[1272] <= mem_n[1272];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1271] <= 1'b0;
    end else if(N1427) begin
      mem_q[1271] <= mem_n[1271];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1270] <= 1'b0;
    end else if(N1427) begin
      mem_q[1270] <= mem_n[1270];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1269] <= 1'b0;
    end else if(N1427) begin
      mem_q[1269] <= mem_n[1269];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1268] <= 1'b0;
    end else if(N1427) begin
      mem_q[1268] <= mem_n[1268];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1267] <= 1'b0;
    end else if(N1427) begin
      mem_q[1267] <= mem_n[1267];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1266] <= 1'b0;
    end else if(N1427) begin
      mem_q[1266] <= mem_n[1266];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1265] <= 1'b0;
    end else if(N1427) begin
      mem_q[1265] <= mem_n[1265];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1264] <= 1'b0;
    end else if(N1427) begin
      mem_q[1264] <= mem_n[1264];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1263] <= 1'b0;
    end else if(N1427) begin
      mem_q[1263] <= mem_n[1263];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1262] <= 1'b0;
    end else if(N1427) begin
      mem_q[1262] <= mem_n[1262];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1261] <= 1'b0;
    end else if(N1427) begin
      mem_q[1261] <= mem_n[1261];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1260] <= 1'b0;
    end else if(N1427) begin
      mem_q[1260] <= mem_n[1260];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1259] <= 1'b0;
    end else if(N1427) begin
      mem_q[1259] <= mem_n[1259];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1258] <= 1'b0;
    end else if(N1427) begin
      mem_q[1258] <= mem_n[1258];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1257] <= 1'b0;
    end else if(N1427) begin
      mem_q[1257] <= mem_n[1257];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1256] <= 1'b0;
    end else if(N1427) begin
      mem_q[1256] <= mem_n[1256];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1255] <= 1'b0;
    end else if(N1427) begin
      mem_q[1255] <= mem_n[1255];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1254] <= 1'b0;
    end else if(N1427) begin
      mem_q[1254] <= mem_n[1254];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1253] <= 1'b0;
    end else if(N1427) begin
      mem_q[1253] <= mem_n[1253];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1252] <= 1'b0;
    end else if(N1427) begin
      mem_q[1252] <= mem_n[1252];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1251] <= 1'b0;
    end else if(N1427) begin
      mem_q[1251] <= mem_n[1251];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1250] <= 1'b0;
    end else if(N1427) begin
      mem_q[1250] <= mem_n[1250];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1249] <= 1'b0;
    end else if(N1427) begin
      mem_q[1249] <= mem_n[1249];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1248] <= 1'b0;
    end else if(N1427) begin
      mem_q[1248] <= mem_n[1248];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1247] <= 1'b0;
    end else if(N1427) begin
      mem_q[1247] <= mem_n[1247];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1246] <= 1'b0;
    end else if(N1427) begin
      mem_q[1246] <= mem_n[1246];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1245] <= 1'b0;
    end else if(N1427) begin
      mem_q[1245] <= mem_n[1245];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1244] <= 1'b0;
    end else if(N1427) begin
      mem_q[1244] <= mem_n[1244];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1243] <= 1'b0;
    end else if(N1427) begin
      mem_q[1243] <= mem_n[1243];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1242] <= 1'b0;
    end else if(N1427) begin
      mem_q[1242] <= mem_n[1242];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1241] <= 1'b0;
    end else if(N1427) begin
      mem_q[1241] <= mem_n[1241];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1240] <= 1'b0;
    end else if(N1427) begin
      mem_q[1240] <= mem_n[1240];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1239] <= 1'b0;
    end else if(N1427) begin
      mem_q[1239] <= mem_n[1239];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1238] <= 1'b0;
    end else if(N1427) begin
      mem_q[1238] <= mem_n[1238];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1237] <= 1'b0;
    end else if(N1427) begin
      mem_q[1237] <= mem_n[1237];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1236] <= 1'b0;
    end else if(N1427) begin
      mem_q[1236] <= mem_n[1236];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1235] <= 1'b0;
    end else if(N1427) begin
      mem_q[1235] <= mem_n[1235];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1234] <= 1'b0;
    end else if(N1427) begin
      mem_q[1234] <= mem_n[1234];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1233] <= 1'b0;
    end else if(N1427) begin
      mem_q[1233] <= mem_n[1233];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1232] <= 1'b0;
    end else if(N1427) begin
      mem_q[1232] <= mem_n[1232];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1231] <= 1'b0;
    end else if(N1427) begin
      mem_q[1231] <= mem_n[1231];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1230] <= 1'b0;
    end else if(N1427) begin
      mem_q[1230] <= mem_n[1230];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1229] <= 1'b0;
    end else if(N1427) begin
      mem_q[1229] <= mem_n[1229];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1228] <= 1'b0;
    end else if(N1427) begin
      mem_q[1228] <= mem_n[1228];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1227] <= 1'b0;
    end else if(N1427) begin
      mem_q[1227] <= mem_n[1227];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1226] <= 1'b0;
    end else if(N1427) begin
      mem_q[1226] <= mem_n[1226];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1225] <= 1'b0;
    end else if(N1427) begin
      mem_q[1225] <= mem_n[1225];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1224] <= 1'b0;
    end else if(N1427) begin
      mem_q[1224] <= mem_n[1224];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1223] <= 1'b0;
    end else if(N1427) begin
      mem_q[1223] <= mem_n[1223];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1222] <= 1'b0;
    end else if(N1427) begin
      mem_q[1222] <= mem_n[1222];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1221] <= 1'b0;
    end else if(N1427) begin
      mem_q[1221] <= mem_n[1221];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1220] <= 1'b0;
    end else if(N1427) begin
      mem_q[1220] <= mem_n[1220];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1219] <= 1'b0;
    end else if(N1427) begin
      mem_q[1219] <= mem_n[1219];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1218] <= 1'b0;
    end else if(N1427) begin
      mem_q[1218] <= mem_n[1218];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1217] <= 1'b0;
    end else if(N1427) begin
      mem_q[1217] <= mem_n[1217];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1216] <= 1'b0;
    end else if(N1427) begin
      mem_q[1216] <= mem_n[1216];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1215] <= 1'b0;
    end else if(N1427) begin
      mem_q[1215] <= mem_n[1215];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1214] <= 1'b0;
    end else if(N1427) begin
      mem_q[1214] <= mem_n[1214];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1213] <= 1'b0;
    end else if(N1427) begin
      mem_q[1213] <= mem_n[1213];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1212] <= 1'b0;
    end else if(N1427) begin
      mem_q[1212] <= mem_n[1212];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1211] <= 1'b0;
    end else if(N1427) begin
      mem_q[1211] <= mem_n[1211];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1210] <= 1'b0;
    end else if(N1427) begin
      mem_q[1210] <= mem_n[1210];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1209] <= 1'b0;
    end else if(N1427) begin
      mem_q[1209] <= mem_n[1209];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1208] <= 1'b0;
    end else if(N1427) begin
      mem_q[1208] <= mem_n[1208];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1207] <= 1'b0;
    end else if(N1427) begin
      mem_q[1207] <= mem_n[1207];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1206] <= 1'b0;
    end else if(N1427) begin
      mem_q[1206] <= mem_n[1206];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1205] <= 1'b0;
    end else if(N1427) begin
      mem_q[1205] <= mem_n[1205];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1204] <= 1'b0;
    end else if(N1427) begin
      mem_q[1204] <= mem_n[1204];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1203] <= 1'b0;
    end else if(N1427) begin
      mem_q[1203] <= mem_n[1203];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1202] <= 1'b0;
    end else if(N1427) begin
      mem_q[1202] <= mem_n[1202];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1201] <= 1'b0;
    end else if(N1427) begin
      mem_q[1201] <= mem_n[1201];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1200] <= 1'b0;
    end else if(N1427) begin
      mem_q[1200] <= mem_n[1200];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1199] <= 1'b0;
    end else if(N1427) begin
      mem_q[1199] <= mem_n[1199];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1198] <= 1'b0;
    end else if(N1427) begin
      mem_q[1198] <= mem_n[1198];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1197] <= 1'b0;
    end else if(N1427) begin
      mem_q[1197] <= mem_n[1197];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1196] <= 1'b0;
    end else if(N1427) begin
      mem_q[1196] <= mem_n[1196];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1195] <= 1'b0;
    end else if(N1427) begin
      mem_q[1195] <= mem_n[1195];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1194] <= 1'b0;
    end else if(N1427) begin
      mem_q[1194] <= mem_n[1194];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1193] <= 1'b0;
    end else if(N1427) begin
      mem_q[1193] <= mem_n[1193];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1192] <= 1'b0;
    end else if(N1427) begin
      mem_q[1192] <= mem_n[1192];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1191] <= 1'b0;
    end else if(N1427) begin
      mem_q[1191] <= mem_n[1191];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1190] <= 1'b0;
    end else if(N1427) begin
      mem_q[1190] <= mem_n[1190];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1189] <= 1'b0;
    end else if(N1427) begin
      mem_q[1189] <= mem_n[1189];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1188] <= 1'b0;
    end else if(N1427) begin
      mem_q[1188] <= mem_n[1188];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1187] <= 1'b0;
    end else if(N1427) begin
      mem_q[1187] <= mem_n[1187];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1186] <= 1'b0;
    end else if(N1427) begin
      mem_q[1186] <= mem_n[1186];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1185] <= 1'b0;
    end else if(N1427) begin
      mem_q[1185] <= mem_n[1185];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1184] <= 1'b0;
    end else if(N1427) begin
      mem_q[1184] <= mem_n[1184];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1183] <= 1'b0;
    end else if(N1427) begin
      mem_q[1183] <= mem_n[1183];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1182] <= 1'b0;
    end else if(N1427) begin
      mem_q[1182] <= mem_n[1182];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1181] <= 1'b0;
    end else if(N1427) begin
      mem_q[1181] <= mem_n[1181];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1180] <= 1'b0;
    end else if(N1427) begin
      mem_q[1180] <= mem_n[1180];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1179] <= 1'b0;
    end else if(N1427) begin
      mem_q[1179] <= mem_n[1179];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1178] <= 1'b0;
    end else if(N1427) begin
      mem_q[1178] <= mem_n[1178];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1177] <= 1'b0;
    end else if(N1427) begin
      mem_q[1177] <= mem_n[1177];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1176] <= 1'b0;
    end else if(N1427) begin
      mem_q[1176] <= mem_n[1176];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1175] <= 1'b0;
    end else if(N1427) begin
      mem_q[1175] <= mem_n[1175];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1174] <= 1'b0;
    end else if(N1427) begin
      mem_q[1174] <= mem_n[1174];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1173] <= 1'b0;
    end else if(N1427) begin
      mem_q[1173] <= mem_n[1173];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1172] <= 1'b0;
    end else if(N1427) begin
      mem_q[1172] <= mem_n[1172];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1171] <= 1'b0;
    end else if(N1427) begin
      mem_q[1171] <= mem_n[1171];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1170] <= 1'b0;
    end else if(N1427) begin
      mem_q[1170] <= mem_n[1170];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1169] <= 1'b0;
    end else if(N1427) begin
      mem_q[1169] <= mem_n[1169];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1168] <= 1'b0;
    end else if(N1427) begin
      mem_q[1168] <= mem_n[1168];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1167] <= 1'b0;
    end else if(N1427) begin
      mem_q[1167] <= mem_n[1167];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1166] <= 1'b0;
    end else if(N1427) begin
      mem_q[1166] <= mem_n[1166];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1165] <= 1'b0;
    end else if(N1427) begin
      mem_q[1165] <= mem_n[1165];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1164] <= 1'b0;
    end else if(N1427) begin
      mem_q[1164] <= mem_n[1164];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1163] <= 1'b0;
    end else if(N1427) begin
      mem_q[1163] <= mem_n[1163];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1162] <= 1'b0;
    end else if(N1427) begin
      mem_q[1162] <= mem_n[1162];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1161] <= 1'b0;
    end else if(N1427) begin
      mem_q[1161] <= mem_n[1161];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1160] <= 1'b0;
    end else if(N1427) begin
      mem_q[1160] <= mem_n[1160];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1159] <= 1'b0;
    end else if(N1427) begin
      mem_q[1159] <= mem_n[1159];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1158] <= 1'b0;
    end else if(N1427) begin
      mem_q[1158] <= mem_n[1158];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1157] <= 1'b0;
    end else if(N1427) begin
      mem_q[1157] <= mem_n[1157];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1156] <= 1'b0;
    end else if(N1427) begin
      mem_q[1156] <= mem_n[1156];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1155] <= 1'b0;
    end else if(N1427) begin
      mem_q[1155] <= mem_n[1155];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1154] <= 1'b0;
    end else if(N1427) begin
      mem_q[1154] <= mem_n[1154];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1153] <= 1'b0;
    end else if(N1427) begin
      mem_q[1153] <= mem_n[1153];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1152] <= 1'b0;
    end else if(N1427) begin
      mem_q[1152] <= mem_n[1152];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1151] <= 1'b0;
    end else if(N1427) begin
      mem_q[1151] <= mem_n[1151];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1150] <= 1'b0;
    end else if(N1427) begin
      mem_q[1150] <= mem_n[1150];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1149] <= 1'b0;
    end else if(N1427) begin
      mem_q[1149] <= mem_n[1149];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1148] <= 1'b0;
    end else if(N1427) begin
      mem_q[1148] <= mem_n[1148];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1147] <= 1'b0;
    end else if(N1427) begin
      mem_q[1147] <= mem_n[1147];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1146] <= 1'b0;
    end else if(N1427) begin
      mem_q[1146] <= mem_n[1146];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1145] <= 1'b0;
    end else if(N1427) begin
      mem_q[1145] <= mem_n[1145];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1144] <= 1'b0;
    end else if(N1427) begin
      mem_q[1144] <= mem_n[1144];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1143] <= 1'b0;
    end else if(N1427) begin
      mem_q[1143] <= mem_n[1143];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1142] <= 1'b0;
    end else if(N1427) begin
      mem_q[1142] <= mem_n[1142];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1141] <= 1'b0;
    end else if(N1427) begin
      mem_q[1141] <= mem_n[1141];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1140] <= 1'b0;
    end else if(N1427) begin
      mem_q[1140] <= mem_n[1140];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1139] <= 1'b0;
    end else if(N1427) begin
      mem_q[1139] <= mem_n[1139];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1138] <= 1'b0;
    end else if(N1427) begin
      mem_q[1138] <= mem_n[1138];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1137] <= 1'b0;
    end else if(N1427) begin
      mem_q[1137] <= mem_n[1137];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1136] <= 1'b0;
    end else if(N1427) begin
      mem_q[1136] <= mem_n[1136];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1135] <= 1'b0;
    end else if(N1427) begin
      mem_q[1135] <= mem_n[1135];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1134] <= 1'b0;
    end else if(N1427) begin
      mem_q[1134] <= mem_n[1134];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1133] <= 1'b0;
    end else if(N1427) begin
      mem_q[1133] <= mem_n[1133];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1132] <= 1'b0;
    end else if(N1427) begin
      mem_q[1132] <= mem_n[1132];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1131] <= 1'b0;
    end else if(N1427) begin
      mem_q[1131] <= mem_n[1131];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1130] <= 1'b0;
    end else if(N1427) begin
      mem_q[1130] <= mem_n[1130];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1129] <= 1'b0;
    end else if(N1427) begin
      mem_q[1129] <= mem_n[1129];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1128] <= 1'b0;
    end else if(N1427) begin
      mem_q[1128] <= mem_n[1128];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1127] <= 1'b0;
    end else if(N1427) begin
      mem_q[1127] <= mem_n[1127];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1126] <= 1'b0;
    end else if(N1427) begin
      mem_q[1126] <= mem_n[1126];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1125] <= 1'b0;
    end else if(N1427) begin
      mem_q[1125] <= mem_n[1125];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1124] <= 1'b0;
    end else if(N1427) begin
      mem_q[1124] <= mem_n[1124];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1123] <= 1'b0;
    end else if(N1427) begin
      mem_q[1123] <= mem_n[1123];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1122] <= 1'b0;
    end else if(N1427) begin
      mem_q[1122] <= mem_n[1122];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1121] <= 1'b0;
    end else if(N1427) begin
      mem_q[1121] <= mem_n[1121];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1120] <= 1'b0;
    end else if(N1427) begin
      mem_q[1120] <= mem_n[1120];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1119] <= 1'b0;
    end else if(N1427) begin
      mem_q[1119] <= mem_n[1119];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1118] <= 1'b0;
    end else if(N1427) begin
      mem_q[1118] <= mem_n[1118];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1117] <= 1'b0;
    end else if(N1427) begin
      mem_q[1117] <= mem_n[1117];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1116] <= 1'b0;
    end else if(N1427) begin
      mem_q[1116] <= mem_n[1116];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1115] <= 1'b0;
    end else if(N1427) begin
      mem_q[1115] <= mem_n[1115];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1114] <= 1'b0;
    end else if(N1427) begin
      mem_q[1114] <= mem_n[1114];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1113] <= 1'b0;
    end else if(N1427) begin
      mem_q[1113] <= mem_n[1113];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1112] <= 1'b0;
    end else if(N1427) begin
      mem_q[1112] <= mem_n[1112];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1111] <= 1'b0;
    end else if(N1427) begin
      mem_q[1111] <= mem_n[1111];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1110] <= 1'b0;
    end else if(N1427) begin
      mem_q[1110] <= mem_n[1110];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1109] <= 1'b0;
    end else if(N1427) begin
      mem_q[1109] <= mem_n[1109];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1108] <= 1'b0;
    end else if(N1427) begin
      mem_q[1108] <= mem_n[1108];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1107] <= 1'b0;
    end else if(N1427) begin
      mem_q[1107] <= mem_n[1107];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1106] <= 1'b0;
    end else if(N1427) begin
      mem_q[1106] <= mem_n[1106];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1105] <= 1'b0;
    end else if(N1427) begin
      mem_q[1105] <= mem_n[1105];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1104] <= 1'b0;
    end else if(N1427) begin
      mem_q[1104] <= mem_n[1104];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1103] <= 1'b0;
    end else if(N1427) begin
      mem_q[1103] <= mem_n[1103];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1102] <= 1'b0;
    end else if(N1427) begin
      mem_q[1102] <= mem_n[1102];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1101] <= 1'b0;
    end else if(N1427) begin
      mem_q[1101] <= mem_n[1101];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1100] <= 1'b0;
    end else if(N1427) begin
      mem_q[1100] <= mem_n[1100];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1099] <= 1'b0;
    end else if(N1427) begin
      mem_q[1099] <= mem_n[1099];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1098] <= 1'b0;
    end else if(N1427) begin
      mem_q[1098] <= mem_n[1098];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1097] <= 1'b0;
    end else if(N1427) begin
      mem_q[1097] <= mem_n[1097];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1096] <= 1'b0;
    end else if(N1427) begin
      mem_q[1096] <= mem_n[1096];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1095] <= 1'b0;
    end else if(N1427) begin
      mem_q[1095] <= mem_n[1095];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1094] <= 1'b0;
    end else if(N1427) begin
      mem_q[1094] <= mem_n[1094];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1093] <= 1'b0;
    end else if(N1427) begin
      mem_q[1093] <= mem_n[1093];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1092] <= 1'b0;
    end else if(N1427) begin
      mem_q[1092] <= mem_n[1092];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1091] <= 1'b0;
    end else if(N1427) begin
      mem_q[1091] <= mem_n[1091];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1090] <= 1'b0;
    end else if(N1427) begin
      mem_q[1090] <= mem_n[1090];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1089] <= 1'b0;
    end else if(N1427) begin
      mem_q[1089] <= mem_n[1089];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1088] <= 1'b0;
    end else if(N1427) begin
      mem_q[1088] <= mem_n[1088];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1087] <= 1'b0;
    end else if(N1427) begin
      mem_q[1087] <= mem_n[1087];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1086] <= 1'b0;
    end else if(N1427) begin
      mem_q[1086] <= mem_n[1086];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1085] <= 1'b0;
    end else if(N1427) begin
      mem_q[1085] <= mem_n[1085];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1084] <= 1'b0;
    end else if(N1427) begin
      mem_q[1084] <= mem_n[1084];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1083] <= 1'b0;
    end else if(N1427) begin
      mem_q[1083] <= mem_n[1083];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1082] <= 1'b0;
    end else if(N1427) begin
      mem_q[1082] <= mem_n[1082];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1081] <= 1'b0;
    end else if(N1427) begin
      mem_q[1081] <= mem_n[1081];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1080] <= 1'b0;
    end else if(N1427) begin
      mem_q[1080] <= mem_n[1080];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1079] <= 1'b0;
    end else if(N1427) begin
      mem_q[1079] <= mem_n[1079];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1078] <= 1'b0;
    end else if(N1427) begin
      mem_q[1078] <= mem_n[1078];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1077] <= 1'b0;
    end else if(N1427) begin
      mem_q[1077] <= mem_n[1077];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1076] <= 1'b0;
    end else if(N1427) begin
      mem_q[1076] <= mem_n[1076];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1075] <= 1'b0;
    end else if(N1427) begin
      mem_q[1075] <= mem_n[1075];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1074] <= 1'b0;
    end else if(N1427) begin
      mem_q[1074] <= mem_n[1074];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1073] <= 1'b0;
    end else if(N1427) begin
      mem_q[1073] <= mem_n[1073];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1072] <= 1'b0;
    end else if(N1427) begin
      mem_q[1072] <= mem_n[1072];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1071] <= 1'b0;
    end else if(N1427) begin
      mem_q[1071] <= mem_n[1071];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1070] <= 1'b0;
    end else if(N1427) begin
      mem_q[1070] <= mem_n[1070];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1069] <= 1'b0;
    end else if(N1427) begin
      mem_q[1069] <= mem_n[1069];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1068] <= 1'b0;
    end else if(N1427) begin
      mem_q[1068] <= mem_n[1068];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1067] <= 1'b0;
    end else if(N1427) begin
      mem_q[1067] <= mem_n[1067];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1066] <= 1'b0;
    end else if(N1427) begin
      mem_q[1066] <= mem_n[1066];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1065] <= 1'b0;
    end else if(N1427) begin
      mem_q[1065] <= mem_n[1065];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1064] <= 1'b0;
    end else if(N1427) begin
      mem_q[1064] <= mem_n[1064];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1063] <= 1'b0;
    end else if(N1427) begin
      mem_q[1063] <= mem_n[1063];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1062] <= 1'b0;
    end else if(N1427) begin
      mem_q[1062] <= mem_n[1062];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1061] <= 1'b0;
    end else if(N1427) begin
      mem_q[1061] <= mem_n[1061];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1060] <= 1'b0;
    end else if(N1427) begin
      mem_q[1060] <= mem_n[1060];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1059] <= 1'b0;
    end else if(N1427) begin
      mem_q[1059] <= mem_n[1059];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1058] <= 1'b0;
    end else if(N1427) begin
      mem_q[1058] <= mem_n[1058];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1057] <= 1'b0;
    end else if(N1427) begin
      mem_q[1057] <= mem_n[1057];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1056] <= 1'b0;
    end else if(N1427) begin
      mem_q[1056] <= mem_n[1056];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1055] <= 1'b0;
    end else if(N1427) begin
      mem_q[1055] <= mem_n[1055];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1054] <= 1'b0;
    end else if(N1427) begin
      mem_q[1054] <= mem_n[1054];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1053] <= 1'b0;
    end else if(N1427) begin
      mem_q[1053] <= mem_n[1053];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1052] <= 1'b0;
    end else if(N1427) begin
      mem_q[1052] <= mem_n[1052];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1051] <= 1'b0;
    end else if(N1427) begin
      mem_q[1051] <= mem_n[1051];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1050] <= 1'b0;
    end else if(N1427) begin
      mem_q[1050] <= mem_n[1050];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1049] <= 1'b0;
    end else if(N1427) begin
      mem_q[1049] <= mem_n[1049];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1048] <= 1'b0;
    end else if(N1427) begin
      mem_q[1048] <= mem_n[1048];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1047] <= 1'b0;
    end else if(N1427) begin
      mem_q[1047] <= mem_n[1047];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1046] <= 1'b0;
    end else if(N1427) begin
      mem_q[1046] <= mem_n[1046];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1045] <= 1'b0;
    end else if(N1427) begin
      mem_q[1045] <= mem_n[1045];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1044] <= 1'b0;
    end else if(N1427) begin
      mem_q[1044] <= mem_n[1044];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1043] <= 1'b0;
    end else if(N1427) begin
      mem_q[1043] <= mem_n[1043];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1042] <= 1'b0;
    end else if(N1427) begin
      mem_q[1042] <= mem_n[1042];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1041] <= 1'b0;
    end else if(N1427) begin
      mem_q[1041] <= mem_n[1041];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1040] <= 1'b0;
    end else if(N1427) begin
      mem_q[1040] <= mem_n[1040];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1039] <= 1'b0;
    end else if(N1427) begin
      mem_q[1039] <= mem_n[1039];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1038] <= 1'b0;
    end else if(N1427) begin
      mem_q[1038] <= mem_n[1038];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1037] <= 1'b0;
    end else if(N1427) begin
      mem_q[1037] <= mem_n[1037];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1036] <= 1'b0;
    end else if(N1427) begin
      mem_q[1036] <= mem_n[1036];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1035] <= 1'b0;
    end else if(N1427) begin
      mem_q[1035] <= mem_n[1035];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1034] <= 1'b0;
    end else if(N1427) begin
      mem_q[1034] <= mem_n[1034];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1033] <= 1'b0;
    end else if(N1427) begin
      mem_q[1033] <= mem_n[1033];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1032] <= 1'b0;
    end else if(N1427) begin
      mem_q[1032] <= mem_n[1032];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1031] <= 1'b0;
    end else if(N1427) begin
      mem_q[1031] <= mem_n[1031];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1030] <= 1'b0;
    end else if(N1427) begin
      mem_q[1030] <= mem_n[1030];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1029] <= 1'b0;
    end else if(N1427) begin
      mem_q[1029] <= mem_n[1029];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1028] <= 1'b0;
    end else if(N1427) begin
      mem_q[1028] <= mem_n[1028];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1027] <= 1'b0;
    end else if(N1427) begin
      mem_q[1027] <= mem_n[1027];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1026] <= 1'b0;
    end else if(N1427) begin
      mem_q[1026] <= mem_n[1026];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1025] <= 1'b0;
    end else if(N1427) begin
      mem_q[1025] <= mem_n[1025];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1024] <= 1'b0;
    end else if(N1427) begin
      mem_q[1024] <= mem_n[1024];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1023] <= 1'b0;
    end else if(N1427) begin
      mem_q[1023] <= mem_n[1023];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1022] <= 1'b0;
    end else if(N1427) begin
      mem_q[1022] <= mem_n[1022];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1021] <= 1'b0;
    end else if(N1427) begin
      mem_q[1021] <= mem_n[1021];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1020] <= 1'b0;
    end else if(N1427) begin
      mem_q[1020] <= mem_n[1020];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1019] <= 1'b0;
    end else if(N1427) begin
      mem_q[1019] <= mem_n[1019];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1018] <= 1'b0;
    end else if(N1427) begin
      mem_q[1018] <= mem_n[1018];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1017] <= 1'b0;
    end else if(N1427) begin
      mem_q[1017] <= mem_n[1017];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1016] <= 1'b0;
    end else if(N1427) begin
      mem_q[1016] <= mem_n[1016];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1015] <= 1'b0;
    end else if(N1427) begin
      mem_q[1015] <= mem_n[1015];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1014] <= 1'b0;
    end else if(N1427) begin
      mem_q[1014] <= mem_n[1014];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1013] <= 1'b0;
    end else if(N1427) begin
      mem_q[1013] <= mem_n[1013];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1012] <= 1'b0;
    end else if(N1427) begin
      mem_q[1012] <= mem_n[1012];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1011] <= 1'b0;
    end else if(N1427) begin
      mem_q[1011] <= mem_n[1011];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1010] <= 1'b0;
    end else if(N1427) begin
      mem_q[1010] <= mem_n[1010];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1009] <= 1'b0;
    end else if(N1427) begin
      mem_q[1009] <= mem_n[1009];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1008] <= 1'b0;
    end else if(N1427) begin
      mem_q[1008] <= mem_n[1008];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1007] <= 1'b0;
    end else if(N1427) begin
      mem_q[1007] <= mem_n[1007];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1006] <= 1'b0;
    end else if(N1427) begin
      mem_q[1006] <= mem_n[1006];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1005] <= 1'b0;
    end else if(N1427) begin
      mem_q[1005] <= mem_n[1005];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1004] <= 1'b0;
    end else if(N1427) begin
      mem_q[1004] <= mem_n[1004];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1003] <= 1'b0;
    end else if(N1427) begin
      mem_q[1003] <= mem_n[1003];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1002] <= 1'b0;
    end else if(N1427) begin
      mem_q[1002] <= mem_n[1002];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1001] <= 1'b0;
    end else if(N1427) begin
      mem_q[1001] <= mem_n[1001];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1000] <= 1'b0;
    end else if(N1427) begin
      mem_q[1000] <= mem_n[1000];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[999] <= 1'b0;
    end else if(N1427) begin
      mem_q[999] <= mem_n[999];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[998] <= 1'b0;
    end else if(N1427) begin
      mem_q[998] <= mem_n[998];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[997] <= 1'b0;
    end else if(N1427) begin
      mem_q[997] <= mem_n[997];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[996] <= 1'b0;
    end else if(N1427) begin
      mem_q[996] <= mem_n[996];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[995] <= 1'b0;
    end else if(N1427) begin
      mem_q[995] <= mem_n[995];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[994] <= 1'b0;
    end else if(N1427) begin
      mem_q[994] <= mem_n[994];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[993] <= 1'b0;
    end else if(N1427) begin
      mem_q[993] <= mem_n[993];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[992] <= 1'b0;
    end else if(N1427) begin
      mem_q[992] <= mem_n[992];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[991] <= 1'b0;
    end else if(N1427) begin
      mem_q[991] <= mem_n[991];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[990] <= 1'b0;
    end else if(N1427) begin
      mem_q[990] <= mem_n[990];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[989] <= 1'b0;
    end else if(N1427) begin
      mem_q[989] <= mem_n[989];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[988] <= 1'b0;
    end else if(N1427) begin
      mem_q[988] <= mem_n[988];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[987] <= 1'b0;
    end else if(N1427) begin
      mem_q[987] <= mem_n[987];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[986] <= 1'b0;
    end else if(N1427) begin
      mem_q[986] <= mem_n[986];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[985] <= 1'b0;
    end else if(N1427) begin
      mem_q[985] <= mem_n[985];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[984] <= 1'b0;
    end else if(N1427) begin
      mem_q[984] <= mem_n[984];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[983] <= 1'b0;
    end else if(N1427) begin
      mem_q[983] <= mem_n[983];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[982] <= 1'b0;
    end else if(N1427) begin
      mem_q[982] <= mem_n[982];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[981] <= 1'b0;
    end else if(N1427) begin
      mem_q[981] <= mem_n[981];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[980] <= 1'b0;
    end else if(N1427) begin
      mem_q[980] <= mem_n[980];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[979] <= 1'b0;
    end else if(N1427) begin
      mem_q[979] <= mem_n[979];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[978] <= 1'b0;
    end else if(N1427) begin
      mem_q[978] <= mem_n[978];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[977] <= 1'b0;
    end else if(N1427) begin
      mem_q[977] <= mem_n[977];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[976] <= 1'b0;
    end else if(N1427) begin
      mem_q[976] <= mem_n[976];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[975] <= 1'b0;
    end else if(N1427) begin
      mem_q[975] <= mem_n[975];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[974] <= 1'b0;
    end else if(N1427) begin
      mem_q[974] <= mem_n[974];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[973] <= 1'b0;
    end else if(N1427) begin
      mem_q[973] <= mem_n[973];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[972] <= 1'b0;
    end else if(N1427) begin
      mem_q[972] <= mem_n[972];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[971] <= 1'b0;
    end else if(N1427) begin
      mem_q[971] <= mem_n[971];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[970] <= 1'b0;
    end else if(N1427) begin
      mem_q[970] <= mem_n[970];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[969] <= 1'b0;
    end else if(N1427) begin
      mem_q[969] <= mem_n[969];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[968] <= 1'b0;
    end else if(N1427) begin
      mem_q[968] <= mem_n[968];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[967] <= 1'b0;
    end else if(N1427) begin
      mem_q[967] <= mem_n[967];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[966] <= 1'b0;
    end else if(N1427) begin
      mem_q[966] <= mem_n[966];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[965] <= 1'b0;
    end else if(N1427) begin
      mem_q[965] <= mem_n[965];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[964] <= 1'b0;
    end else if(N1427) begin
      mem_q[964] <= mem_n[964];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[963] <= 1'b0;
    end else if(N1427) begin
      mem_q[963] <= mem_n[963];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[962] <= 1'b0;
    end else if(N1427) begin
      mem_q[962] <= mem_n[962];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[961] <= 1'b0;
    end else if(N1427) begin
      mem_q[961] <= mem_n[961];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[960] <= 1'b0;
    end else if(N1427) begin
      mem_q[960] <= mem_n[960];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[959] <= 1'b0;
    end else if(N1427) begin
      mem_q[959] <= mem_n[959];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[958] <= 1'b0;
    end else if(N1427) begin
      mem_q[958] <= mem_n[958];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[957] <= 1'b0;
    end else if(N1427) begin
      mem_q[957] <= mem_n[957];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[956] <= 1'b0;
    end else if(N1427) begin
      mem_q[956] <= mem_n[956];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[955] <= 1'b0;
    end else if(N1427) begin
      mem_q[955] <= mem_n[955];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[954] <= 1'b0;
    end else if(N1427) begin
      mem_q[954] <= mem_n[954];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[953] <= 1'b0;
    end else if(N1427) begin
      mem_q[953] <= mem_n[953];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[952] <= 1'b0;
    end else if(N1427) begin
      mem_q[952] <= mem_n[952];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[951] <= 1'b0;
    end else if(N1427) begin
      mem_q[951] <= mem_n[951];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[950] <= 1'b0;
    end else if(N1427) begin
      mem_q[950] <= mem_n[950];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[949] <= 1'b0;
    end else if(N1427) begin
      mem_q[949] <= mem_n[949];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[948] <= 1'b0;
    end else if(N1427) begin
      mem_q[948] <= mem_n[948];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[947] <= 1'b0;
    end else if(N1427) begin
      mem_q[947] <= mem_n[947];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[946] <= 1'b0;
    end else if(N1427) begin
      mem_q[946] <= mem_n[946];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[945] <= 1'b0;
    end else if(N1427) begin
      mem_q[945] <= mem_n[945];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[944] <= 1'b0;
    end else if(N1427) begin
      mem_q[944] <= mem_n[944];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[943] <= 1'b0;
    end else if(N1427) begin
      mem_q[943] <= mem_n[943];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[942] <= 1'b0;
    end else if(N1427) begin
      mem_q[942] <= mem_n[942];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[941] <= 1'b0;
    end else if(N1427) begin
      mem_q[941] <= mem_n[941];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[940] <= 1'b0;
    end else if(N1427) begin
      mem_q[940] <= mem_n[940];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[939] <= 1'b0;
    end else if(N1427) begin
      mem_q[939] <= mem_n[939];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[938] <= 1'b0;
    end else if(N1427) begin
      mem_q[938] <= mem_n[938];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[937] <= 1'b0;
    end else if(N1427) begin
      mem_q[937] <= mem_n[937];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[936] <= 1'b0;
    end else if(N1427) begin
      mem_q[936] <= mem_n[936];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[935] <= 1'b0;
    end else if(N1427) begin
      mem_q[935] <= mem_n[935];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[934] <= 1'b0;
    end else if(N1427) begin
      mem_q[934] <= mem_n[934];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[933] <= 1'b0;
    end else if(N1427) begin
      mem_q[933] <= mem_n[933];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[932] <= 1'b0;
    end else if(N1427) begin
      mem_q[932] <= mem_n[932];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[931] <= 1'b0;
    end else if(N1427) begin
      mem_q[931] <= mem_n[931];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[930] <= 1'b0;
    end else if(N1427) begin
      mem_q[930] <= mem_n[930];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[929] <= 1'b0;
    end else if(N1427) begin
      mem_q[929] <= mem_n[929];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[928] <= 1'b0;
    end else if(N1427) begin
      mem_q[928] <= mem_n[928];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[927] <= 1'b0;
    end else if(N1427) begin
      mem_q[927] <= mem_n[927];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[926] <= 1'b0;
    end else if(N1427) begin
      mem_q[926] <= mem_n[926];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[925] <= 1'b0;
    end else if(N1427) begin
      mem_q[925] <= mem_n[925];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[924] <= 1'b0;
    end else if(N1427) begin
      mem_q[924] <= mem_n[924];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[923] <= 1'b0;
    end else if(N1427) begin
      mem_q[923] <= mem_n[923];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[922] <= 1'b0;
    end else if(N1427) begin
      mem_q[922] <= mem_n[922];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[921] <= 1'b0;
    end else if(N1427) begin
      mem_q[921] <= mem_n[921];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[920] <= 1'b0;
    end else if(N1427) begin
      mem_q[920] <= mem_n[920];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[919] <= 1'b0;
    end else if(N1427) begin
      mem_q[919] <= mem_n[919];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[918] <= 1'b0;
    end else if(N1427) begin
      mem_q[918] <= mem_n[918];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[917] <= 1'b0;
    end else if(N1427) begin
      mem_q[917] <= mem_n[917];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[916] <= 1'b0;
    end else if(N1427) begin
      mem_q[916] <= mem_n[916];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[915] <= 1'b0;
    end else if(N1427) begin
      mem_q[915] <= mem_n[915];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[914] <= 1'b0;
    end else if(N1427) begin
      mem_q[914] <= mem_n[914];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[913] <= 1'b0;
    end else if(N1427) begin
      mem_q[913] <= mem_n[913];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[912] <= 1'b0;
    end else if(N1427) begin
      mem_q[912] <= mem_n[912];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[911] <= 1'b0;
    end else if(N1427) begin
      mem_q[911] <= mem_n[911];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[910] <= 1'b0;
    end else if(N1427) begin
      mem_q[910] <= mem_n[910];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[909] <= 1'b0;
    end else if(N1427) begin
      mem_q[909] <= mem_n[909];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[908] <= 1'b0;
    end else if(N1427) begin
      mem_q[908] <= mem_n[908];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[907] <= 1'b0;
    end else if(N1427) begin
      mem_q[907] <= mem_n[907];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[906] <= 1'b0;
    end else if(N1427) begin
      mem_q[906] <= mem_n[906];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[905] <= 1'b0;
    end else if(N1427) begin
      mem_q[905] <= mem_n[905];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[904] <= 1'b0;
    end else if(N1427) begin
      mem_q[904] <= mem_n[904];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[903] <= 1'b0;
    end else if(N1427) begin
      mem_q[903] <= mem_n[903];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[902] <= 1'b0;
    end else if(N1427) begin
      mem_q[902] <= mem_n[902];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[901] <= 1'b0;
    end else if(N1427) begin
      mem_q[901] <= mem_n[901];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[900] <= 1'b0;
    end else if(N1427) begin
      mem_q[900] <= mem_n[900];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[899] <= 1'b0;
    end else if(N1427) begin
      mem_q[899] <= mem_n[899];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[898] <= 1'b0;
    end else if(N1427) begin
      mem_q[898] <= mem_n[898];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[897] <= 1'b0;
    end else if(N1427) begin
      mem_q[897] <= mem_n[897];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[896] <= 1'b0;
    end else if(N1427) begin
      mem_q[896] <= mem_n[896];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[895] <= 1'b0;
    end else if(N1427) begin
      mem_q[895] <= mem_n[895];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[894] <= 1'b0;
    end else if(N1427) begin
      mem_q[894] <= mem_n[894];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[893] <= 1'b0;
    end else if(N1427) begin
      mem_q[893] <= mem_n[893];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[892] <= 1'b0;
    end else if(N1427) begin
      mem_q[892] <= mem_n[892];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[891] <= 1'b0;
    end else if(N1427) begin
      mem_q[891] <= mem_n[891];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[890] <= 1'b0;
    end else if(N1427) begin
      mem_q[890] <= mem_n[890];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[889] <= 1'b0;
    end else if(N1427) begin
      mem_q[889] <= mem_n[889];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[888] <= 1'b0;
    end else if(N1427) begin
      mem_q[888] <= mem_n[888];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[887] <= 1'b0;
    end else if(N1427) begin
      mem_q[887] <= mem_n[887];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[886] <= 1'b0;
    end else if(N1427) begin
      mem_q[886] <= mem_n[886];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[885] <= 1'b0;
    end else if(N1427) begin
      mem_q[885] <= mem_n[885];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[884] <= 1'b0;
    end else if(N1427) begin
      mem_q[884] <= mem_n[884];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[883] <= 1'b0;
    end else if(N1427) begin
      mem_q[883] <= mem_n[883];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[882] <= 1'b0;
    end else if(N1427) begin
      mem_q[882] <= mem_n[882];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[881] <= 1'b0;
    end else if(N1427) begin
      mem_q[881] <= mem_n[881];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[880] <= 1'b0;
    end else if(N1427) begin
      mem_q[880] <= mem_n[880];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[879] <= 1'b0;
    end else if(N1427) begin
      mem_q[879] <= mem_n[879];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[878] <= 1'b0;
    end else if(N1427) begin
      mem_q[878] <= mem_n[878];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[877] <= 1'b0;
    end else if(N1427) begin
      mem_q[877] <= mem_n[877];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[876] <= 1'b0;
    end else if(N1427) begin
      mem_q[876] <= mem_n[876];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[875] <= 1'b0;
    end else if(N1427) begin
      mem_q[875] <= mem_n[875];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[874] <= 1'b0;
    end else if(N1427) begin
      mem_q[874] <= mem_n[874];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[873] <= 1'b0;
    end else if(N1427) begin
      mem_q[873] <= mem_n[873];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[872] <= 1'b0;
    end else if(N1427) begin
      mem_q[872] <= mem_n[872];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[871] <= 1'b0;
    end else if(N1427) begin
      mem_q[871] <= mem_n[871];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[870] <= 1'b0;
    end else if(N1427) begin
      mem_q[870] <= mem_n[870];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[869] <= 1'b0;
    end else if(N1427) begin
      mem_q[869] <= mem_n[869];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[868] <= 1'b0;
    end else if(N1427) begin
      mem_q[868] <= mem_n[868];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[867] <= 1'b0;
    end else if(N1427) begin
      mem_q[867] <= mem_n[867];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[866] <= 1'b0;
    end else if(N1427) begin
      mem_q[866] <= mem_n[866];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[865] <= 1'b0;
    end else if(N1427) begin
      mem_q[865] <= mem_n[865];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[864] <= 1'b0;
    end else if(N1427) begin
      mem_q[864] <= mem_n[864];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[863] <= 1'b0;
    end else if(N1427) begin
      mem_q[863] <= mem_n[863];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[862] <= 1'b0;
    end else if(N1427) begin
      mem_q[862] <= mem_n[862];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[861] <= 1'b0;
    end else if(N1427) begin
      mem_q[861] <= mem_n[861];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[860] <= 1'b0;
    end else if(N1427) begin
      mem_q[860] <= mem_n[860];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[859] <= 1'b0;
    end else if(N1427) begin
      mem_q[859] <= mem_n[859];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[858] <= 1'b0;
    end else if(N1427) begin
      mem_q[858] <= mem_n[858];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[857] <= 1'b0;
    end else if(N1427) begin
      mem_q[857] <= mem_n[857];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[856] <= 1'b0;
    end else if(N1427) begin
      mem_q[856] <= mem_n[856];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[855] <= 1'b0;
    end else if(N1427) begin
      mem_q[855] <= mem_n[855];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[854] <= 1'b0;
    end else if(N1427) begin
      mem_q[854] <= mem_n[854];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[853] <= 1'b0;
    end else if(N1427) begin
      mem_q[853] <= mem_n[853];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[852] <= 1'b0;
    end else if(N1427) begin
      mem_q[852] <= mem_n[852];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[851] <= 1'b0;
    end else if(N1427) begin
      mem_q[851] <= mem_n[851];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[850] <= 1'b0;
    end else if(N1427) begin
      mem_q[850] <= mem_n[850];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[849] <= 1'b0;
    end else if(N1427) begin
      mem_q[849] <= mem_n[849];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[848] <= 1'b0;
    end else if(N1427) begin
      mem_q[848] <= mem_n[848];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[847] <= 1'b0;
    end else if(N1427) begin
      mem_q[847] <= mem_n[847];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[846] <= 1'b0;
    end else if(N1427) begin
      mem_q[846] <= mem_n[846];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[845] <= 1'b0;
    end else if(N1427) begin
      mem_q[845] <= mem_n[845];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[844] <= 1'b0;
    end else if(N1427) begin
      mem_q[844] <= mem_n[844];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[843] <= 1'b0;
    end else if(N1427) begin
      mem_q[843] <= mem_n[843];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[842] <= 1'b0;
    end else if(N1427) begin
      mem_q[842] <= mem_n[842];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[841] <= 1'b0;
    end else if(N1427) begin
      mem_q[841] <= mem_n[841];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[840] <= 1'b0;
    end else if(N1427) begin
      mem_q[840] <= mem_n[840];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[839] <= 1'b0;
    end else if(N1427) begin
      mem_q[839] <= mem_n[839];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[838] <= 1'b0;
    end else if(N1427) begin
      mem_q[838] <= mem_n[838];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[837] <= 1'b0;
    end else if(N1427) begin
      mem_q[837] <= mem_n[837];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[836] <= 1'b0;
    end else if(N1427) begin
      mem_q[836] <= mem_n[836];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[835] <= 1'b0;
    end else if(N1427) begin
      mem_q[835] <= mem_n[835];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[834] <= 1'b0;
    end else if(N1427) begin
      mem_q[834] <= mem_n[834];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[833] <= 1'b0;
    end else if(N1427) begin
      mem_q[833] <= mem_n[833];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[832] <= 1'b0;
    end else if(N1427) begin
      mem_q[832] <= mem_n[832];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[831] <= 1'b0;
    end else if(N1427) begin
      mem_q[831] <= mem_n[831];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[830] <= 1'b0;
    end else if(N1427) begin
      mem_q[830] <= mem_n[830];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[829] <= 1'b0;
    end else if(N1427) begin
      mem_q[829] <= mem_n[829];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[828] <= 1'b0;
    end else if(N1427) begin
      mem_q[828] <= mem_n[828];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[827] <= 1'b0;
    end else if(N1427) begin
      mem_q[827] <= mem_n[827];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[826] <= 1'b0;
    end else if(N1427) begin
      mem_q[826] <= mem_n[826];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[825] <= 1'b0;
    end else if(N1427) begin
      mem_q[825] <= mem_n[825];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[824] <= 1'b0;
    end else if(N1427) begin
      mem_q[824] <= mem_n[824];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[823] <= 1'b0;
    end else if(N1427) begin
      mem_q[823] <= mem_n[823];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[822] <= 1'b0;
    end else if(N1427) begin
      mem_q[822] <= mem_n[822];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[821] <= 1'b0;
    end else if(N1427) begin
      mem_q[821] <= mem_n[821];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[820] <= 1'b0;
    end else if(N1427) begin
      mem_q[820] <= mem_n[820];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[819] <= 1'b0;
    end else if(N1427) begin
      mem_q[819] <= mem_n[819];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[818] <= 1'b0;
    end else if(N1427) begin
      mem_q[818] <= mem_n[818];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[817] <= 1'b0;
    end else if(N1427) begin
      mem_q[817] <= mem_n[817];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[816] <= 1'b0;
    end else if(N1427) begin
      mem_q[816] <= mem_n[816];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[815] <= 1'b0;
    end else if(N1427) begin
      mem_q[815] <= mem_n[815];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[814] <= 1'b0;
    end else if(N1427) begin
      mem_q[814] <= mem_n[814];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[813] <= 1'b0;
    end else if(N1427) begin
      mem_q[813] <= mem_n[813];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[812] <= 1'b0;
    end else if(N1427) begin
      mem_q[812] <= mem_n[812];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[811] <= 1'b0;
    end else if(N1427) begin
      mem_q[811] <= mem_n[811];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[810] <= 1'b0;
    end else if(N1427) begin
      mem_q[810] <= mem_n[810];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[809] <= 1'b0;
    end else if(N1427) begin
      mem_q[809] <= mem_n[809];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[808] <= 1'b0;
    end else if(N1427) begin
      mem_q[808] <= mem_n[808];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[807] <= 1'b0;
    end else if(N1427) begin
      mem_q[807] <= mem_n[807];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[806] <= 1'b0;
    end else if(N1427) begin
      mem_q[806] <= mem_n[806];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[805] <= 1'b0;
    end else if(N1427) begin
      mem_q[805] <= mem_n[805];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[804] <= 1'b0;
    end else if(N1427) begin
      mem_q[804] <= mem_n[804];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[803] <= 1'b0;
    end else if(N1427) begin
      mem_q[803] <= mem_n[803];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[802] <= 1'b0;
    end else if(N1427) begin
      mem_q[802] <= mem_n[802];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[801] <= 1'b0;
    end else if(N1427) begin
      mem_q[801] <= mem_n[801];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[800] <= 1'b0;
    end else if(N1427) begin
      mem_q[800] <= mem_n[800];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[799] <= 1'b0;
    end else if(N1427) begin
      mem_q[799] <= mem_n[799];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[798] <= 1'b0;
    end else if(N1427) begin
      mem_q[798] <= mem_n[798];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[797] <= 1'b0;
    end else if(N1427) begin
      mem_q[797] <= mem_n[797];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[796] <= 1'b0;
    end else if(N1427) begin
      mem_q[796] <= mem_n[796];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[795] <= 1'b0;
    end else if(N1427) begin
      mem_q[795] <= mem_n[795];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[794] <= 1'b0;
    end else if(N1427) begin
      mem_q[794] <= mem_n[794];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[793] <= 1'b0;
    end else if(N1427) begin
      mem_q[793] <= mem_n[793];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[792] <= 1'b0;
    end else if(N1427) begin
      mem_q[792] <= mem_n[792];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[791] <= 1'b0;
    end else if(N1427) begin
      mem_q[791] <= mem_n[791];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[790] <= 1'b0;
    end else if(N1427) begin
      mem_q[790] <= mem_n[790];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[789] <= 1'b0;
    end else if(N1427) begin
      mem_q[789] <= mem_n[789];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[788] <= 1'b0;
    end else if(N1427) begin
      mem_q[788] <= mem_n[788];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[787] <= 1'b0;
    end else if(N1427) begin
      mem_q[787] <= mem_n[787];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[786] <= 1'b0;
    end else if(N1427) begin
      mem_q[786] <= mem_n[786];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[785] <= 1'b0;
    end else if(N1427) begin
      mem_q[785] <= mem_n[785];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[784] <= 1'b0;
    end else if(N1427) begin
      mem_q[784] <= mem_n[784];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[783] <= 1'b0;
    end else if(N1427) begin
      mem_q[783] <= mem_n[783];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[782] <= 1'b0;
    end else if(N1427) begin
      mem_q[782] <= mem_n[782];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[781] <= 1'b0;
    end else if(N1427) begin
      mem_q[781] <= mem_n[781];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[780] <= 1'b0;
    end else if(N1427) begin
      mem_q[780] <= mem_n[780];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[779] <= 1'b0;
    end else if(N1427) begin
      mem_q[779] <= mem_n[779];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[778] <= 1'b0;
    end else if(N1427) begin
      mem_q[778] <= mem_n[778];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[777] <= 1'b0;
    end else if(N1427) begin
      mem_q[777] <= mem_n[777];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[776] <= 1'b0;
    end else if(N1427) begin
      mem_q[776] <= mem_n[776];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[775] <= 1'b0;
    end else if(N1427) begin
      mem_q[775] <= mem_n[775];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[774] <= 1'b0;
    end else if(N1427) begin
      mem_q[774] <= mem_n[774];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[773] <= 1'b0;
    end else if(N1427) begin
      mem_q[773] <= mem_n[773];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[772] <= 1'b0;
    end else if(N1427) begin
      mem_q[772] <= mem_n[772];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[771] <= 1'b0;
    end else if(N1427) begin
      mem_q[771] <= mem_n[771];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[770] <= 1'b0;
    end else if(N1427) begin
      mem_q[770] <= mem_n[770];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[769] <= 1'b0;
    end else if(N1427) begin
      mem_q[769] <= mem_n[769];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[768] <= 1'b0;
    end else if(N1427) begin
      mem_q[768] <= mem_n[768];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[767] <= 1'b0;
    end else if(N1427) begin
      mem_q[767] <= mem_n[767];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[766] <= 1'b0;
    end else if(N1427) begin
      mem_q[766] <= mem_n[766];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[765] <= 1'b0;
    end else if(N1427) begin
      mem_q[765] <= mem_n[765];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[764] <= 1'b0;
    end else if(N1427) begin
      mem_q[764] <= mem_n[764];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[763] <= 1'b0;
    end else if(N1427) begin
      mem_q[763] <= mem_n[763];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[762] <= 1'b0;
    end else if(N1427) begin
      mem_q[762] <= mem_n[762];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[761] <= 1'b0;
    end else if(N1427) begin
      mem_q[761] <= mem_n[761];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[760] <= 1'b0;
    end else if(N1427) begin
      mem_q[760] <= mem_n[760];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[759] <= 1'b0;
    end else if(N1427) begin
      mem_q[759] <= mem_n[759];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[758] <= 1'b0;
    end else if(N1427) begin
      mem_q[758] <= mem_n[758];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[757] <= 1'b0;
    end else if(N1427) begin
      mem_q[757] <= mem_n[757];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[756] <= 1'b0;
    end else if(N1427) begin
      mem_q[756] <= mem_n[756];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[755] <= 1'b0;
    end else if(N1427) begin
      mem_q[755] <= mem_n[755];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[754] <= 1'b0;
    end else if(N1427) begin
      mem_q[754] <= mem_n[754];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[753] <= 1'b0;
    end else if(N1427) begin
      mem_q[753] <= mem_n[753];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[752] <= 1'b0;
    end else if(N1427) begin
      mem_q[752] <= mem_n[752];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[751] <= 1'b0;
    end else if(N1427) begin
      mem_q[751] <= mem_n[751];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[750] <= 1'b0;
    end else if(N1427) begin
      mem_q[750] <= mem_n[750];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[749] <= 1'b0;
    end else if(N1427) begin
      mem_q[749] <= mem_n[749];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[748] <= 1'b0;
    end else if(N1427) begin
      mem_q[748] <= mem_n[748];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[747] <= 1'b0;
    end else if(N1427) begin
      mem_q[747] <= mem_n[747];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[746] <= 1'b0;
    end else if(N1427) begin
      mem_q[746] <= mem_n[746];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[745] <= 1'b0;
    end else if(N1427) begin
      mem_q[745] <= mem_n[745];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[744] <= 1'b0;
    end else if(N1427) begin
      mem_q[744] <= mem_n[744];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[743] <= 1'b0;
    end else if(N1427) begin
      mem_q[743] <= mem_n[743];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[742] <= 1'b0;
    end else if(N1427) begin
      mem_q[742] <= mem_n[742];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[741] <= 1'b0;
    end else if(N1427) begin
      mem_q[741] <= mem_n[741];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[740] <= 1'b0;
    end else if(N1427) begin
      mem_q[740] <= mem_n[740];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[739] <= 1'b0;
    end else if(N1427) begin
      mem_q[739] <= mem_n[739];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[738] <= 1'b0;
    end else if(N1427) begin
      mem_q[738] <= mem_n[738];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[737] <= 1'b0;
    end else if(N1427) begin
      mem_q[737] <= mem_n[737];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[736] <= 1'b0;
    end else if(N1427) begin
      mem_q[736] <= mem_n[736];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[735] <= 1'b0;
    end else if(N1427) begin
      mem_q[735] <= mem_n[735];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[734] <= 1'b0;
    end else if(N1427) begin
      mem_q[734] <= mem_n[734];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[733] <= 1'b0;
    end else if(N1427) begin
      mem_q[733] <= mem_n[733];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[732] <= 1'b0;
    end else if(N1427) begin
      mem_q[732] <= mem_n[732];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[731] <= 1'b0;
    end else if(N1427) begin
      mem_q[731] <= mem_n[731];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[730] <= 1'b0;
    end else if(N1427) begin
      mem_q[730] <= mem_n[730];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[729] <= 1'b0;
    end else if(N1427) begin
      mem_q[729] <= mem_n[729];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[728] <= 1'b0;
    end else if(N1427) begin
      mem_q[728] <= mem_n[728];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[727] <= 1'b0;
    end else if(N1427) begin
      mem_q[727] <= mem_n[727];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[726] <= 1'b0;
    end else if(N1427) begin
      mem_q[726] <= mem_n[726];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[725] <= 1'b0;
    end else if(N1427) begin
      mem_q[725] <= mem_n[725];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[724] <= 1'b0;
    end else if(N1427) begin
      mem_q[724] <= mem_n[724];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[723] <= 1'b0;
    end else if(N1427) begin
      mem_q[723] <= mem_n[723];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[722] <= 1'b0;
    end else if(N1427) begin
      mem_q[722] <= mem_n[722];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[721] <= 1'b0;
    end else if(N1427) begin
      mem_q[721] <= mem_n[721];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[720] <= 1'b0;
    end else if(N1427) begin
      mem_q[720] <= mem_n[720];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[719] <= 1'b0;
    end else if(N1427) begin
      mem_q[719] <= mem_n[719];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[718] <= 1'b0;
    end else if(N1427) begin
      mem_q[718] <= mem_n[718];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[717] <= 1'b0;
    end else if(N1427) begin
      mem_q[717] <= mem_n[717];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[716] <= 1'b0;
    end else if(N1427) begin
      mem_q[716] <= mem_n[716];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[715] <= 1'b0;
    end else if(N1427) begin
      mem_q[715] <= mem_n[715];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[714] <= 1'b0;
    end else if(N1427) begin
      mem_q[714] <= mem_n[714];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[713] <= 1'b0;
    end else if(N1427) begin
      mem_q[713] <= mem_n[713];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[712] <= 1'b0;
    end else if(N1427) begin
      mem_q[712] <= mem_n[712];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[711] <= 1'b0;
    end else if(N1427) begin
      mem_q[711] <= mem_n[711];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[710] <= 1'b0;
    end else if(N1427) begin
      mem_q[710] <= mem_n[710];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[709] <= 1'b0;
    end else if(N1427) begin
      mem_q[709] <= mem_n[709];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[708] <= 1'b0;
    end else if(N1427) begin
      mem_q[708] <= mem_n[708];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[707] <= 1'b0;
    end else if(N1427) begin
      mem_q[707] <= mem_n[707];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[706] <= 1'b0;
    end else if(N1427) begin
      mem_q[706] <= mem_n[706];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[705] <= 1'b0;
    end else if(N1427) begin
      mem_q[705] <= mem_n[705];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[704] <= 1'b0;
    end else if(N1427) begin
      mem_q[704] <= mem_n[704];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[703] <= 1'b0;
    end else if(N1427) begin
      mem_q[703] <= mem_n[703];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[702] <= 1'b0;
    end else if(N1427) begin
      mem_q[702] <= mem_n[702];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[701] <= 1'b0;
    end else if(N1427) begin
      mem_q[701] <= mem_n[701];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[700] <= 1'b0;
    end else if(N1427) begin
      mem_q[700] <= mem_n[700];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[699] <= 1'b0;
    end else if(N1427) begin
      mem_q[699] <= mem_n[699];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[698] <= 1'b0;
    end else if(N1427) begin
      mem_q[698] <= mem_n[698];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[697] <= 1'b0;
    end else if(N1427) begin
      mem_q[697] <= mem_n[697];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[696] <= 1'b0;
    end else if(N1427) begin
      mem_q[696] <= mem_n[696];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[695] <= 1'b0;
    end else if(N1427) begin
      mem_q[695] <= mem_n[695];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[694] <= 1'b0;
    end else if(N1427) begin
      mem_q[694] <= mem_n[694];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[693] <= 1'b0;
    end else if(N1427) begin
      mem_q[693] <= mem_n[693];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[692] <= 1'b0;
    end else if(N1427) begin
      mem_q[692] <= mem_n[692];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[691] <= 1'b0;
    end else if(N1427) begin
      mem_q[691] <= mem_n[691];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[690] <= 1'b0;
    end else if(N1427) begin
      mem_q[690] <= mem_n[690];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[689] <= 1'b0;
    end else if(N1427) begin
      mem_q[689] <= mem_n[689];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[688] <= 1'b0;
    end else if(N1427) begin
      mem_q[688] <= mem_n[688];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[687] <= 1'b0;
    end else if(N1427) begin
      mem_q[687] <= mem_n[687];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[686] <= 1'b0;
    end else if(N1427) begin
      mem_q[686] <= mem_n[686];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[685] <= 1'b0;
    end else if(N1427) begin
      mem_q[685] <= mem_n[685];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[684] <= 1'b0;
    end else if(N1427) begin
      mem_q[684] <= mem_n[684];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[683] <= 1'b0;
    end else if(N1427) begin
      mem_q[683] <= mem_n[683];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[682] <= 1'b0;
    end else if(N1427) begin
      mem_q[682] <= mem_n[682];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[681] <= 1'b0;
    end else if(N1427) begin
      mem_q[681] <= mem_n[681];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[680] <= 1'b0;
    end else if(N1427) begin
      mem_q[680] <= mem_n[680];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[679] <= 1'b0;
    end else if(N1427) begin
      mem_q[679] <= mem_n[679];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[678] <= 1'b0;
    end else if(N1427) begin
      mem_q[678] <= mem_n[678];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[677] <= 1'b0;
    end else if(N1427) begin
      mem_q[677] <= mem_n[677];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[676] <= 1'b0;
    end else if(N1427) begin
      mem_q[676] <= mem_n[676];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[675] <= 1'b0;
    end else if(N1427) begin
      mem_q[675] <= mem_n[675];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[674] <= 1'b0;
    end else if(N1427) begin
      mem_q[674] <= mem_n[674];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[673] <= 1'b0;
    end else if(N1427) begin
      mem_q[673] <= mem_n[673];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[672] <= 1'b0;
    end else if(N1427) begin
      mem_q[672] <= mem_n[672];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[671] <= 1'b0;
    end else if(N1427) begin
      mem_q[671] <= mem_n[671];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[670] <= 1'b0;
    end else if(N1427) begin
      mem_q[670] <= mem_n[670];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[669] <= 1'b0;
    end else if(N1427) begin
      mem_q[669] <= mem_n[669];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[668] <= 1'b0;
    end else if(N1427) begin
      mem_q[668] <= mem_n[668];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[667] <= 1'b0;
    end else if(N1427) begin
      mem_q[667] <= mem_n[667];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[666] <= 1'b0;
    end else if(N1427) begin
      mem_q[666] <= mem_n[666];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[665] <= 1'b0;
    end else if(N1427) begin
      mem_q[665] <= mem_n[665];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[664] <= 1'b0;
    end else if(N1427) begin
      mem_q[664] <= mem_n[664];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[663] <= 1'b0;
    end else if(N1427) begin
      mem_q[663] <= mem_n[663];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[662] <= 1'b0;
    end else if(N1427) begin
      mem_q[662] <= mem_n[662];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[661] <= 1'b0;
    end else if(N1427) begin
      mem_q[661] <= mem_n[661];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[660] <= 1'b0;
    end else if(N1427) begin
      mem_q[660] <= mem_n[660];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[659] <= 1'b0;
    end else if(N1427) begin
      mem_q[659] <= mem_n[659];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[658] <= 1'b0;
    end else if(N1427) begin
      mem_q[658] <= mem_n[658];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[657] <= 1'b0;
    end else if(N1427) begin
      mem_q[657] <= mem_n[657];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[656] <= 1'b0;
    end else if(N1427) begin
      mem_q[656] <= mem_n[656];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[655] <= 1'b0;
    end else if(N1427) begin
      mem_q[655] <= mem_n[655];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[654] <= 1'b0;
    end else if(N1427) begin
      mem_q[654] <= mem_n[654];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[653] <= 1'b0;
    end else if(N1427) begin
      mem_q[653] <= mem_n[653];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[652] <= 1'b0;
    end else if(N1427) begin
      mem_q[652] <= mem_n[652];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[651] <= 1'b0;
    end else if(N1427) begin
      mem_q[651] <= mem_n[651];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[650] <= 1'b0;
    end else if(N1427) begin
      mem_q[650] <= mem_n[650];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[649] <= 1'b0;
    end else if(N1427) begin
      mem_q[649] <= mem_n[649];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[648] <= 1'b0;
    end else if(N1427) begin
      mem_q[648] <= mem_n[648];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[647] <= 1'b0;
    end else if(N1427) begin
      mem_q[647] <= mem_n[647];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[646] <= 1'b0;
    end else if(N1427) begin
      mem_q[646] <= mem_n[646];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[645] <= 1'b0;
    end else if(N1427) begin
      mem_q[645] <= mem_n[645];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[644] <= 1'b0;
    end else if(N1427) begin
      mem_q[644] <= mem_n[644];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[643] <= 1'b0;
    end else if(N1427) begin
      mem_q[643] <= mem_n[643];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[642] <= 1'b0;
    end else if(N1427) begin
      mem_q[642] <= mem_n[642];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[641] <= 1'b0;
    end else if(N1427) begin
      mem_q[641] <= mem_n[641];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[640] <= 1'b0;
    end else if(N1427) begin
      mem_q[640] <= mem_n[640];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[639] <= 1'b0;
    end else if(N1427) begin
      mem_q[639] <= mem_n[639];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[638] <= 1'b0;
    end else if(N1427) begin
      mem_q[638] <= mem_n[638];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[637] <= 1'b0;
    end else if(N1427) begin
      mem_q[637] <= mem_n[637];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[636] <= 1'b0;
    end else if(N1427) begin
      mem_q[636] <= mem_n[636];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[635] <= 1'b0;
    end else if(N1427) begin
      mem_q[635] <= mem_n[635];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[634] <= 1'b0;
    end else if(N1427) begin
      mem_q[634] <= mem_n[634];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[633] <= 1'b0;
    end else if(N1427) begin
      mem_q[633] <= mem_n[633];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[632] <= 1'b0;
    end else if(N1427) begin
      mem_q[632] <= mem_n[632];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[631] <= 1'b0;
    end else if(N1427) begin
      mem_q[631] <= mem_n[631];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[630] <= 1'b0;
    end else if(N1427) begin
      mem_q[630] <= mem_n[630];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[629] <= 1'b0;
    end else if(N1427) begin
      mem_q[629] <= mem_n[629];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[628] <= 1'b0;
    end else if(N1427) begin
      mem_q[628] <= mem_n[628];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[627] <= 1'b0;
    end else if(N1427) begin
      mem_q[627] <= mem_n[627];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[626] <= 1'b0;
    end else if(N1427) begin
      mem_q[626] <= mem_n[626];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[625] <= 1'b0;
    end else if(N1427) begin
      mem_q[625] <= mem_n[625];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[624] <= 1'b0;
    end else if(N1427) begin
      mem_q[624] <= mem_n[624];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[623] <= 1'b0;
    end else if(N1427) begin
      mem_q[623] <= mem_n[623];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[622] <= 1'b0;
    end else if(N1427) begin
      mem_q[622] <= mem_n[622];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[621] <= 1'b0;
    end else if(N1427) begin
      mem_q[621] <= mem_n[621];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[620] <= 1'b0;
    end else if(N1427) begin
      mem_q[620] <= mem_n[620];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[619] <= 1'b0;
    end else if(N1427) begin
      mem_q[619] <= mem_n[619];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[618] <= 1'b0;
    end else if(N1427) begin
      mem_q[618] <= mem_n[618];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[617] <= 1'b0;
    end else if(N1427) begin
      mem_q[617] <= mem_n[617];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[616] <= 1'b0;
    end else if(N1427) begin
      mem_q[616] <= mem_n[616];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[615] <= 1'b0;
    end else if(N1427) begin
      mem_q[615] <= mem_n[615];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[614] <= 1'b0;
    end else if(N1427) begin
      mem_q[614] <= mem_n[614];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[613] <= 1'b0;
    end else if(N1427) begin
      mem_q[613] <= mem_n[613];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[612] <= 1'b0;
    end else if(N1427) begin
      mem_q[612] <= mem_n[612];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[611] <= 1'b0;
    end else if(N1427) begin
      mem_q[611] <= mem_n[611];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[610] <= 1'b0;
    end else if(N1427) begin
      mem_q[610] <= mem_n[610];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[609] <= 1'b0;
    end else if(N1427) begin
      mem_q[609] <= mem_n[609];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[608] <= 1'b0;
    end else if(N1427) begin
      mem_q[608] <= mem_n[608];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[607] <= 1'b0;
    end else if(N1427) begin
      mem_q[607] <= mem_n[607];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[606] <= 1'b0;
    end else if(N1427) begin
      mem_q[606] <= mem_n[606];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[605] <= 1'b0;
    end else if(N1427) begin
      mem_q[605] <= mem_n[605];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[604] <= 1'b0;
    end else if(N1427) begin
      mem_q[604] <= mem_n[604];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[603] <= 1'b0;
    end else if(N1427) begin
      mem_q[603] <= mem_n[603];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[602] <= 1'b0;
    end else if(N1427) begin
      mem_q[602] <= mem_n[602];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[601] <= 1'b0;
    end else if(N1427) begin
      mem_q[601] <= mem_n[601];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[600] <= 1'b0;
    end else if(N1427) begin
      mem_q[600] <= mem_n[600];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[599] <= 1'b0;
    end else if(N1427) begin
      mem_q[599] <= mem_n[599];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[598] <= 1'b0;
    end else if(N1427) begin
      mem_q[598] <= mem_n[598];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[597] <= 1'b0;
    end else if(N1427) begin
      mem_q[597] <= mem_n[597];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[596] <= 1'b0;
    end else if(N1427) begin
      mem_q[596] <= mem_n[596];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[595] <= 1'b0;
    end else if(N1427) begin
      mem_q[595] <= mem_n[595];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[594] <= 1'b0;
    end else if(N1427) begin
      mem_q[594] <= mem_n[594];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[593] <= 1'b0;
    end else if(N1427) begin
      mem_q[593] <= mem_n[593];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[592] <= 1'b0;
    end else if(N1427) begin
      mem_q[592] <= mem_n[592];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[591] <= 1'b0;
    end else if(N1427) begin
      mem_q[591] <= mem_n[591];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[590] <= 1'b0;
    end else if(N1427) begin
      mem_q[590] <= mem_n[590];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[589] <= 1'b0;
    end else if(N1427) begin
      mem_q[589] <= mem_n[589];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[588] <= 1'b0;
    end else if(N1427) begin
      mem_q[588] <= mem_n[588];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[587] <= 1'b0;
    end else if(N1427) begin
      mem_q[587] <= mem_n[587];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[586] <= 1'b0;
    end else if(N1427) begin
      mem_q[586] <= mem_n[586];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[585] <= 1'b0;
    end else if(N1427) begin
      mem_q[585] <= mem_n[585];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[584] <= 1'b0;
    end else if(N1427) begin
      mem_q[584] <= mem_n[584];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[583] <= 1'b0;
    end else if(N1427) begin
      mem_q[583] <= mem_n[583];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[582] <= 1'b0;
    end else if(N1427) begin
      mem_q[582] <= mem_n[582];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[581] <= 1'b0;
    end else if(N1427) begin
      mem_q[581] <= mem_n[581];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[580] <= 1'b0;
    end else if(N1427) begin
      mem_q[580] <= mem_n[580];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[579] <= 1'b0;
    end else if(N1427) begin
      mem_q[579] <= mem_n[579];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[578] <= 1'b0;
    end else if(N1427) begin
      mem_q[578] <= mem_n[578];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[577] <= 1'b0;
    end else if(N1427) begin
      mem_q[577] <= mem_n[577];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[576] <= 1'b0;
    end else if(N1427) begin
      mem_q[576] <= mem_n[576];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[575] <= 1'b0;
    end else if(N1427) begin
      mem_q[575] <= mem_n[575];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[574] <= 1'b0;
    end else if(N1427) begin
      mem_q[574] <= mem_n[574];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[573] <= 1'b0;
    end else if(N1427) begin
      mem_q[573] <= mem_n[573];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[572] <= 1'b0;
    end else if(N1427) begin
      mem_q[572] <= mem_n[572];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[571] <= 1'b0;
    end else if(N1427) begin
      mem_q[571] <= mem_n[571];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[570] <= 1'b0;
    end else if(N1427) begin
      mem_q[570] <= mem_n[570];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[569] <= 1'b0;
    end else if(N1427) begin
      mem_q[569] <= mem_n[569];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[568] <= 1'b0;
    end else if(N1427) begin
      mem_q[568] <= mem_n[568];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[567] <= 1'b0;
    end else if(N1427) begin
      mem_q[567] <= mem_n[567];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[566] <= 1'b0;
    end else if(N1427) begin
      mem_q[566] <= mem_n[566];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[565] <= 1'b0;
    end else if(N1427) begin
      mem_q[565] <= mem_n[565];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[564] <= 1'b0;
    end else if(N1427) begin
      mem_q[564] <= mem_n[564];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[563] <= 1'b0;
    end else if(N1427) begin
      mem_q[563] <= mem_n[563];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[562] <= 1'b0;
    end else if(N1427) begin
      mem_q[562] <= mem_n[562];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[561] <= 1'b0;
    end else if(N1427) begin
      mem_q[561] <= mem_n[561];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[560] <= 1'b0;
    end else if(N1427) begin
      mem_q[560] <= mem_n[560];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[559] <= 1'b0;
    end else if(N1427) begin
      mem_q[559] <= mem_n[559];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[558] <= 1'b0;
    end else if(N1427) begin
      mem_q[558] <= mem_n[558];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[557] <= 1'b0;
    end else if(N1427) begin
      mem_q[557] <= mem_n[557];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[556] <= 1'b0;
    end else if(N1427) begin
      mem_q[556] <= mem_n[556];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[555] <= 1'b0;
    end else if(N1427) begin
      mem_q[555] <= mem_n[555];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[554] <= 1'b0;
    end else if(N1427) begin
      mem_q[554] <= mem_n[554];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[553] <= 1'b0;
    end else if(N1427) begin
      mem_q[553] <= mem_n[553];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[552] <= 1'b0;
    end else if(N1427) begin
      mem_q[552] <= mem_n[552];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[551] <= 1'b0;
    end else if(N1427) begin
      mem_q[551] <= mem_n[551];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[550] <= 1'b0;
    end else if(N1427) begin
      mem_q[550] <= mem_n[550];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[549] <= 1'b0;
    end else if(N1427) begin
      mem_q[549] <= mem_n[549];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[548] <= 1'b0;
    end else if(N1427) begin
      mem_q[548] <= mem_n[548];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[547] <= 1'b0;
    end else if(N1427) begin
      mem_q[547] <= mem_n[547];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[546] <= 1'b0;
    end else if(N1427) begin
      mem_q[546] <= mem_n[546];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[545] <= 1'b0;
    end else if(N1427) begin
      mem_q[545] <= mem_n[545];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[544] <= 1'b0;
    end else if(N1427) begin
      mem_q[544] <= mem_n[544];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[543] <= 1'b0;
    end else if(N1427) begin
      mem_q[543] <= mem_n[543];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[542] <= 1'b0;
    end else if(N1427) begin
      mem_q[542] <= mem_n[542];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[541] <= 1'b0;
    end else if(N1427) begin
      mem_q[541] <= mem_n[541];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[540] <= 1'b0;
    end else if(N1427) begin
      mem_q[540] <= mem_n[540];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[539] <= 1'b0;
    end else if(N1427) begin
      mem_q[539] <= mem_n[539];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[538] <= 1'b0;
    end else if(N1427) begin
      mem_q[538] <= mem_n[538];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[537] <= 1'b0;
    end else if(N1427) begin
      mem_q[537] <= mem_n[537];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[536] <= 1'b0;
    end else if(N1427) begin
      mem_q[536] <= mem_n[536];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[535] <= 1'b0;
    end else if(N1427) begin
      mem_q[535] <= mem_n[535];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[534] <= 1'b0;
    end else if(N1427) begin
      mem_q[534] <= mem_n[534];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[533] <= 1'b0;
    end else if(N1427) begin
      mem_q[533] <= mem_n[533];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[532] <= 1'b0;
    end else if(N1427) begin
      mem_q[532] <= mem_n[532];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[531] <= 1'b0;
    end else if(N1427) begin
      mem_q[531] <= mem_n[531];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[530] <= 1'b0;
    end else if(N1427) begin
      mem_q[530] <= mem_n[530];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[529] <= 1'b0;
    end else if(N1427) begin
      mem_q[529] <= mem_n[529];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[528] <= 1'b0;
    end else if(N1427) begin
      mem_q[528] <= mem_n[528];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[527] <= 1'b0;
    end else if(N1427) begin
      mem_q[527] <= mem_n[527];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[526] <= 1'b0;
    end else if(N1427) begin
      mem_q[526] <= mem_n[526];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[525] <= 1'b0;
    end else if(N1427) begin
      mem_q[525] <= mem_n[525];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[524] <= 1'b0;
    end else if(N1427) begin
      mem_q[524] <= mem_n[524];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[523] <= 1'b0;
    end else if(N1427) begin
      mem_q[523] <= mem_n[523];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[522] <= 1'b0;
    end else if(N1427) begin
      mem_q[522] <= mem_n[522];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[521] <= 1'b0;
    end else if(N1427) begin
      mem_q[521] <= mem_n[521];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[520] <= 1'b0;
    end else if(N1427) begin
      mem_q[520] <= mem_n[520];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[519] <= 1'b0;
    end else if(N1427) begin
      mem_q[519] <= mem_n[519];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[518] <= 1'b0;
    end else if(N1427) begin
      mem_q[518] <= mem_n[518];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[517] <= 1'b0;
    end else if(N1427) begin
      mem_q[517] <= mem_n[517];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[516] <= 1'b0;
    end else if(N1427) begin
      mem_q[516] <= mem_n[516];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[515] <= 1'b0;
    end else if(N1427) begin
      mem_q[515] <= mem_n[515];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[514] <= 1'b0;
    end else if(N1427) begin
      mem_q[514] <= mem_n[514];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[513] <= 1'b0;
    end else if(N1427) begin
      mem_q[513] <= mem_n[513];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[512] <= 1'b0;
    end else if(N1427) begin
      mem_q[512] <= mem_n[512];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[511] <= 1'b0;
    end else if(N1427) begin
      mem_q[511] <= mem_n[511];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[510] <= 1'b0;
    end else if(N1427) begin
      mem_q[510] <= mem_n[510];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[509] <= 1'b0;
    end else if(N1427) begin
      mem_q[509] <= mem_n[509];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[508] <= 1'b0;
    end else if(N1427) begin
      mem_q[508] <= mem_n[508];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[507] <= 1'b0;
    end else if(N1427) begin
      mem_q[507] <= mem_n[507];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[506] <= 1'b0;
    end else if(N1427) begin
      mem_q[506] <= mem_n[506];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[505] <= 1'b0;
    end else if(N1427) begin
      mem_q[505] <= mem_n[505];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[504] <= 1'b0;
    end else if(N1427) begin
      mem_q[504] <= mem_n[504];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[503] <= 1'b0;
    end else if(N1427) begin
      mem_q[503] <= mem_n[503];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[502] <= 1'b0;
    end else if(N1427) begin
      mem_q[502] <= mem_n[502];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[501] <= 1'b0;
    end else if(N1427) begin
      mem_q[501] <= mem_n[501];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[500] <= 1'b0;
    end else if(N1427) begin
      mem_q[500] <= mem_n[500];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[499] <= 1'b0;
    end else if(N1427) begin
      mem_q[499] <= mem_n[499];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[498] <= 1'b0;
    end else if(N1427) begin
      mem_q[498] <= mem_n[498];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[497] <= 1'b0;
    end else if(N1427) begin
      mem_q[497] <= mem_n[497];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[496] <= 1'b0;
    end else if(N1427) begin
      mem_q[496] <= mem_n[496];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[495] <= 1'b0;
    end else if(N1427) begin
      mem_q[495] <= mem_n[495];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[494] <= 1'b0;
    end else if(N1427) begin
      mem_q[494] <= mem_n[494];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[493] <= 1'b0;
    end else if(N1427) begin
      mem_q[493] <= mem_n[493];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[492] <= 1'b0;
    end else if(N1427) begin
      mem_q[492] <= mem_n[492];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[491] <= 1'b0;
    end else if(N1427) begin
      mem_q[491] <= mem_n[491];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[490] <= 1'b0;
    end else if(N1427) begin
      mem_q[490] <= mem_n[490];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[489] <= 1'b0;
    end else if(N1427) begin
      mem_q[489] <= mem_n[489];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[488] <= 1'b0;
    end else if(N1427) begin
      mem_q[488] <= mem_n[488];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[487] <= 1'b0;
    end else if(N1427) begin
      mem_q[487] <= mem_n[487];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[486] <= 1'b0;
    end else if(N1427) begin
      mem_q[486] <= mem_n[486];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[485] <= 1'b0;
    end else if(N1427) begin
      mem_q[485] <= mem_n[485];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[484] <= 1'b0;
    end else if(N1427) begin
      mem_q[484] <= mem_n[484];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[483] <= 1'b0;
    end else if(N1427) begin
      mem_q[483] <= mem_n[483];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[482] <= 1'b0;
    end else if(N1427) begin
      mem_q[482] <= mem_n[482];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[481] <= 1'b0;
    end else if(N1427) begin
      mem_q[481] <= mem_n[481];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[480] <= 1'b0;
    end else if(N1427) begin
      mem_q[480] <= mem_n[480];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[479] <= 1'b0;
    end else if(N1427) begin
      mem_q[479] <= mem_n[479];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[478] <= 1'b0;
    end else if(N1427) begin
      mem_q[478] <= mem_n[478];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[477] <= 1'b0;
    end else if(N1427) begin
      mem_q[477] <= mem_n[477];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[476] <= 1'b0;
    end else if(N1427) begin
      mem_q[476] <= mem_n[476];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[475] <= 1'b0;
    end else if(N1427) begin
      mem_q[475] <= mem_n[475];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[474] <= 1'b0;
    end else if(N1427) begin
      mem_q[474] <= mem_n[474];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[473] <= 1'b0;
    end else if(N1427) begin
      mem_q[473] <= mem_n[473];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[472] <= 1'b0;
    end else if(N1427) begin
      mem_q[472] <= mem_n[472];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[471] <= 1'b0;
    end else if(N1427) begin
      mem_q[471] <= mem_n[471];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[470] <= 1'b0;
    end else if(N1427) begin
      mem_q[470] <= mem_n[470];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[469] <= 1'b0;
    end else if(N1427) begin
      mem_q[469] <= mem_n[469];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[468] <= 1'b0;
    end else if(N1427) begin
      mem_q[468] <= mem_n[468];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[467] <= 1'b0;
    end else if(N1427) begin
      mem_q[467] <= mem_n[467];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[466] <= 1'b0;
    end else if(N1427) begin
      mem_q[466] <= mem_n[466];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[465] <= 1'b0;
    end else if(N1427) begin
      mem_q[465] <= mem_n[465];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[464] <= 1'b0;
    end else if(N1427) begin
      mem_q[464] <= mem_n[464];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[463] <= 1'b0;
    end else if(N1427) begin
      mem_q[463] <= mem_n[463];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[462] <= 1'b0;
    end else if(N1427) begin
      mem_q[462] <= mem_n[462];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[461] <= 1'b0;
    end else if(N1427) begin
      mem_q[461] <= mem_n[461];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[460] <= 1'b0;
    end else if(N1427) begin
      mem_q[460] <= mem_n[460];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[459] <= 1'b0;
    end else if(N1427) begin
      mem_q[459] <= mem_n[459];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[458] <= 1'b0;
    end else if(N1427) begin
      mem_q[458] <= mem_n[458];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[457] <= 1'b0;
    end else if(N1427) begin
      mem_q[457] <= mem_n[457];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[456] <= 1'b0;
    end else if(N1427) begin
      mem_q[456] <= mem_n[456];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[455] <= 1'b0;
    end else if(N1427) begin
      mem_q[455] <= mem_n[455];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[454] <= 1'b0;
    end else if(N1427) begin
      mem_q[454] <= mem_n[454];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[453] <= 1'b0;
    end else if(N1427) begin
      mem_q[453] <= mem_n[453];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[452] <= 1'b0;
    end else if(N1427) begin
      mem_q[452] <= mem_n[452];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[451] <= 1'b0;
    end else if(N1427) begin
      mem_q[451] <= mem_n[451];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[450] <= 1'b0;
    end else if(N1427) begin
      mem_q[450] <= mem_n[450];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[449] <= 1'b0;
    end else if(N1427) begin
      mem_q[449] <= mem_n[449];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[448] <= 1'b0;
    end else if(N1427) begin
      mem_q[448] <= mem_n[448];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[447] <= 1'b0;
    end else if(N1427) begin
      mem_q[447] <= mem_n[447];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[446] <= 1'b0;
    end else if(N1427) begin
      mem_q[446] <= mem_n[446];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[445] <= 1'b0;
    end else if(N1427) begin
      mem_q[445] <= mem_n[445];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[444] <= 1'b0;
    end else if(N1427) begin
      mem_q[444] <= mem_n[444];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[443] <= 1'b0;
    end else if(N1427) begin
      mem_q[443] <= mem_n[443];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[442] <= 1'b0;
    end else if(N1427) begin
      mem_q[442] <= mem_n[442];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[441] <= 1'b0;
    end else if(N1427) begin
      mem_q[441] <= mem_n[441];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[440] <= 1'b0;
    end else if(N1427) begin
      mem_q[440] <= mem_n[440];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[439] <= 1'b0;
    end else if(N1427) begin
      mem_q[439] <= mem_n[439];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[438] <= 1'b0;
    end else if(N1427) begin
      mem_q[438] <= mem_n[438];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[437] <= 1'b0;
    end else if(N1427) begin
      mem_q[437] <= mem_n[437];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[436] <= 1'b0;
    end else if(N1427) begin
      mem_q[436] <= mem_n[436];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[435] <= 1'b0;
    end else if(N1427) begin
      mem_q[435] <= mem_n[435];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[434] <= 1'b0;
    end else if(N1427) begin
      mem_q[434] <= mem_n[434];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[433] <= 1'b0;
    end else if(N1427) begin
      mem_q[433] <= mem_n[433];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[432] <= 1'b0;
    end else if(N1427) begin
      mem_q[432] <= mem_n[432];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[431] <= 1'b0;
    end else if(N1427) begin
      mem_q[431] <= mem_n[431];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[430] <= 1'b0;
    end else if(N1427) begin
      mem_q[430] <= mem_n[430];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[429] <= 1'b0;
    end else if(N1427) begin
      mem_q[429] <= mem_n[429];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[428] <= 1'b0;
    end else if(N1427) begin
      mem_q[428] <= mem_n[428];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[427] <= 1'b0;
    end else if(N1427) begin
      mem_q[427] <= mem_n[427];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[426] <= 1'b0;
    end else if(N1427) begin
      mem_q[426] <= mem_n[426];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[425] <= 1'b0;
    end else if(N1427) begin
      mem_q[425] <= mem_n[425];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[424] <= 1'b0;
    end else if(N1427) begin
      mem_q[424] <= mem_n[424];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[423] <= 1'b0;
    end else if(N1427) begin
      mem_q[423] <= mem_n[423];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[422] <= 1'b0;
    end else if(N1427) begin
      mem_q[422] <= mem_n[422];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[421] <= 1'b0;
    end else if(N1427) begin
      mem_q[421] <= mem_n[421];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[420] <= 1'b0;
    end else if(N1427) begin
      mem_q[420] <= mem_n[420];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[419] <= 1'b0;
    end else if(N1427) begin
      mem_q[419] <= mem_n[419];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[418] <= 1'b0;
    end else if(N1427) begin
      mem_q[418] <= mem_n[418];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[417] <= 1'b0;
    end else if(N1427) begin
      mem_q[417] <= mem_n[417];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[416] <= 1'b0;
    end else if(N1427) begin
      mem_q[416] <= mem_n[416];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[415] <= 1'b0;
    end else if(N1427) begin
      mem_q[415] <= mem_n[415];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[414] <= 1'b0;
    end else if(N1427) begin
      mem_q[414] <= mem_n[414];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[413] <= 1'b0;
    end else if(N1427) begin
      mem_q[413] <= mem_n[413];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[412] <= 1'b0;
    end else if(N1427) begin
      mem_q[412] <= mem_n[412];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[411] <= 1'b0;
    end else if(N1427) begin
      mem_q[411] <= mem_n[411];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[410] <= 1'b0;
    end else if(N1427) begin
      mem_q[410] <= mem_n[410];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[409] <= 1'b0;
    end else if(N1427) begin
      mem_q[409] <= mem_n[409];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[408] <= 1'b0;
    end else if(N1427) begin
      mem_q[408] <= mem_n[408];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[407] <= 1'b0;
    end else if(N1427) begin
      mem_q[407] <= mem_n[407];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[406] <= 1'b0;
    end else if(N1427) begin
      mem_q[406] <= mem_n[406];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[405] <= 1'b0;
    end else if(N1427) begin
      mem_q[405] <= mem_n[405];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[404] <= 1'b0;
    end else if(N1427) begin
      mem_q[404] <= mem_n[404];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[403] <= 1'b0;
    end else if(N1427) begin
      mem_q[403] <= mem_n[403];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[402] <= 1'b0;
    end else if(N1427) begin
      mem_q[402] <= mem_n[402];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[401] <= 1'b0;
    end else if(N1427) begin
      mem_q[401] <= mem_n[401];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[400] <= 1'b0;
    end else if(N1427) begin
      mem_q[400] <= mem_n[400];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[399] <= 1'b0;
    end else if(N1427) begin
      mem_q[399] <= mem_n[399];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[398] <= 1'b0;
    end else if(N1427) begin
      mem_q[398] <= mem_n[398];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[397] <= 1'b0;
    end else if(N1427) begin
      mem_q[397] <= mem_n[397];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[396] <= 1'b0;
    end else if(N1427) begin
      mem_q[396] <= mem_n[396];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[395] <= 1'b0;
    end else if(N1427) begin
      mem_q[395] <= mem_n[395];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[394] <= 1'b0;
    end else if(N1427) begin
      mem_q[394] <= mem_n[394];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[393] <= 1'b0;
    end else if(N1427) begin
      mem_q[393] <= mem_n[393];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[392] <= 1'b0;
    end else if(N1427) begin
      mem_q[392] <= mem_n[392];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[391] <= 1'b0;
    end else if(N1427) begin
      mem_q[391] <= mem_n[391];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[390] <= 1'b0;
    end else if(N1427) begin
      mem_q[390] <= mem_n[390];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[389] <= 1'b0;
    end else if(N1427) begin
      mem_q[389] <= mem_n[389];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[388] <= 1'b0;
    end else if(N1427) begin
      mem_q[388] <= mem_n[388];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[387] <= 1'b0;
    end else if(N1427) begin
      mem_q[387] <= mem_n[387];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[386] <= 1'b0;
    end else if(N1427) begin
      mem_q[386] <= mem_n[386];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[385] <= 1'b0;
    end else if(N1427) begin
      mem_q[385] <= mem_n[385];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[384] <= 1'b0;
    end else if(N1427) begin
      mem_q[384] <= mem_n[384];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[383] <= 1'b0;
    end else if(N1427) begin
      mem_q[383] <= mem_n[383];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[382] <= 1'b0;
    end else if(N1427) begin
      mem_q[382] <= mem_n[382];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[381] <= 1'b0;
    end else if(N1427) begin
      mem_q[381] <= mem_n[381];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[380] <= 1'b0;
    end else if(N1427) begin
      mem_q[380] <= mem_n[380];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[379] <= 1'b0;
    end else if(N1427) begin
      mem_q[379] <= mem_n[379];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[378] <= 1'b0;
    end else if(N1427) begin
      mem_q[378] <= mem_n[378];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[377] <= 1'b0;
    end else if(N1427) begin
      mem_q[377] <= mem_n[377];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[376] <= 1'b0;
    end else if(N1427) begin
      mem_q[376] <= mem_n[376];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[375] <= 1'b0;
    end else if(N1427) begin
      mem_q[375] <= mem_n[375];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[374] <= 1'b0;
    end else if(N1427) begin
      mem_q[374] <= mem_n[374];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[373] <= 1'b0;
    end else if(N1427) begin
      mem_q[373] <= mem_n[373];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[372] <= 1'b0;
    end else if(N1427) begin
      mem_q[372] <= mem_n[372];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[371] <= 1'b0;
    end else if(N1427) begin
      mem_q[371] <= mem_n[371];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[370] <= 1'b0;
    end else if(N1427) begin
      mem_q[370] <= mem_n[370];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[369] <= 1'b0;
    end else if(N1427) begin
      mem_q[369] <= mem_n[369];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[368] <= 1'b0;
    end else if(N1427) begin
      mem_q[368] <= mem_n[368];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[367] <= 1'b0;
    end else if(N1427) begin
      mem_q[367] <= mem_n[367];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[366] <= 1'b0;
    end else if(N1427) begin
      mem_q[366] <= mem_n[366];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[365] <= 1'b0;
    end else if(N1427) begin
      mem_q[365] <= mem_n[365];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[364] <= 1'b0;
    end else if(N1427) begin
      mem_q[364] <= mem_n[364];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[363] <= 1'b0;
    end else if(N1427) begin
      mem_q[363] <= mem_n[363];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[362] <= 1'b0;
    end else if(N1427) begin
      mem_q[362] <= mem_n[362];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[361] <= 1'b0;
    end else if(N1427) begin
      mem_q[361] <= mem_n[361];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[360] <= 1'b0;
    end else if(N1427) begin
      mem_q[360] <= mem_n[360];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[359] <= 1'b0;
    end else if(N1427) begin
      mem_q[359] <= mem_n[359];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[358] <= 1'b0;
    end else if(N1427) begin
      mem_q[358] <= mem_n[358];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[357] <= 1'b0;
    end else if(N1427) begin
      mem_q[357] <= mem_n[357];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[356] <= 1'b0;
    end else if(N1427) begin
      mem_q[356] <= mem_n[356];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[355] <= 1'b0;
    end else if(N1427) begin
      mem_q[355] <= mem_n[355];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[354] <= 1'b0;
    end else if(N1427) begin
      mem_q[354] <= mem_n[354];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[353] <= 1'b0;
    end else if(N1427) begin
      mem_q[353] <= mem_n[353];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[352] <= 1'b0;
    end else if(N1427) begin
      mem_q[352] <= mem_n[352];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[351] <= 1'b0;
    end else if(N1427) begin
      mem_q[351] <= mem_n[351];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[350] <= 1'b0;
    end else if(N1427) begin
      mem_q[350] <= mem_n[350];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[349] <= 1'b0;
    end else if(N1427) begin
      mem_q[349] <= mem_n[349];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[348] <= 1'b0;
    end else if(N1427) begin
      mem_q[348] <= mem_n[348];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[347] <= 1'b0;
    end else if(N1427) begin
      mem_q[347] <= mem_n[347];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[346] <= 1'b0;
    end else if(N1427) begin
      mem_q[346] <= mem_n[346];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[345] <= 1'b0;
    end else if(N1427) begin
      mem_q[345] <= mem_n[345];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[344] <= 1'b0;
    end else if(N1427) begin
      mem_q[344] <= mem_n[344];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[343] <= 1'b0;
    end else if(N1427) begin
      mem_q[343] <= mem_n[343];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[342] <= 1'b0;
    end else if(N1427) begin
      mem_q[342] <= mem_n[342];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[341] <= 1'b0;
    end else if(N1427) begin
      mem_q[341] <= mem_n[341];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[340] <= 1'b0;
    end else if(N1427) begin
      mem_q[340] <= mem_n[340];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[339] <= 1'b0;
    end else if(N1427) begin
      mem_q[339] <= mem_n[339];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[338] <= 1'b0;
    end else if(N1427) begin
      mem_q[338] <= mem_n[338];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[337] <= 1'b0;
    end else if(N1427) begin
      mem_q[337] <= mem_n[337];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[336] <= 1'b0;
    end else if(N1427) begin
      mem_q[336] <= mem_n[336];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[335] <= 1'b0;
    end else if(N1427) begin
      mem_q[335] <= mem_n[335];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[334] <= 1'b0;
    end else if(N1427) begin
      mem_q[334] <= mem_n[334];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[333] <= 1'b0;
    end else if(N1427) begin
      mem_q[333] <= mem_n[333];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[332] <= 1'b0;
    end else if(N1427) begin
      mem_q[332] <= mem_n[332];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[331] <= 1'b0;
    end else if(N1427) begin
      mem_q[331] <= mem_n[331];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[330] <= 1'b0;
    end else if(N1427) begin
      mem_q[330] <= mem_n[330];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[329] <= 1'b0;
    end else if(N1427) begin
      mem_q[329] <= mem_n[329];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[328] <= 1'b0;
    end else if(N1427) begin
      mem_q[328] <= mem_n[328];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[327] <= 1'b0;
    end else if(N1427) begin
      mem_q[327] <= mem_n[327];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[326] <= 1'b0;
    end else if(N1427) begin
      mem_q[326] <= mem_n[326];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[325] <= 1'b0;
    end else if(N1427) begin
      mem_q[325] <= mem_n[325];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[324] <= 1'b0;
    end else if(N1427) begin
      mem_q[324] <= mem_n[324];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[323] <= 1'b0;
    end else if(N1427) begin
      mem_q[323] <= mem_n[323];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[322] <= 1'b0;
    end else if(N1427) begin
      mem_q[322] <= mem_n[322];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[321] <= 1'b0;
    end else if(N1427) begin
      mem_q[321] <= mem_n[321];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[320] <= 1'b0;
    end else if(N1427) begin
      mem_q[320] <= mem_n[320];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[319] <= 1'b0;
    end else if(N1427) begin
      mem_q[319] <= mem_n[319];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[318] <= 1'b0;
    end else if(N1427) begin
      mem_q[318] <= mem_n[318];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[317] <= 1'b0;
    end else if(N1427) begin
      mem_q[317] <= mem_n[317];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[316] <= 1'b0;
    end else if(N1427) begin
      mem_q[316] <= mem_n[316];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[315] <= 1'b0;
    end else if(N1427) begin
      mem_q[315] <= mem_n[315];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[314] <= 1'b0;
    end else if(N1427) begin
      mem_q[314] <= mem_n[314];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[313] <= 1'b0;
    end else if(N1427) begin
      mem_q[313] <= mem_n[313];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[312] <= 1'b0;
    end else if(N1427) begin
      mem_q[312] <= mem_n[312];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[311] <= 1'b0;
    end else if(N1427) begin
      mem_q[311] <= mem_n[311];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[310] <= 1'b0;
    end else if(N1427) begin
      mem_q[310] <= mem_n[310];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[309] <= 1'b0;
    end else if(N1427) begin
      mem_q[309] <= mem_n[309];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[308] <= 1'b0;
    end else if(N1427) begin
      mem_q[308] <= mem_n[308];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[307] <= 1'b0;
    end else if(N1427) begin
      mem_q[307] <= mem_n[307];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[306] <= 1'b0;
    end else if(N1427) begin
      mem_q[306] <= mem_n[306];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[305] <= 1'b0;
    end else if(N1427) begin
      mem_q[305] <= mem_n[305];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[304] <= 1'b0;
    end else if(N1427) begin
      mem_q[304] <= mem_n[304];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[303] <= 1'b0;
    end else if(N1427) begin
      mem_q[303] <= mem_n[303];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[302] <= 1'b0;
    end else if(N1427) begin
      mem_q[302] <= mem_n[302];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[301] <= 1'b0;
    end else if(N1427) begin
      mem_q[301] <= mem_n[301];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[300] <= 1'b0;
    end else if(N1427) begin
      mem_q[300] <= mem_n[300];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[299] <= 1'b0;
    end else if(N1427) begin
      mem_q[299] <= mem_n[299];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[298] <= 1'b0;
    end else if(N1427) begin
      mem_q[298] <= mem_n[298];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[297] <= 1'b0;
    end else if(N1427) begin
      mem_q[297] <= mem_n[297];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[296] <= 1'b0;
    end else if(N1427) begin
      mem_q[296] <= mem_n[296];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[295] <= 1'b0;
    end else if(N1427) begin
      mem_q[295] <= mem_n[295];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[294] <= 1'b0;
    end else if(N1427) begin
      mem_q[294] <= mem_n[294];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[293] <= 1'b0;
    end else if(N1427) begin
      mem_q[293] <= mem_n[293];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[292] <= 1'b0;
    end else if(N1427) begin
      mem_q[292] <= mem_n[292];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[291] <= 1'b0;
    end else if(N1427) begin
      mem_q[291] <= mem_n[291];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[290] <= 1'b0;
    end else if(N1427) begin
      mem_q[290] <= mem_n[290];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[289] <= 1'b0;
    end else if(N1427) begin
      mem_q[289] <= mem_n[289];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[288] <= 1'b0;
    end else if(N1427) begin
      mem_q[288] <= mem_n[288];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[287] <= 1'b0;
    end else if(N1427) begin
      mem_q[287] <= mem_n[287];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[286] <= 1'b0;
    end else if(N1427) begin
      mem_q[286] <= mem_n[286];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[285] <= 1'b0;
    end else if(N1427) begin
      mem_q[285] <= mem_n[285];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[284] <= 1'b0;
    end else if(N1427) begin
      mem_q[284] <= mem_n[284];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[283] <= 1'b0;
    end else if(N1427) begin
      mem_q[283] <= mem_n[283];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[282] <= 1'b0;
    end else if(N1427) begin
      mem_q[282] <= mem_n[282];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[281] <= 1'b0;
    end else if(N1427) begin
      mem_q[281] <= mem_n[281];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[280] <= 1'b0;
    end else if(N1427) begin
      mem_q[280] <= mem_n[280];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[279] <= 1'b0;
    end else if(N1427) begin
      mem_q[279] <= mem_n[279];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[278] <= 1'b0;
    end else if(N1427) begin
      mem_q[278] <= mem_n[278];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[277] <= 1'b0;
    end else if(N1427) begin
      mem_q[277] <= mem_n[277];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[276] <= 1'b0;
    end else if(N1427) begin
      mem_q[276] <= mem_n[276];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[275] <= 1'b0;
    end else if(N1427) begin
      mem_q[275] <= mem_n[275];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[274] <= 1'b0;
    end else if(N1427) begin
      mem_q[274] <= mem_n[274];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[273] <= 1'b0;
    end else if(N1427) begin
      mem_q[273] <= mem_n[273];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[272] <= 1'b0;
    end else if(N1427) begin
      mem_q[272] <= mem_n[272];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[271] <= 1'b0;
    end else if(N1427) begin
      mem_q[271] <= mem_n[271];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[270] <= 1'b0;
    end else if(N1427) begin
      mem_q[270] <= mem_n[270];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[269] <= 1'b0;
    end else if(N1427) begin
      mem_q[269] <= mem_n[269];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[268] <= 1'b0;
    end else if(N1427) begin
      mem_q[268] <= mem_n[268];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[267] <= 1'b0;
    end else if(N1427) begin
      mem_q[267] <= mem_n[267];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[266] <= 1'b0;
    end else if(N1427) begin
      mem_q[266] <= mem_n[266];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[265] <= 1'b0;
    end else if(N1427) begin
      mem_q[265] <= mem_n[265];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[264] <= 1'b0;
    end else if(N1427) begin
      mem_q[264] <= mem_n[264];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[263] <= 1'b0;
    end else if(N1427) begin
      mem_q[263] <= mem_n[263];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[262] <= 1'b0;
    end else if(N1427) begin
      mem_q[262] <= mem_n[262];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[261] <= 1'b0;
    end else if(N1427) begin
      mem_q[261] <= mem_n[261];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[260] <= 1'b0;
    end else if(N1427) begin
      mem_q[260] <= mem_n[260];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[259] <= 1'b0;
    end else if(N1427) begin
      mem_q[259] <= mem_n[259];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[258] <= 1'b0;
    end else if(N1427) begin
      mem_q[258] <= mem_n[258];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[257] <= 1'b0;
    end else if(N1427) begin
      mem_q[257] <= mem_n[257];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[256] <= 1'b0;
    end else if(N1427) begin
      mem_q[256] <= mem_n[256];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[255] <= 1'b0;
    end else if(N1427) begin
      mem_q[255] <= mem_n[255];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[254] <= 1'b0;
    end else if(N1427) begin
      mem_q[254] <= mem_n[254];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[253] <= 1'b0;
    end else if(N1427) begin
      mem_q[253] <= mem_n[253];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[252] <= 1'b0;
    end else if(N1427) begin
      mem_q[252] <= mem_n[252];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[251] <= 1'b0;
    end else if(N1427) begin
      mem_q[251] <= mem_n[251];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[250] <= 1'b0;
    end else if(N1427) begin
      mem_q[250] <= mem_n[250];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[249] <= 1'b0;
    end else if(N1427) begin
      mem_q[249] <= mem_n[249];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[248] <= 1'b0;
    end else if(N1427) begin
      mem_q[248] <= mem_n[248];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[247] <= 1'b0;
    end else if(N1427) begin
      mem_q[247] <= mem_n[247];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[246] <= 1'b0;
    end else if(N1427) begin
      mem_q[246] <= mem_n[246];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[245] <= 1'b0;
    end else if(N1427) begin
      mem_q[245] <= mem_n[245];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[244] <= 1'b0;
    end else if(N1427) begin
      mem_q[244] <= mem_n[244];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[243] <= 1'b0;
    end else if(N1427) begin
      mem_q[243] <= mem_n[243];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[242] <= 1'b0;
    end else if(N1427) begin
      mem_q[242] <= mem_n[242];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[241] <= 1'b0;
    end else if(N1427) begin
      mem_q[241] <= mem_n[241];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[240] <= 1'b0;
    end else if(N1427) begin
      mem_q[240] <= mem_n[240];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[239] <= 1'b0;
    end else if(N1427) begin
      mem_q[239] <= mem_n[239];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[238] <= 1'b0;
    end else if(N1427) begin
      mem_q[238] <= mem_n[238];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[237] <= 1'b0;
    end else if(N1427) begin
      mem_q[237] <= mem_n[237];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[236] <= 1'b0;
    end else if(N1427) begin
      mem_q[236] <= mem_n[236];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[235] <= 1'b0;
    end else if(N1427) begin
      mem_q[235] <= mem_n[235];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[234] <= 1'b0;
    end else if(N1427) begin
      mem_q[234] <= mem_n[234];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[233] <= 1'b0;
    end else if(N1427) begin
      mem_q[233] <= mem_n[233];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[232] <= 1'b0;
    end else if(N1427) begin
      mem_q[232] <= mem_n[232];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[231] <= 1'b0;
    end else if(N1427) begin
      mem_q[231] <= mem_n[231];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[230] <= 1'b0;
    end else if(N1427) begin
      mem_q[230] <= mem_n[230];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[229] <= 1'b0;
    end else if(N1427) begin
      mem_q[229] <= mem_n[229];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[228] <= 1'b0;
    end else if(N1427) begin
      mem_q[228] <= mem_n[228];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[227] <= 1'b0;
    end else if(N1427) begin
      mem_q[227] <= mem_n[227];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[226] <= 1'b0;
    end else if(N1427) begin
      mem_q[226] <= mem_n[226];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[225] <= 1'b0;
    end else if(N1427) begin
      mem_q[225] <= mem_n[225];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[224] <= 1'b0;
    end else if(N1427) begin
      mem_q[224] <= mem_n[224];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[223] <= 1'b0;
    end else if(N1427) begin
      mem_q[223] <= mem_n[223];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[222] <= 1'b0;
    end else if(N1427) begin
      mem_q[222] <= mem_n[222];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[221] <= 1'b0;
    end else if(N1427) begin
      mem_q[221] <= mem_n[221];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[220] <= 1'b0;
    end else if(N1427) begin
      mem_q[220] <= mem_n[220];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[219] <= 1'b0;
    end else if(N1427) begin
      mem_q[219] <= mem_n[219];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[218] <= 1'b0;
    end else if(N1427) begin
      mem_q[218] <= mem_n[218];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[217] <= 1'b0;
    end else if(N1427) begin
      mem_q[217] <= mem_n[217];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[216] <= 1'b0;
    end else if(N1427) begin
      mem_q[216] <= mem_n[216];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[215] <= 1'b0;
    end else if(N1427) begin
      mem_q[215] <= mem_n[215];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[214] <= 1'b0;
    end else if(N1427) begin
      mem_q[214] <= mem_n[214];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[213] <= 1'b0;
    end else if(N1427) begin
      mem_q[213] <= mem_n[213];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[212] <= 1'b0;
    end else if(N1427) begin
      mem_q[212] <= mem_n[212];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[211] <= 1'b0;
    end else if(N1427) begin
      mem_q[211] <= mem_n[211];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[210] <= 1'b0;
    end else if(N1427) begin
      mem_q[210] <= mem_n[210];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[209] <= 1'b0;
    end else if(N1427) begin
      mem_q[209] <= mem_n[209];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[208] <= 1'b0;
    end else if(N1427) begin
      mem_q[208] <= mem_n[208];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[207] <= 1'b0;
    end else if(N1427) begin
      mem_q[207] <= mem_n[207];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[206] <= 1'b0;
    end else if(N1427) begin
      mem_q[206] <= mem_n[206];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[205] <= 1'b0;
    end else if(N1427) begin
      mem_q[205] <= mem_n[205];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[204] <= 1'b0;
    end else if(N1427) begin
      mem_q[204] <= mem_n[204];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[203] <= 1'b0;
    end else if(N1427) begin
      mem_q[203] <= mem_n[203];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[202] <= 1'b0;
    end else if(N1427) begin
      mem_q[202] <= mem_n[202];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[201] <= 1'b0;
    end else if(N1427) begin
      mem_q[201] <= mem_n[201];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[200] <= 1'b0;
    end else if(N1427) begin
      mem_q[200] <= mem_n[200];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[199] <= 1'b0;
    end else if(N1427) begin
      mem_q[199] <= mem_n[199];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[198] <= 1'b0;
    end else if(N1427) begin
      mem_q[198] <= mem_n[198];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[197] <= 1'b0;
    end else if(N1427) begin
      mem_q[197] <= mem_n[197];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[196] <= 1'b0;
    end else if(N1427) begin
      mem_q[196] <= mem_n[196];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[195] <= 1'b0;
    end else if(N1427) begin
      mem_q[195] <= mem_n[195];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[194] <= 1'b0;
    end else if(N1427) begin
      mem_q[194] <= mem_n[194];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[193] <= 1'b0;
    end else if(N1427) begin
      mem_q[193] <= mem_n[193];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[192] <= 1'b0;
    end else if(N1427) begin
      mem_q[192] <= mem_n[192];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[191] <= 1'b0;
    end else if(N1427) begin
      mem_q[191] <= mem_n[191];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[190] <= 1'b0;
    end else if(N1427) begin
      mem_q[190] <= mem_n[190];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[189] <= 1'b0;
    end else if(N1427) begin
      mem_q[189] <= mem_n[189];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[188] <= 1'b0;
    end else if(N1427) begin
      mem_q[188] <= mem_n[188];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[187] <= 1'b0;
    end else if(N1427) begin
      mem_q[187] <= mem_n[187];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[186] <= 1'b0;
    end else if(N1427) begin
      mem_q[186] <= mem_n[186];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[185] <= 1'b0;
    end else if(N1427) begin
      mem_q[185] <= mem_n[185];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[184] <= 1'b0;
    end else if(N1427) begin
      mem_q[184] <= mem_n[184];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[183] <= 1'b0;
    end else if(N1427) begin
      mem_q[183] <= mem_n[183];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[182] <= 1'b0;
    end else if(N1427) begin
      mem_q[182] <= mem_n[182];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[181] <= 1'b0;
    end else if(N1427) begin
      mem_q[181] <= mem_n[181];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[180] <= 1'b0;
    end else if(N1427) begin
      mem_q[180] <= mem_n[180];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[179] <= 1'b0;
    end else if(N1427) begin
      mem_q[179] <= mem_n[179];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[178] <= 1'b0;
    end else if(N1427) begin
      mem_q[178] <= mem_n[178];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[177] <= 1'b0;
    end else if(N1427) begin
      mem_q[177] <= mem_n[177];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[176] <= 1'b0;
    end else if(N1427) begin
      mem_q[176] <= mem_n[176];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[175] <= 1'b0;
    end else if(N1427) begin
      mem_q[175] <= mem_n[175];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[174] <= 1'b0;
    end else if(N1427) begin
      mem_q[174] <= mem_n[174];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[173] <= 1'b0;
    end else if(N1427) begin
      mem_q[173] <= mem_n[173];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[172] <= 1'b0;
    end else if(N1427) begin
      mem_q[172] <= mem_n[172];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[171] <= 1'b0;
    end else if(N1427) begin
      mem_q[171] <= mem_n[171];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[170] <= 1'b0;
    end else if(N1427) begin
      mem_q[170] <= mem_n[170];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[169] <= 1'b0;
    end else if(N1427) begin
      mem_q[169] <= mem_n[169];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[168] <= 1'b0;
    end else if(N1427) begin
      mem_q[168] <= mem_n[168];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[167] <= 1'b0;
    end else if(N1427) begin
      mem_q[167] <= mem_n[167];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[166] <= 1'b0;
    end else if(N1427) begin
      mem_q[166] <= mem_n[166];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[165] <= 1'b0;
    end else if(N1427) begin
      mem_q[165] <= mem_n[165];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[164] <= 1'b0;
    end else if(N1427) begin
      mem_q[164] <= mem_n[164];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[163] <= 1'b0;
    end else if(N1427) begin
      mem_q[163] <= mem_n[163];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[162] <= 1'b0;
    end else if(N1427) begin
      mem_q[162] <= mem_n[162];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[161] <= 1'b0;
    end else if(N1427) begin
      mem_q[161] <= mem_n[161];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[160] <= 1'b0;
    end else if(N1427) begin
      mem_q[160] <= mem_n[160];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[159] <= 1'b0;
    end else if(N1427) begin
      mem_q[159] <= mem_n[159];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[158] <= 1'b0;
    end else if(N1427) begin
      mem_q[158] <= mem_n[158];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[157] <= 1'b0;
    end else if(N1427) begin
      mem_q[157] <= mem_n[157];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[156] <= 1'b0;
    end else if(N1427) begin
      mem_q[156] <= mem_n[156];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[155] <= 1'b0;
    end else if(N1427) begin
      mem_q[155] <= mem_n[155];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[154] <= 1'b0;
    end else if(N1427) begin
      mem_q[154] <= mem_n[154];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[153] <= 1'b0;
    end else if(N1427) begin
      mem_q[153] <= mem_n[153];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[152] <= 1'b0;
    end else if(N1427) begin
      mem_q[152] <= mem_n[152];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[151] <= 1'b0;
    end else if(N1427) begin
      mem_q[151] <= mem_n[151];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[150] <= 1'b0;
    end else if(N1427) begin
      mem_q[150] <= mem_n[150];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[149] <= 1'b0;
    end else if(N1427) begin
      mem_q[149] <= mem_n[149];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[148] <= 1'b0;
    end else if(N1427) begin
      mem_q[148] <= mem_n[148];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[147] <= 1'b0;
    end else if(N1427) begin
      mem_q[147] <= mem_n[147];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[146] <= 1'b0;
    end else if(N1427) begin
      mem_q[146] <= mem_n[146];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[145] <= 1'b0;
    end else if(N1427) begin
      mem_q[145] <= mem_n[145];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[144] <= 1'b0;
    end else if(N1427) begin
      mem_q[144] <= mem_n[144];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[143] <= 1'b0;
    end else if(N1427) begin
      mem_q[143] <= mem_n[143];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[142] <= 1'b0;
    end else if(N1427) begin
      mem_q[142] <= mem_n[142];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[141] <= 1'b0;
    end else if(N1427) begin
      mem_q[141] <= mem_n[141];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[140] <= 1'b0;
    end else if(N1427) begin
      mem_q[140] <= mem_n[140];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[139] <= 1'b0;
    end else if(N1427) begin
      mem_q[139] <= mem_n[139];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[138] <= 1'b0;
    end else if(N1427) begin
      mem_q[138] <= mem_n[138];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[137] <= 1'b0;
    end else if(N1427) begin
      mem_q[137] <= mem_n[137];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[136] <= 1'b0;
    end else if(N1427) begin
      mem_q[136] <= mem_n[136];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[135] <= 1'b0;
    end else if(N1427) begin
      mem_q[135] <= mem_n[135];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[134] <= 1'b0;
    end else if(N1427) begin
      mem_q[134] <= mem_n[134];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[133] <= 1'b0;
    end else if(N1427) begin
      mem_q[133] <= mem_n[133];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[132] <= 1'b0;
    end else if(N1427) begin
      mem_q[132] <= mem_n[132];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[131] <= 1'b0;
    end else if(N1427) begin
      mem_q[131] <= mem_n[131];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[130] <= 1'b0;
    end else if(N1427) begin
      mem_q[130] <= mem_n[130];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[129] <= 1'b0;
    end else if(N1427) begin
      mem_q[129] <= mem_n[129];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[128] <= 1'b0;
    end else if(N1427) begin
      mem_q[128] <= mem_n[128];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[127] <= 1'b0;
    end else if(N1427) begin
      mem_q[127] <= mem_n[127];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[126] <= 1'b0;
    end else if(N1427) begin
      mem_q[126] <= mem_n[126];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[125] <= 1'b0;
    end else if(N1427) begin
      mem_q[125] <= mem_n[125];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[124] <= 1'b0;
    end else if(N1427) begin
      mem_q[124] <= mem_n[124];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[123] <= 1'b0;
    end else if(N1427) begin
      mem_q[123] <= mem_n[123];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[122] <= 1'b0;
    end else if(N1427) begin
      mem_q[122] <= mem_n[122];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[121] <= 1'b0;
    end else if(N1427) begin
      mem_q[121] <= mem_n[121];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[120] <= 1'b0;
    end else if(N1427) begin
      mem_q[120] <= mem_n[120];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[119] <= 1'b0;
    end else if(N1427) begin
      mem_q[119] <= mem_n[119];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[118] <= 1'b0;
    end else if(N1427) begin
      mem_q[118] <= mem_n[118];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[117] <= 1'b0;
    end else if(N1427) begin
      mem_q[117] <= mem_n[117];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[116] <= 1'b0;
    end else if(N1427) begin
      mem_q[116] <= mem_n[116];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[115] <= 1'b0;
    end else if(N1427) begin
      mem_q[115] <= mem_n[115];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[114] <= 1'b0;
    end else if(N1427) begin
      mem_q[114] <= mem_n[114];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[113] <= 1'b0;
    end else if(N1427) begin
      mem_q[113] <= mem_n[113];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[112] <= 1'b0;
    end else if(N1427) begin
      mem_q[112] <= mem_n[112];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[111] <= 1'b0;
    end else if(N1427) begin
      mem_q[111] <= mem_n[111];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[110] <= 1'b0;
    end else if(N1427) begin
      mem_q[110] <= mem_n[110];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[109] <= 1'b0;
    end else if(N1427) begin
      mem_q[109] <= mem_n[109];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[108] <= 1'b0;
    end else if(N1427) begin
      mem_q[108] <= mem_n[108];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[107] <= 1'b0;
    end else if(N1427) begin
      mem_q[107] <= mem_n[107];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[106] <= 1'b0;
    end else if(N1427) begin
      mem_q[106] <= mem_n[106];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[105] <= 1'b0;
    end else if(N1427) begin
      mem_q[105] <= mem_n[105];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[104] <= 1'b0;
    end else if(N1427) begin
      mem_q[104] <= mem_n[104];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[103] <= 1'b0;
    end else if(N1427) begin
      mem_q[103] <= mem_n[103];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[102] <= 1'b0;
    end else if(N1427) begin
      mem_q[102] <= mem_n[102];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[101] <= 1'b0;
    end else if(N1427) begin
      mem_q[101] <= mem_n[101];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[100] <= 1'b0;
    end else if(N1427) begin
      mem_q[100] <= mem_n[100];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[99] <= 1'b0;
    end else if(N1427) begin
      mem_q[99] <= mem_n[99];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[98] <= 1'b0;
    end else if(N1427) begin
      mem_q[98] <= mem_n[98];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[97] <= 1'b0;
    end else if(N1427) begin
      mem_q[97] <= mem_n[97];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[96] <= 1'b0;
    end else if(N1427) begin
      mem_q[96] <= mem_n[96];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[95] <= 1'b0;
    end else if(N1427) begin
      mem_q[95] <= mem_n[95];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[94] <= 1'b0;
    end else if(N1427) begin
      mem_q[94] <= mem_n[94];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[93] <= 1'b0;
    end else if(N1427) begin
      mem_q[93] <= mem_n[93];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[92] <= 1'b0;
    end else if(N1427) begin
      mem_q[92] <= mem_n[92];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[91] <= 1'b0;
    end else if(N1427) begin
      mem_q[91] <= mem_n[91];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[90] <= 1'b0;
    end else if(N1427) begin
      mem_q[90] <= mem_n[90];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[89] <= 1'b0;
    end else if(N1427) begin
      mem_q[89] <= mem_n[89];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[88] <= 1'b0;
    end else if(N1427) begin
      mem_q[88] <= mem_n[88];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[87] <= 1'b0;
    end else if(N1427) begin
      mem_q[87] <= mem_n[87];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[86] <= 1'b0;
    end else if(N1427) begin
      mem_q[86] <= mem_n[86];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[85] <= 1'b0;
    end else if(N1427) begin
      mem_q[85] <= mem_n[85];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[84] <= 1'b0;
    end else if(N1427) begin
      mem_q[84] <= mem_n[84];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[83] <= 1'b0;
    end else if(N1427) begin
      mem_q[83] <= mem_n[83];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[82] <= 1'b0;
    end else if(N1427) begin
      mem_q[82] <= mem_n[82];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[81] <= 1'b0;
    end else if(N1427) begin
      mem_q[81] <= mem_n[81];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[80] <= 1'b0;
    end else if(N1427) begin
      mem_q[80] <= mem_n[80];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[79] <= 1'b0;
    end else if(N1427) begin
      mem_q[79] <= mem_n[79];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[78] <= 1'b0;
    end else if(N1427) begin
      mem_q[78] <= mem_n[78];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[77] <= 1'b0;
    end else if(N1427) begin
      mem_q[77] <= mem_n[77];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[76] <= 1'b0;
    end else if(N1427) begin
      mem_q[76] <= mem_n[76];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[75] <= 1'b0;
    end else if(N1427) begin
      mem_q[75] <= mem_n[75];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[74] <= 1'b0;
    end else if(N1427) begin
      mem_q[74] <= mem_n[74];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[73] <= 1'b0;
    end else if(N1427) begin
      mem_q[73] <= mem_n[73];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[72] <= 1'b0;
    end else if(N1427) begin
      mem_q[72] <= mem_n[72];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[71] <= 1'b0;
    end else if(N1427) begin
      mem_q[71] <= mem_n[71];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[70] <= 1'b0;
    end else if(N1427) begin
      mem_q[70] <= mem_n[70];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[69] <= 1'b0;
    end else if(N1427) begin
      mem_q[69] <= mem_n[69];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[68] <= 1'b0;
    end else if(N1427) begin
      mem_q[68] <= mem_n[68];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[67] <= 1'b0;
    end else if(N1427) begin
      mem_q[67] <= mem_n[67];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[66] <= 1'b0;
    end else if(N1427) begin
      mem_q[66] <= mem_n[66];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[65] <= 1'b0;
    end else if(N1427) begin
      mem_q[65] <= mem_n[65];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[64] <= 1'b0;
    end else if(N1427) begin
      mem_q[64] <= mem_n[64];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[63] <= 1'b0;
    end else if(N1427) begin
      mem_q[63] <= mem_n[63];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[62] <= 1'b0;
    end else if(N1427) begin
      mem_q[62] <= mem_n[62];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[61] <= 1'b0;
    end else if(N1427) begin
      mem_q[61] <= mem_n[61];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[60] <= 1'b0;
    end else if(N1427) begin
      mem_q[60] <= mem_n[60];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[59] <= 1'b0;
    end else if(N1427) begin
      mem_q[59] <= mem_n[59];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[58] <= 1'b0;
    end else if(N1427) begin
      mem_q[58] <= mem_n[58];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[57] <= 1'b0;
    end else if(N1427) begin
      mem_q[57] <= mem_n[57];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[56] <= 1'b0;
    end else if(N1427) begin
      mem_q[56] <= mem_n[56];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[55] <= 1'b0;
    end else if(N1427) begin
      mem_q[55] <= mem_n[55];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[54] <= 1'b0;
    end else if(N1427) begin
      mem_q[54] <= mem_n[54];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[53] <= 1'b0;
    end else if(N1427) begin
      mem_q[53] <= mem_n[53];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[52] <= 1'b0;
    end else if(N1427) begin
      mem_q[52] <= mem_n[52];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[51] <= 1'b0;
    end else if(N1427) begin
      mem_q[51] <= mem_n[51];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[50] <= 1'b0;
    end else if(N1427) begin
      mem_q[50] <= mem_n[50];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[49] <= 1'b0;
    end else if(N1427) begin
      mem_q[49] <= mem_n[49];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[48] <= 1'b0;
    end else if(N1427) begin
      mem_q[48] <= mem_n[48];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[47] <= 1'b0;
    end else if(N1427) begin
      mem_q[47] <= mem_n[47];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[46] <= 1'b0;
    end else if(N1427) begin
      mem_q[46] <= mem_n[46];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[45] <= 1'b0;
    end else if(N1427) begin
      mem_q[45] <= mem_n[45];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[44] <= 1'b0;
    end else if(N1427) begin
      mem_q[44] <= mem_n[44];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[43] <= 1'b0;
    end else if(N1427) begin
      mem_q[43] <= mem_n[43];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[42] <= 1'b0;
    end else if(N1427) begin
      mem_q[42] <= mem_n[42];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[41] <= 1'b0;
    end else if(N1427) begin
      mem_q[41] <= mem_n[41];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[40] <= 1'b0;
    end else if(N1427) begin
      mem_q[40] <= mem_n[40];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[39] <= 1'b0;
    end else if(N1427) begin
      mem_q[39] <= mem_n[39];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[38] <= 1'b0;
    end else if(N1427) begin
      mem_q[38] <= mem_n[38];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[37] <= 1'b0;
    end else if(N1427) begin
      mem_q[37] <= mem_n[37];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[36] <= 1'b0;
    end else if(N1427) begin
      mem_q[36] <= mem_n[36];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[35] <= 1'b0;
    end else if(N1427) begin
      mem_q[35] <= mem_n[35];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[34] <= 1'b0;
    end else if(N1427) begin
      mem_q[34] <= mem_n[34];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[33] <= 1'b0;
    end else if(N1427) begin
      mem_q[33] <= mem_n[33];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[32] <= 1'b0;
    end else if(N1427) begin
      mem_q[32] <= mem_n[32];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[31] <= 1'b0;
    end else if(N1427) begin
      mem_q[31] <= mem_n[31];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[30] <= 1'b0;
    end else if(N1427) begin
      mem_q[30] <= mem_n[30];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[29] <= 1'b0;
    end else if(N1427) begin
      mem_q[29] <= mem_n[29];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[28] <= 1'b0;
    end else if(N1427) begin
      mem_q[28] <= mem_n[28];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[27] <= 1'b0;
    end else if(N1427) begin
      mem_q[27] <= mem_n[27];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[26] <= 1'b0;
    end else if(N1427) begin
      mem_q[26] <= mem_n[26];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[25] <= 1'b0;
    end else if(N1427) begin
      mem_q[25] <= mem_n[25];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[24] <= 1'b0;
    end else if(N1427) begin
      mem_q[24] <= mem_n[24];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[23] <= 1'b0;
    end else if(N1427) begin
      mem_q[23] <= mem_n[23];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[22] <= 1'b0;
    end else if(N1427) begin
      mem_q[22] <= mem_n[22];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[21] <= 1'b0;
    end else if(N1427) begin
      mem_q[21] <= mem_n[21];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[20] <= 1'b0;
    end else if(N1427) begin
      mem_q[20] <= mem_n[20];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[19] <= 1'b0;
    end else if(N1427) begin
      mem_q[19] <= mem_n[19];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[18] <= 1'b0;
    end else if(N1427) begin
      mem_q[18] <= mem_n[18];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[17] <= 1'b0;
    end else if(N1427) begin
      mem_q[17] <= mem_n[17];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[16] <= 1'b0;
    end else if(N1427) begin
      mem_q[16] <= mem_n[16];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[15] <= 1'b0;
    end else if(N1427) begin
      mem_q[15] <= mem_n[15];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[14] <= 1'b0;
    end else if(N1427) begin
      mem_q[14] <= mem_n[14];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[13] <= 1'b0;
    end else if(N1427) begin
      mem_q[13] <= mem_n[13];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[12] <= 1'b0;
    end else if(N1427) begin
      mem_q[12] <= mem_n[12];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[11] <= 1'b0;
    end else if(N1427) begin
      mem_q[11] <= mem_n[11];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[10] <= 1'b0;
    end else if(N1427) begin
      mem_q[10] <= mem_n[10];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[9] <= 1'b0;
    end else if(N1427) begin
      mem_q[9] <= mem_n[9];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[8] <= 1'b0;
    end else if(N1427) begin
      mem_q[8] <= mem_n[8];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[7] <= 1'b0;
    end else if(N1427) begin
      mem_q[7] <= mem_n[7];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[6] <= 1'b0;
    end else if(N1427) begin
      mem_q[6] <= mem_n[6];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[5] <= 1'b0;
    end else if(N1427) begin
      mem_q[5] <= mem_n[5];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[4] <= 1'b0;
    end else if(N1427) begin
      mem_q[4] <= mem_n[4];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[3] <= 1'b0;
    end else if(N1427) begin
      mem_q[3] <= mem_n[3];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[2] <= 1'b0;
    end else if(N1427) begin
      mem_q[2] <= mem_n[2];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[1] <= 1'b0;
    end else if(N1427) begin
      mem_q[1] <= mem_n[1];
    end 
  end


  always @(posedge clk_i or posedge N1415) begin
    if(N1415) begin
      mem_q[0] <= 1'b0;
    end else if(N1427) begin
      mem_q[0] <= mem_n[0];
    end 
  end

  assign N1438 = usage_o[2] | status_cnt_q[3];
  assign N1439 = usage_o[1] | N1438;
  assign N1440 = usage_o[0] | N1439;
  assign empty_o = ~N1440;
  assign N1442 = ~status_cnt_q[3];
  assign N1443 = usage_o[2] | N1442;
  assign N1444 = usage_o[1] | N1443;
  assign N1445 = usage_o[0] | N1444;
  assign full_o = ~N1445;
  assign { N1404, N1403, N1402 } = read_pointer_q + 1'b1;
  assign { N1408, N1407, N1406, N1405 } = { status_cnt_q[3:3], usage_o } - 1'b1;
  assign { N1395, N1394, N1393 } = write_pointer_q + 1'b1;
  assign { N1399, N1398, N1397, N1396 } = { status_cnt_q[3:3], usage_o } + 1'b1;
  assign N1447 = write_pointer_q[0] & write_pointer_q[1];
  assign N48 = N1447 & write_pointer_q[2];
  assign N1448 = N0 & write_pointer_q[1];
  assign N0 = ~write_pointer_q[0];
  assign N47 = N1448 & write_pointer_q[2];
  assign N1449 = write_pointer_q[0] & N1;
  assign N1 = ~write_pointer_q[1];
  assign N46 = N1449 & write_pointer_q[2];
  assign N1450 = N2 & N3;
  assign N2 = ~write_pointer_q[0];
  assign N3 = ~write_pointer_q[1];
  assign N45 = N1450 & write_pointer_q[2];
  assign N1451 = write_pointer_q[0] & write_pointer_q[1];
  assign N44 = N1451 & N4;
  assign N4 = ~write_pointer_q[2];
  assign N1452 = N5 & write_pointer_q[1];
  assign N5 = ~write_pointer_q[0];
  assign N43 = N1452 & N6;
  assign N6 = ~write_pointer_q[2];
  assign N1453 = write_pointer_q[0] & N7;
  assign N7 = ~write_pointer_q[1];
  assign N42 = N1453 & N8;
  assign N8 = ~write_pointer_q[2];
  assign N1454 = N9 & N10;
  assign N9 = ~write_pointer_q[0];
  assign N10 = ~write_pointer_q[1];
  assign N41 = N1454 & N11;
  assign N11 = ~write_pointer_q[2];
  assign { N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50 } = (N12)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N49)? { mem_q[0:0], mem_q[1:1], mem_q[2:2], mem_q[3:3], mem_q[4:4], mem_q[5:5], mem_q[6:6], mem_q[7:7], mem_q[8:8], mem_q[9:9], mem_q[10:10], mem_q[11:11], mem_q[12:12], mem_q[13:13], mem_q[14:14], mem_q[15:15], mem_q[16:16], mem_q[17:17], mem_q[18:18], mem_q[19:19], mem_q[20:20], mem_q[21:21], mem_q[22:22], mem_q[23:23], mem_q[24:24], mem_q[25:25], mem_q[26:26], mem_q[27:27], mem_q[28:28], mem_q[29:29], mem_q[30:30], mem_q[31:31], mem_q[32:32], mem_q[33:33], mem_q[34:34], mem_q[35:35], mem_q[36:36], mem_q[37:37], mem_q[38:38], mem_q[39:39], mem_q[40:40], mem_q[41:41], mem_q[42:42], mem_q[43:43], mem_q[44:44], mem_q[45:45], mem_q[46:46], mem_q[47:47], mem_q[48:48], mem_q[49:49], mem_q[50:50], mem_q[51:51], mem_q[52:52], mem_q[53:53], mem_q[54:54], mem_q[55:55], mem_q[56:56], mem_q[57:57], mem_q[58:58], mem_q[59:59], mem_q[60:60], mem_q[61:61], mem_q[62:62], mem_q[63:63], mem_q[64:64], mem_q[65:65], mem_q[66:66], mem_q[67:67], mem_q[68:68], mem_q[69:69], mem_q[70:70], mem_q[71:71], mem_q[72:72], mem_q[73:73], mem_q[74:74], mem_q[75:75], mem_q[76:76], mem_q[77:77], mem_q[78:78], mem_q[79:79], mem_q[80:80], mem_q[81:81], mem_q[82:82], mem_q[83:83], mem_q[84:84], mem_q[85:85], mem_q[86:86], mem_q[87:87], mem_q[88:88], mem_q[89:89], mem_q[90:90], mem_q[91:91], mem_q[92:92], mem_q[93:93], mem_q[94:94], mem_q[95:95], mem_q[96:96], mem_q[97:97], mem_q[98:98], mem_q[99:99], mem_q[100:100], mem_q[101:101], mem_q[102:102], mem_q[103:103], mem_q[104:104], mem_q[105:105], mem_q[106:106], mem_q[107:107], mem_q[108:108], mem_q[109:109], mem_q[110:110], mem_q[111:111], mem_q[112:112], mem_q[113:113], mem_q[114:114], mem_q[115:115], mem_q[116:116], mem_q[117:117], mem_q[118:118], mem_q[119:119], mem_q[120:120], mem_q[121:121], mem_q[122:122], mem_q[123:123], mem_q[124:124], mem_q[125:125], mem_q[126:126], mem_q[127:127], mem_q[128:128], mem_q[129:129], mem_q[130:130], mem_q[131:131], mem_q[132:132], mem_q[133:133], mem_q[134:134], mem_q[135:135], mem_q[136:136], mem_q[137:137], mem_q[138:138], mem_q[139:139], mem_q[140:140], mem_q[141:141], mem_q[142:142], mem_q[143:143], mem_q[144:144], mem_q[145:145], mem_q[146:146], mem_q[147:147], mem_q[148:148], mem_q[149:149], mem_q[150:150], mem_q[151:151], mem_q[152:152], mem_q[153:153], mem_q[154:154], mem_q[155:155], mem_q[156:156], mem_q[157:157], mem_q[158:158], mem_q[159:159], mem_q[160:160], mem_q[161:161], mem_q[162:162], mem_q[163:163], mem_q[164:164], mem_q[165:165], mem_q[166:166] } : 1'b0;
  assign N12 = N41;
  assign { N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218 } = (N13)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N217)? { mem_q[167:167], mem_q[168:168], mem_q[169:169], mem_q[170:170], mem_q[171:171], mem_q[172:172], mem_q[173:173], mem_q[174:174], mem_q[175:175], mem_q[176:176], mem_q[177:177], mem_q[178:178], mem_q[179:179], mem_q[180:180], mem_q[181:181], mem_q[182:182], mem_q[183:183], mem_q[184:184], mem_q[185:185], mem_q[186:186], mem_q[187:187], mem_q[188:188], mem_q[189:189], mem_q[190:190], mem_q[191:191], mem_q[192:192], mem_q[193:193], mem_q[194:194], mem_q[195:195], mem_q[196:196], mem_q[197:197], mem_q[198:198], mem_q[199:199], mem_q[200:200], mem_q[201:201], mem_q[202:202], mem_q[203:203], mem_q[204:204], mem_q[205:205], mem_q[206:206], mem_q[207:207], mem_q[208:208], mem_q[209:209], mem_q[210:210], mem_q[211:211], mem_q[212:212], mem_q[213:213], mem_q[214:214], mem_q[215:215], mem_q[216:216], mem_q[217:217], mem_q[218:218], mem_q[219:219], mem_q[220:220], mem_q[221:221], mem_q[222:222], mem_q[223:223], mem_q[224:224], mem_q[225:225], mem_q[226:226], mem_q[227:227], mem_q[228:228], mem_q[229:229], mem_q[230:230], mem_q[231:231], mem_q[232:232], mem_q[233:233], mem_q[234:234], mem_q[235:235], mem_q[236:236], mem_q[237:237], mem_q[238:238], mem_q[239:239], mem_q[240:240], mem_q[241:241], mem_q[242:242], mem_q[243:243], mem_q[244:244], mem_q[245:245], mem_q[246:246], mem_q[247:247], mem_q[248:248], mem_q[249:249], mem_q[250:250], mem_q[251:251], mem_q[252:252], mem_q[253:253], mem_q[254:254], mem_q[255:255], mem_q[256:256], mem_q[257:257], mem_q[258:258], mem_q[259:259], mem_q[260:260], mem_q[261:261], mem_q[262:262], mem_q[263:263], mem_q[264:264], mem_q[265:265], mem_q[266:266], mem_q[267:267], mem_q[268:268], mem_q[269:269], mem_q[270:270], mem_q[271:271], mem_q[272:272], mem_q[273:273], mem_q[274:274], mem_q[275:275], mem_q[276:276], mem_q[277:277], mem_q[278:278], mem_q[279:279], mem_q[280:280], mem_q[281:281], mem_q[282:282], mem_q[283:283], mem_q[284:284], mem_q[285:285], mem_q[286:286], mem_q[287:287], mem_q[288:288], mem_q[289:289], mem_q[290:290], mem_q[291:291], mem_q[292:292], mem_q[293:293], mem_q[294:294], mem_q[295:295], mem_q[296:296], mem_q[297:297], mem_q[298:298], mem_q[299:299], mem_q[300:300], mem_q[301:301], mem_q[302:302], mem_q[303:303], mem_q[304:304], mem_q[305:305], mem_q[306:306], mem_q[307:307], mem_q[308:308], mem_q[309:309], mem_q[310:310], mem_q[311:311], mem_q[312:312], mem_q[313:313], mem_q[314:314], mem_q[315:315], mem_q[316:316], mem_q[317:317], mem_q[318:318], mem_q[319:319], mem_q[320:320], mem_q[321:321], mem_q[322:322], mem_q[323:323], mem_q[324:324], mem_q[325:325], mem_q[326:326], mem_q[327:327], mem_q[328:328], mem_q[329:329], mem_q[330:330], mem_q[331:331], mem_q[332:332], mem_q[333:333] } : 1'b0;
  assign N13 = N42;
  assign { N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386 } = (N14)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N385)? { mem_q[334:334], mem_q[335:335], mem_q[336:336], mem_q[337:337], mem_q[338:338], mem_q[339:339], mem_q[340:340], mem_q[341:341], mem_q[342:342], mem_q[343:343], mem_q[344:344], mem_q[345:345], mem_q[346:346], mem_q[347:347], mem_q[348:348], mem_q[349:349], mem_q[350:350], mem_q[351:351], mem_q[352:352], mem_q[353:353], mem_q[354:354], mem_q[355:355], mem_q[356:356], mem_q[357:357], mem_q[358:358], mem_q[359:359], mem_q[360:360], mem_q[361:361], mem_q[362:362], mem_q[363:363], mem_q[364:364], mem_q[365:365], mem_q[366:366], mem_q[367:367], mem_q[368:368], mem_q[369:369], mem_q[370:370], mem_q[371:371], mem_q[372:372], mem_q[373:373], mem_q[374:374], mem_q[375:375], mem_q[376:376], mem_q[377:377], mem_q[378:378], mem_q[379:379], mem_q[380:380], mem_q[381:381], mem_q[382:382], mem_q[383:383], mem_q[384:384], mem_q[385:385], mem_q[386:386], mem_q[387:387], mem_q[388:388], mem_q[389:389], mem_q[390:390], mem_q[391:391], mem_q[392:392], mem_q[393:393], mem_q[394:394], mem_q[395:395], mem_q[396:396], mem_q[397:397], mem_q[398:398], mem_q[399:399], mem_q[400:400], mem_q[401:401], mem_q[402:402], mem_q[403:403], mem_q[404:404], mem_q[405:405], mem_q[406:406], mem_q[407:407], mem_q[408:408], mem_q[409:409], mem_q[410:410], mem_q[411:411], mem_q[412:412], mem_q[413:413], mem_q[414:414], mem_q[415:415], mem_q[416:416], mem_q[417:417], mem_q[418:418], mem_q[419:419], mem_q[420:420], mem_q[421:421], mem_q[422:422], mem_q[423:423], mem_q[424:424], mem_q[425:425], mem_q[426:426], mem_q[427:427], mem_q[428:428], mem_q[429:429], mem_q[430:430], mem_q[431:431], mem_q[432:432], mem_q[433:433], mem_q[434:434], mem_q[435:435], mem_q[436:436], mem_q[437:437], mem_q[438:438], mem_q[439:439], mem_q[440:440], mem_q[441:441], mem_q[442:442], mem_q[443:443], mem_q[444:444], mem_q[445:445], mem_q[446:446], mem_q[447:447], mem_q[448:448], mem_q[449:449], mem_q[450:450], mem_q[451:451], mem_q[452:452], mem_q[453:453], mem_q[454:454], mem_q[455:455], mem_q[456:456], mem_q[457:457], mem_q[458:458], mem_q[459:459], mem_q[460:460], mem_q[461:461], mem_q[462:462], mem_q[463:463], mem_q[464:464], mem_q[465:465], mem_q[466:466], mem_q[467:467], mem_q[468:468], mem_q[469:469], mem_q[470:470], mem_q[471:471], mem_q[472:472], mem_q[473:473], mem_q[474:474], mem_q[475:475], mem_q[476:476], mem_q[477:477], mem_q[478:478], mem_q[479:479], mem_q[480:480], mem_q[481:481], mem_q[482:482], mem_q[483:483], mem_q[484:484], mem_q[485:485], mem_q[486:486], mem_q[487:487], mem_q[488:488], mem_q[489:489], mem_q[490:490], mem_q[491:491], mem_q[492:492], mem_q[493:493], mem_q[494:494], mem_q[495:495], mem_q[496:496], mem_q[497:497], mem_q[498:498], mem_q[499:499], mem_q[500:500] } : 1'b0;
  assign N14 = N43;
  assign { N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554 } = (N15)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N553)? { mem_q[501:501], mem_q[502:502], mem_q[503:503], mem_q[504:504], mem_q[505:505], mem_q[506:506], mem_q[507:507], mem_q[508:508], mem_q[509:509], mem_q[510:510], mem_q[511:511], mem_q[512:512], mem_q[513:513], mem_q[514:514], mem_q[515:515], mem_q[516:516], mem_q[517:517], mem_q[518:518], mem_q[519:519], mem_q[520:520], mem_q[521:521], mem_q[522:522], mem_q[523:523], mem_q[524:524], mem_q[525:525], mem_q[526:526], mem_q[527:527], mem_q[528:528], mem_q[529:529], mem_q[530:530], mem_q[531:531], mem_q[532:532], mem_q[533:533], mem_q[534:534], mem_q[535:535], mem_q[536:536], mem_q[537:537], mem_q[538:538], mem_q[539:539], mem_q[540:540], mem_q[541:541], mem_q[542:542], mem_q[543:543], mem_q[544:544], mem_q[545:545], mem_q[546:546], mem_q[547:547], mem_q[548:548], mem_q[549:549], mem_q[550:550], mem_q[551:551], mem_q[552:552], mem_q[553:553], mem_q[554:554], mem_q[555:555], mem_q[556:556], mem_q[557:557], mem_q[558:558], mem_q[559:559], mem_q[560:560], mem_q[561:561], mem_q[562:562], mem_q[563:563], mem_q[564:564], mem_q[565:565], mem_q[566:566], mem_q[567:567], mem_q[568:568], mem_q[569:569], mem_q[570:570], mem_q[571:571], mem_q[572:572], mem_q[573:573], mem_q[574:574], mem_q[575:575], mem_q[576:576], mem_q[577:577], mem_q[578:578], mem_q[579:579], mem_q[580:580], mem_q[581:581], mem_q[582:582], mem_q[583:583], mem_q[584:584], mem_q[585:585], mem_q[586:586], mem_q[587:587], mem_q[588:588], mem_q[589:589], mem_q[590:590], mem_q[591:591], mem_q[592:592], mem_q[593:593], mem_q[594:594], mem_q[595:595], mem_q[596:596], mem_q[597:597], mem_q[598:598], mem_q[599:599], mem_q[600:600], mem_q[601:601], mem_q[602:602], mem_q[603:603], mem_q[604:604], mem_q[605:605], mem_q[606:606], mem_q[607:607], mem_q[608:608], mem_q[609:609], mem_q[610:610], mem_q[611:611], mem_q[612:612], mem_q[613:613], mem_q[614:614], mem_q[615:615], mem_q[616:616], mem_q[617:617], mem_q[618:618], mem_q[619:619], mem_q[620:620], mem_q[621:621], mem_q[622:622], mem_q[623:623], mem_q[624:624], mem_q[625:625], mem_q[626:626], mem_q[627:627], mem_q[628:628], mem_q[629:629], mem_q[630:630], mem_q[631:631], mem_q[632:632], mem_q[633:633], mem_q[634:634], mem_q[635:635], mem_q[636:636], mem_q[637:637], mem_q[638:638], mem_q[639:639], mem_q[640:640], mem_q[641:641], mem_q[642:642], mem_q[643:643], mem_q[644:644], mem_q[645:645], mem_q[646:646], mem_q[647:647], mem_q[648:648], mem_q[649:649], mem_q[650:650], mem_q[651:651], mem_q[652:652], mem_q[653:653], mem_q[654:654], mem_q[655:655], mem_q[656:656], mem_q[657:657], mem_q[658:658], mem_q[659:659], mem_q[660:660], mem_q[661:661], mem_q[662:662], mem_q[663:663], mem_q[664:664], mem_q[665:665], mem_q[666:666], mem_q[667:667] } : 1'b0;
  assign N15 = N44;
  assign { N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722 } = (N16)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N721)? { mem_q[668:668], mem_q[669:669], mem_q[670:670], mem_q[671:671], mem_q[672:672], mem_q[673:673], mem_q[674:674], mem_q[675:675], mem_q[676:676], mem_q[677:677], mem_q[678:678], mem_q[679:679], mem_q[680:680], mem_q[681:681], mem_q[682:682], mem_q[683:683], mem_q[684:684], mem_q[685:685], mem_q[686:686], mem_q[687:687], mem_q[688:688], mem_q[689:689], mem_q[690:690], mem_q[691:691], mem_q[692:692], mem_q[693:693], mem_q[694:694], mem_q[695:695], mem_q[696:696], mem_q[697:697], mem_q[698:698], mem_q[699:699], mem_q[700:700], mem_q[701:701], mem_q[702:702], mem_q[703:703], mem_q[704:704], mem_q[705:705], mem_q[706:706], mem_q[707:707], mem_q[708:708], mem_q[709:709], mem_q[710:710], mem_q[711:711], mem_q[712:712], mem_q[713:713], mem_q[714:714], mem_q[715:715], mem_q[716:716], mem_q[717:717], mem_q[718:718], mem_q[719:719], mem_q[720:720], mem_q[721:721], mem_q[722:722], mem_q[723:723], mem_q[724:724], mem_q[725:725], mem_q[726:726], mem_q[727:727], mem_q[728:728], mem_q[729:729], mem_q[730:730], mem_q[731:731], mem_q[732:732], mem_q[733:733], mem_q[734:734], mem_q[735:735], mem_q[736:736], mem_q[737:737], mem_q[738:738], mem_q[739:739], mem_q[740:740], mem_q[741:741], mem_q[742:742], mem_q[743:743], mem_q[744:744], mem_q[745:745], mem_q[746:746], mem_q[747:747], mem_q[748:748], mem_q[749:749], mem_q[750:750], mem_q[751:751], mem_q[752:752], mem_q[753:753], mem_q[754:754], mem_q[755:755], mem_q[756:756], mem_q[757:757], mem_q[758:758], mem_q[759:759], mem_q[760:760], mem_q[761:761], mem_q[762:762], mem_q[763:763], mem_q[764:764], mem_q[765:765], mem_q[766:766], mem_q[767:767], mem_q[768:768], mem_q[769:769], mem_q[770:770], mem_q[771:771], mem_q[772:772], mem_q[773:773], mem_q[774:774], mem_q[775:775], mem_q[776:776], mem_q[777:777], mem_q[778:778], mem_q[779:779], mem_q[780:780], mem_q[781:781], mem_q[782:782], mem_q[783:783], mem_q[784:784], mem_q[785:785], mem_q[786:786], mem_q[787:787], mem_q[788:788], mem_q[789:789], mem_q[790:790], mem_q[791:791], mem_q[792:792], mem_q[793:793], mem_q[794:794], mem_q[795:795], mem_q[796:796], mem_q[797:797], mem_q[798:798], mem_q[799:799], mem_q[800:800], mem_q[801:801], mem_q[802:802], mem_q[803:803], mem_q[804:804], mem_q[805:805], mem_q[806:806], mem_q[807:807], mem_q[808:808], mem_q[809:809], mem_q[810:810], mem_q[811:811], mem_q[812:812], mem_q[813:813], mem_q[814:814], mem_q[815:815], mem_q[816:816], mem_q[817:817], mem_q[818:818], mem_q[819:819], mem_q[820:820], mem_q[821:821], mem_q[822:822], mem_q[823:823], mem_q[824:824], mem_q[825:825], mem_q[826:826], mem_q[827:827], mem_q[828:828], mem_q[829:829], mem_q[830:830], mem_q[831:831], mem_q[832:832], mem_q[833:833], mem_q[834:834] } : 1'b0;
  assign N16 = N45;
  assign { N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890 } = (N17)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (N889)? { mem_q[835:835], mem_q[836:836], mem_q[837:837], mem_q[838:838], mem_q[839:839], mem_q[840:840], mem_q[841:841], mem_q[842:842], mem_q[843:843], mem_q[844:844], mem_q[845:845], mem_q[846:846], mem_q[847:847], mem_q[848:848], mem_q[849:849], mem_q[850:850], mem_q[851:851], mem_q[852:852], mem_q[853:853], mem_q[854:854], mem_q[855:855], mem_q[856:856], mem_q[857:857], mem_q[858:858], mem_q[859:859], mem_q[860:860], mem_q[861:861], mem_q[862:862], mem_q[863:863], mem_q[864:864], mem_q[865:865], mem_q[866:866], mem_q[867:867], mem_q[868:868], mem_q[869:869], mem_q[870:870], mem_q[871:871], mem_q[872:872], mem_q[873:873], mem_q[874:874], mem_q[875:875], mem_q[876:876], mem_q[877:877], mem_q[878:878], mem_q[879:879], mem_q[880:880], mem_q[881:881], mem_q[882:882], mem_q[883:883], mem_q[884:884], mem_q[885:885], mem_q[886:886], mem_q[887:887], mem_q[888:888], mem_q[889:889], mem_q[890:890], mem_q[891:891], mem_q[892:892], mem_q[893:893], mem_q[894:894], mem_q[895:895], mem_q[896:896], mem_q[897:897], mem_q[898:898], mem_q[899:899], mem_q[900:900], mem_q[901:901], mem_q[902:902], mem_q[903:903], mem_q[904:904], mem_q[905:905], mem_q[906:906], mem_q[907:907], mem_q[908:908], mem_q[909:909], mem_q[910:910], mem_q[911:911], mem_q[912:912], mem_q[913:913], mem_q[914:914], mem_q[915:915], mem_q[916:916], mem_q[917:917], mem_q[918:918], mem_q[919:919], mem_q[920:920], mem_q[921:921], mem_q[922:922], mem_q[923:923], mem_q[924:924], mem_q[925:925], mem_q[926:926], mem_q[927:927], mem_q[928:928], mem_q[929:929], mem_q[930:930], mem_q[931:931], mem_q[932:932], mem_q[933:933], mem_q[934:934], mem_q[935:935], mem_q[936:936], mem_q[937:937], mem_q[938:938], mem_q[939:939], mem_q[940:940], mem_q[941:941], mem_q[942:942], mem_q[943:943], mem_q[944:944], mem_q[945:945], mem_q[946:946], mem_q[947:947], mem_q[948:948], mem_q[949:949], mem_q[950:950], mem_q[951:951], mem_q[952:952], mem_q[953:953], mem_q[954:954], mem_q[955:955], mem_q[956:956], mem_q[957:957], mem_q[958:958], mem_q[959:959], mem_q[960:960], mem_q[961:961], mem_q[962:962], mem_q[963:963], mem_q[964:964], mem_q[965:965], mem_q[966:966], mem_q[967:967], mem_q[968:968], mem_q[969:969], mem_q[970:970], mem_q[971:971], mem_q[972:972], mem_q[973:973], mem_q[974:974], mem_q[975:975], mem_q[976:976], mem_q[977:977], mem_q[978:978], mem_q[979:979], mem_q[980:980], mem_q[981:981], mem_q[982:982], mem_q[983:983], mem_q[984:984], mem_q[985:985], mem_q[986:986], mem_q[987:987], mem_q[988:988], mem_q[989:989], mem_q[990:990], mem_q[991:991], mem_q[992:992], mem_q[993:993], mem_q[994:994], mem_q[995:995], mem_q[996:996], mem_q[997:997], mem_q[998:998], mem_q[999:999], mem_q[1000:1000], mem_q[1001:1001] } : 1'b0;
  assign N17 = N46;
  assign { N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058 } = (N18)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (N1057)? { mem_q[1002:1002], mem_q[1003:1003], mem_q[1004:1004], mem_q[1005:1005], mem_q[1006:1006], mem_q[1007:1007], mem_q[1008:1008], mem_q[1009:1009], mem_q[1010:1010], mem_q[1011:1011], mem_q[1012:1012], mem_q[1013:1013], mem_q[1014:1014], mem_q[1015:1015], mem_q[1016:1016], mem_q[1017:1017], mem_q[1018:1018], mem_q[1019:1019], mem_q[1020:1020], mem_q[1021:1021], mem_q[1022:1022], mem_q[1023:1023], mem_q[1024:1024], mem_q[1025:1025], mem_q[1026:1026], mem_q[1027:1027], mem_q[1028:1028], mem_q[1029:1029], mem_q[1030:1030], mem_q[1031:1031], mem_q[1032:1032], mem_q[1033:1033], mem_q[1034:1034], mem_q[1035:1035], mem_q[1036:1036], mem_q[1037:1037], mem_q[1038:1038], mem_q[1039:1039], mem_q[1040:1040], mem_q[1041:1041], mem_q[1042:1042], mem_q[1043:1043], mem_q[1044:1044], mem_q[1045:1045], mem_q[1046:1046], mem_q[1047:1047], mem_q[1048:1048], mem_q[1049:1049], mem_q[1050:1050], mem_q[1051:1051], mem_q[1052:1052], mem_q[1053:1053], mem_q[1054:1054], mem_q[1055:1055], mem_q[1056:1056], mem_q[1057:1057], mem_q[1058:1058], mem_q[1059:1059], mem_q[1060:1060], mem_q[1061:1061], mem_q[1062:1062], mem_q[1063:1063], mem_q[1064:1064], mem_q[1065:1065], mem_q[1066:1066], mem_q[1067:1067], mem_q[1068:1068], mem_q[1069:1069], mem_q[1070:1070], mem_q[1071:1071], mem_q[1072:1072], mem_q[1073:1073], mem_q[1074:1074], mem_q[1075:1075], mem_q[1076:1076], mem_q[1077:1077], mem_q[1078:1078], mem_q[1079:1079], mem_q[1080:1080], mem_q[1081:1081], mem_q[1082:1082], mem_q[1083:1083], mem_q[1084:1084], mem_q[1085:1085], mem_q[1086:1086], mem_q[1087:1087], mem_q[1088:1088], mem_q[1089:1089], mem_q[1090:1090], mem_q[1091:1091], mem_q[1092:1092], mem_q[1093:1093], mem_q[1094:1094], mem_q[1095:1095], mem_q[1096:1096], mem_q[1097:1097], mem_q[1098:1098], mem_q[1099:1099], mem_q[1100:1100], mem_q[1101:1101], mem_q[1102:1102], mem_q[1103:1103], mem_q[1104:1104], mem_q[1105:1105], mem_q[1106:1106], mem_q[1107:1107], mem_q[1108:1108], mem_q[1109:1109], mem_q[1110:1110], mem_q[1111:1111], mem_q[1112:1112], mem_q[1113:1113], mem_q[1114:1114], mem_q[1115:1115], mem_q[1116:1116], mem_q[1117:1117], mem_q[1118:1118], mem_q[1119:1119], mem_q[1120:1120], mem_q[1121:1121], mem_q[1122:1122], mem_q[1123:1123], mem_q[1124:1124], mem_q[1125:1125], mem_q[1126:1126], mem_q[1127:1127], mem_q[1128:1128], mem_q[1129:1129], mem_q[1130:1130], mem_q[1131:1131], mem_q[1132:1132], mem_q[1133:1133], mem_q[1134:1134], mem_q[1135:1135], mem_q[1136:1136], mem_q[1137:1137], mem_q[1138:1138], mem_q[1139:1139], mem_q[1140:1140], mem_q[1141:1141], mem_q[1142:1142], mem_q[1143:1143], mem_q[1144:1144], mem_q[1145:1145], mem_q[1146:1146], mem_q[1147:1147], mem_q[1148:1148], mem_q[1149:1149], mem_q[1150:1150], mem_q[1151:1151], mem_q[1152:1152], mem_q[1153:1153], mem_q[1154:1154], mem_q[1155:1155], mem_q[1156:1156], mem_q[1157:1157], mem_q[1158:1158], mem_q[1159:1159], mem_q[1160:1160], mem_q[1161:1161], mem_q[1162:1162], mem_q[1163:1163], mem_q[1164:1164], mem_q[1165:1165], mem_q[1166:1166], mem_q[1167:1167], mem_q[1168:1168] } : 1'b0;
  assign N18 = N47;
  assign { N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226 } = (N19)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63], data_i[64:64], data_i[65:65], data_i[66:66], data_i[67:67], data_i[68:68], data_i[69:69], data_i[70:70], data_i[71:71], data_i[72:72], data_i[73:73], data_i[74:74], data_i[75:75], data_i[76:76], data_i[77:77], data_i[78:78], data_i[79:79], data_i[80:80], data_i[81:81], data_i[82:82], data_i[83:83], data_i[84:84], data_i[85:85], data_i[86:86], data_i[87:87], data_i[88:88], data_i[89:89], data_i[90:90], data_i[91:91], data_i[92:92], data_i[93:93], data_i[94:94], data_i[95:95], data_i[96:96], data_i[97:97], data_i[98:98], data_i[99:99], data_i[100:100], data_i[101:101], data_i[102:102], data_i[103:103], data_i[104:104], data_i[105:105], data_i[106:106], data_i[107:107], data_i[108:108], data_i[109:109], data_i[110:110], data_i[111:111], data_i[112:112], data_i[113:113], data_i[114:114], data_i[115:115], data_i[116:116], data_i[117:117], data_i[118:118], data_i[119:119], data_i[120:120], data_i[121:121], data_i[122:122], data_i[123:123], data_i[124:124], data_i[125:125], data_i[126:126], data_i[127:127], data_i[128:128], data_i[129:129], data_i[130:130], data_i[131:131], data_i[132:132], data_i[133:133], data_i[134:134], data_i[135:135], data_i[136:136], data_i[137:137], data_i[138:138], data_i[139:139], data_i[140:140], data_i[141:141], data_i[142:142], data_i[143:143], data_i[144:144], data_i[145:145], data_i[146:146], data_i[147:147], data_i[148:148], data_i[149:149], data_i[150:150], data_i[151:151], data_i[152:152], data_i[153:153], data_i[154:154], data_i[155:155], data_i[156:156], data_i[157:157], data_i[158:158], data_i[159:159], data_i[160:160], data_i[161:161], data_i[162:162], data_i[163:163], data_i[164:164], data_i[165:165], data_i[166:166] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               (N1225)? { mem_q[1169:1169], mem_q[1170:1170], mem_q[1171:1171], mem_q[1172:1172], mem_q[1173:1173], mem_q[1174:1174], mem_q[1175:1175], mem_q[1176:1176], mem_q[1177:1177], mem_q[1178:1178], mem_q[1179:1179], mem_q[1180:1180], mem_q[1181:1181], mem_q[1182:1182], mem_q[1183:1183], mem_q[1184:1184], mem_q[1185:1185], mem_q[1186:1186], mem_q[1187:1187], mem_q[1188:1188], mem_q[1189:1189], mem_q[1190:1190], mem_q[1191:1191], mem_q[1192:1192], mem_q[1193:1193], mem_q[1194:1194], mem_q[1195:1195], mem_q[1196:1196], mem_q[1197:1197], mem_q[1198:1198], mem_q[1199:1199], mem_q[1200:1200], mem_q[1201:1201], mem_q[1202:1202], mem_q[1203:1203], mem_q[1204:1204], mem_q[1205:1205], mem_q[1206:1206], mem_q[1207:1207], mem_q[1208:1208], mem_q[1209:1209], mem_q[1210:1210], mem_q[1211:1211], mem_q[1212:1212], mem_q[1213:1213], mem_q[1214:1214], mem_q[1215:1215], mem_q[1216:1216], mem_q[1217:1217], mem_q[1218:1218], mem_q[1219:1219], mem_q[1220:1220], mem_q[1221:1221], mem_q[1222:1222], mem_q[1223:1223], mem_q[1224:1224], mem_q[1225:1225], mem_q[1226:1226], mem_q[1227:1227], mem_q[1228:1228], mem_q[1229:1229], mem_q[1230:1230], mem_q[1231:1231], mem_q[1232:1232], mem_q[1233:1233], mem_q[1234:1234], mem_q[1235:1235], mem_q[1236:1236], mem_q[1237:1237], mem_q[1238:1238], mem_q[1239:1239], mem_q[1240:1240], mem_q[1241:1241], mem_q[1242:1242], mem_q[1243:1243], mem_q[1244:1244], mem_q[1245:1245], mem_q[1246:1246], mem_q[1247:1247], mem_q[1248:1248], mem_q[1249:1249], mem_q[1250:1250], mem_q[1251:1251], mem_q[1252:1252], mem_q[1253:1253], mem_q[1254:1254], mem_q[1255:1255], mem_q[1256:1256], mem_q[1257:1257], mem_q[1258:1258], mem_q[1259:1259], mem_q[1260:1260], mem_q[1261:1261], mem_q[1262:1262], mem_q[1263:1263], mem_q[1264:1264], mem_q[1265:1265], mem_q[1266:1266], mem_q[1267:1267], mem_q[1268:1268], mem_q[1269:1269], mem_q[1270:1270], mem_q[1271:1271], mem_q[1272:1272], mem_q[1273:1273], mem_q[1274:1274], mem_q[1275:1275], mem_q[1276:1276], mem_q[1277:1277], mem_q[1278:1278], mem_q[1279:1279], mem_q[1280:1280], mem_q[1281:1281], mem_q[1282:1282], mem_q[1283:1283], mem_q[1284:1284], mem_q[1285:1285], mem_q[1286:1286], mem_q[1287:1287], mem_q[1288:1288], mem_q[1289:1289], mem_q[1290:1290], mem_q[1291:1291], mem_q[1292:1292], mem_q[1293:1293], mem_q[1294:1294], mem_q[1295:1295], mem_q[1296:1296], mem_q[1297:1297], mem_q[1298:1298], mem_q[1299:1299], mem_q[1300:1300], mem_q[1301:1301], mem_q[1302:1302], mem_q[1303:1303], mem_q[1304:1304], mem_q[1305:1305], mem_q[1306:1306], mem_q[1307:1307], mem_q[1308:1308], mem_q[1309:1309], mem_q[1310:1310], mem_q[1311:1311], mem_q[1312:1312], mem_q[1313:1313], mem_q[1314:1314], mem_q[1315:1315], mem_q[1316:1316], mem_q[1317:1317], mem_q[1318:1318], mem_q[1319:1319], mem_q[1320:1320], mem_q[1321:1321], mem_q[1322:1322], mem_q[1323:1323], mem_q[1324:1324], mem_q[1325:1325], mem_q[1326:1326], mem_q[1327:1327], mem_q[1328:1328], mem_q[1329:1329], mem_q[1330:1330], mem_q[1331:1331], mem_q[1332:1332], mem_q[1333:1333], mem_q[1334:1334], mem_q[1335:1335] } : 1'b0;
  assign N19 = N48;
  assign mem_n = (N20)? { N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216 } : 
                 (N40)? mem_q : 1'b0;
  assign N20 = N39;
  assign gate_clock = ~N39;
  assign { N1412, N1411, N1410, N1409 } = (N21)? { N1408, N1407, N1406, N1405 } : 
                                          (N1401)? { N1399, N1398, N1397, N1396 } : 1'b0;
  assign N21 = N1400;
  assign { N1419, N1418, N1417 } = (N22)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N23)? { N1404, N1403, N1402 } : 1'b0;
  assign N22 = flush_i;
  assign N23 = N1416;
  assign { N1422, N1421, N1420 } = (N22)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N23)? { N1395, N1394, N1393 } : 1'b0;
  assign { N1426, N1425, N1424, N1423 } = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                          (N23)? { N1412, N1411, N1410, N1409 } : 1'b0;
  assign N24 = ~read_pointer_q[0];
  assign N25 = ~read_pointer_q[1];
  assign N26 = N24 & N25;
  assign N27 = N24 & read_pointer_q[1];
  assign N28 = read_pointer_q[0] & N25;
  assign N29 = read_pointer_q[0] & read_pointer_q[1];
  assign N30 = ~read_pointer_q[2];
  assign N31 = N26 & N30;
  assign N32 = N26 & read_pointer_q[2];
  assign N33 = N28 & N30;
  assign N34 = N28 & read_pointer_q[2];
  assign N35 = N27 & N30;
  assign N36 = N27 & read_pointer_q[2];
  assign N37 = N29 & N30;
  assign N38 = N29 & read_pointer_q[2];
  assign N39 = push_i & N1445;
  assign N40 = ~N39;
  assign N49 = ~N41;
  assign N217 = ~N42;
  assign N385 = ~N43;
  assign N553 = ~N44;
  assign N721 = ~N45;
  assign N889 = ~N46;
  assign N1057 = ~N47;
  assign N1225 = ~N48;
  assign N1400 = pop_i & N1440;
  assign N1401 = ~N1400;
  assign N1413 = N1456 & N1440;
  assign N1456 = N1455 & N1445;
  assign N1455 = push_i & pop_i;
  assign N1414 = ~N1413;
  assign N1415 = ~rst_ni;
  assign N1416 = ~flush_i;
  assign N1427 = ~gate_clock;
  assign N1428 = N1413 & N1416;
  assign N1429 = N1414 & N1416;
  assign N1430 = N1401 & N1429;
  assign N1431 = N40 & N1430;
  assign N1432 = N1428 | N1431;
  assign N1433 = ~N1432;
  assign N1434 = N1401 & N1416;
  assign N1435 = ~N1434;
  assign N1436 = N40 & N1416;
  assign N1437 = ~N1436;

endmodule