module load_unit
(
  clk_i,
  rst_ni,
  flush_i,
  valid_i,
  lsu_ctrl_i,
  pop_ld_o,
  valid_o,
  trans_id_o,
  result_o,
  ex_o,
  translation_req_o,
  vaddr_o,
  paddr_i,
  ex_i,
  dtlb_hit_i,
  page_offset_o,
  page_offset_matches_i,
  req_port_i,
  req_port_o
);

  input [150:0] lsu_ctrl_i;
  output [2:0] trans_id_o;
  output [63:0] result_o;
  output [128:0] ex_o;
  output [63:0] vaddr_o;
  input [63:0] paddr_i;
  input [128:0] ex_i;
  output [11:0] page_offset_o;
  input [65:0] req_port_i;
  output [133:0] req_port_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input valid_i;
  input dtlb_hit_i;
  input page_offset_matches_i;
  output pop_ld_o;
  output valid_o;
  output translation_req_o;
  wire [2:0] trans_id_o,state_d,idx_d;
  wire [63:0] result_o,vaddr_o;
  wire [128:0] ex_o;
  wire [11:0] page_offset_o;
  wire [133:0] req_port_o;
  wire pop_ld_o,valid_o,translation_req_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,
  N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,
  N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,
  N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,
  N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,
  N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,
  N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,
  N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,
  N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,
  N223,N224,N225,N226,N227,N228,signed_d,N229,N230,N231,N232,N233,N234,N235,N236,
  N237,N238,N239,fp_sign_d,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,sign_bit,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487;
  wire [12:0] load_data_d;
  wire [63:8] shifted_data;
  reg [12:0] load_data_q;
  reg [2:0] state_q,idx_q;
  reg n__tmp493,signed_q,fp_sign_q;
  assign req_port_o[14] = 1'b0;
  assign req_port_o[15] = 1'b0;
  assign req_port_o[16] = 1'b0;
  assign req_port_o[17] = 1'b0;
  assign req_port_o[18] = 1'b0;
  assign req_port_o[19] = 1'b0;
  assign req_port_o[20] = 1'b0;
  assign req_port_o[21] = 1'b0;
  assign req_port_o[22] = 1'b0;
  assign req_port_o[23] = 1'b0;
  assign req_port_o[24] = 1'b0;
  assign req_port_o[25] = 1'b0;
  assign req_port_o[26] = 1'b0;
  assign req_port_o[27] = 1'b0;
  assign req_port_o[28] = 1'b0;
  assign req_port_o[29] = 1'b0;
  assign req_port_o[30] = 1'b0;
  assign req_port_o[31] = 1'b0;
  assign req_port_o[32] = 1'b0;
  assign req_port_o[33] = 1'b0;
  assign req_port_o[34] = 1'b0;
  assign req_port_o[35] = 1'b0;
  assign req_port_o[36] = 1'b0;
  assign req_port_o[37] = 1'b0;
  assign req_port_o[38] = 1'b0;
  assign req_port_o[39] = 1'b0;
  assign req_port_o[40] = 1'b0;
  assign req_port_o[41] = 1'b0;
  assign req_port_o[42] = 1'b0;
  assign req_port_o[43] = 1'b0;
  assign req_port_o[44] = 1'b0;
  assign req_port_o[45] = 1'b0;
  assign req_port_o[46] = 1'b0;
  assign req_port_o[47] = 1'b0;
  assign req_port_o[48] = 1'b0;
  assign req_port_o[49] = 1'b0;
  assign req_port_o[50] = 1'b0;
  assign req_port_o[51] = 1'b0;
  assign req_port_o[52] = 1'b0;
  assign req_port_o[53] = 1'b0;
  assign req_port_o[54] = 1'b0;
  assign req_port_o[55] = 1'b0;
  assign req_port_o[56] = 1'b0;
  assign req_port_o[57] = 1'b0;
  assign req_port_o[58] = 1'b0;
  assign req_port_o[59] = 1'b0;
  assign req_port_o[60] = 1'b0;
  assign req_port_o[61] = 1'b0;
  assign req_port_o[62] = 1'b0;
  assign req_port_o[63] = 1'b0;
  assign req_port_o[64] = 1'b0;
  assign req_port_o[65] = 1'b0;
  assign req_port_o[66] = 1'b0;
  assign req_port_o[67] = 1'b0;
  assign req_port_o[68] = 1'b0;
  assign req_port_o[69] = 1'b0;
  assign req_port_o[70] = 1'b0;
  assign req_port_o[71] = 1'b0;
  assign req_port_o[72] = 1'b0;
  assign req_port_o[73] = 1'b0;
  assign req_port_o[74] = 1'b0;
  assign req_port_o[75] = 1'b0;
  assign req_port_o[76] = 1'b0;
  assign req_port_o[77] = 1'b0;
  assign req_port_o[12] = 1'b0;
  assign req_port_o[133] = lsu_ctrl_i[97];
  assign vaddr_o[11] = lsu_ctrl_i[97];
  assign page_offset_o[11] = lsu_ctrl_i[97];
  assign req_port_o[132] = lsu_ctrl_i[96];
  assign vaddr_o[10] = lsu_ctrl_i[96];
  assign page_offset_o[10] = lsu_ctrl_i[96];
  assign req_port_o[131] = lsu_ctrl_i[95];
  assign vaddr_o[9] = lsu_ctrl_i[95];
  assign page_offset_o[9] = lsu_ctrl_i[95];
  assign req_port_o[130] = lsu_ctrl_i[94];
  assign vaddr_o[8] = lsu_ctrl_i[94];
  assign page_offset_o[8] = lsu_ctrl_i[94];
  assign req_port_o[129] = lsu_ctrl_i[93];
  assign vaddr_o[7] = lsu_ctrl_i[93];
  assign page_offset_o[7] = lsu_ctrl_i[93];
  assign req_port_o[128] = lsu_ctrl_i[92];
  assign vaddr_o[6] = lsu_ctrl_i[92];
  assign page_offset_o[6] = lsu_ctrl_i[92];
  assign req_port_o[127] = lsu_ctrl_i[91];
  assign vaddr_o[5] = lsu_ctrl_i[91];
  assign page_offset_o[5] = lsu_ctrl_i[91];
  assign req_port_o[126] = lsu_ctrl_i[90];
  assign vaddr_o[4] = lsu_ctrl_i[90];
  assign page_offset_o[4] = lsu_ctrl_i[90];
  assign req_port_o[125] = lsu_ctrl_i[89];
  assign vaddr_o[3] = lsu_ctrl_i[89];
  assign page_offset_o[3] = lsu_ctrl_i[89];
  assign req_port_o[124] = lsu_ctrl_i[88];
  assign vaddr_o[2] = lsu_ctrl_i[88];
  assign page_offset_o[2] = lsu_ctrl_i[88];
  assign req_port_o[123] = lsu_ctrl_i[87];
  assign vaddr_o[1] = lsu_ctrl_i[87];
  assign page_offset_o[1] = lsu_ctrl_i[87];
  assign req_port_o[122] = lsu_ctrl_i[86];
  assign vaddr_o[0] = lsu_ctrl_i[86];
  assign page_offset_o[0] = lsu_ctrl_i[86];
  assign vaddr_o[63] = lsu_ctrl_i[149];
  assign vaddr_o[62] = lsu_ctrl_i[148];
  assign vaddr_o[61] = lsu_ctrl_i[147];
  assign vaddr_o[60] = lsu_ctrl_i[146];
  assign vaddr_o[59] = lsu_ctrl_i[145];
  assign vaddr_o[58] = lsu_ctrl_i[144];
  assign vaddr_o[57] = lsu_ctrl_i[143];
  assign vaddr_o[56] = lsu_ctrl_i[142];
  assign vaddr_o[55] = lsu_ctrl_i[141];
  assign vaddr_o[54] = lsu_ctrl_i[140];
  assign vaddr_o[53] = lsu_ctrl_i[139];
  assign vaddr_o[52] = lsu_ctrl_i[138];
  assign vaddr_o[51] = lsu_ctrl_i[137];
  assign vaddr_o[50] = lsu_ctrl_i[136];
  assign vaddr_o[49] = lsu_ctrl_i[135];
  assign vaddr_o[48] = lsu_ctrl_i[134];
  assign vaddr_o[47] = lsu_ctrl_i[133];
  assign vaddr_o[46] = lsu_ctrl_i[132];
  assign vaddr_o[45] = lsu_ctrl_i[131];
  assign vaddr_o[44] = lsu_ctrl_i[130];
  assign vaddr_o[43] = lsu_ctrl_i[129];
  assign vaddr_o[42] = lsu_ctrl_i[128];
  assign vaddr_o[41] = lsu_ctrl_i[127];
  assign vaddr_o[40] = lsu_ctrl_i[126];
  assign vaddr_o[39] = lsu_ctrl_i[125];
  assign vaddr_o[38] = lsu_ctrl_i[124];
  assign vaddr_o[37] = lsu_ctrl_i[123];
  assign vaddr_o[36] = lsu_ctrl_i[122];
  assign vaddr_o[35] = lsu_ctrl_i[121];
  assign vaddr_o[34] = lsu_ctrl_i[120];
  assign vaddr_o[33] = lsu_ctrl_i[119];
  assign vaddr_o[32] = lsu_ctrl_i[118];
  assign vaddr_o[31] = lsu_ctrl_i[117];
  assign vaddr_o[30] = lsu_ctrl_i[116];
  assign vaddr_o[29] = lsu_ctrl_i[115];
  assign vaddr_o[28] = lsu_ctrl_i[114];
  assign vaddr_o[27] = lsu_ctrl_i[113];
  assign vaddr_o[26] = lsu_ctrl_i[112];
  assign vaddr_o[25] = lsu_ctrl_i[111];
  assign vaddr_o[24] = lsu_ctrl_i[110];
  assign vaddr_o[23] = lsu_ctrl_i[109];
  assign vaddr_o[22] = lsu_ctrl_i[108];
  assign vaddr_o[21] = lsu_ctrl_i[107];
  assign vaddr_o[20] = lsu_ctrl_i[106];
  assign vaddr_o[19] = lsu_ctrl_i[105];
  assign vaddr_o[18] = lsu_ctrl_i[104];
  assign vaddr_o[17] = lsu_ctrl_i[103];
  assign vaddr_o[16] = lsu_ctrl_i[102];
  assign vaddr_o[15] = lsu_ctrl_i[101];
  assign vaddr_o[14] = lsu_ctrl_i[100];
  assign vaddr_o[13] = lsu_ctrl_i[99];
  assign vaddr_o[12] = lsu_ctrl_i[98];
  assign req_port_o[11] = lsu_ctrl_i[21];
  assign req_port_o[10] = lsu_ctrl_i[20];
  assign req_port_o[9] = lsu_ctrl_i[19];
  assign req_port_o[8] = lsu_ctrl_i[18];
  assign req_port_o[7] = lsu_ctrl_i[17];
  assign req_port_o[6] = lsu_ctrl_i[16];
  assign req_port_o[5] = lsu_ctrl_i[15];
  assign req_port_o[4] = lsu_ctrl_i[14];
  assign ex_o[128] = ex_i[128];
  assign ex_o[127] = ex_i[127];
  assign ex_o[126] = ex_i[126];
  assign ex_o[125] = ex_i[125];
  assign ex_o[124] = ex_i[124];
  assign ex_o[123] = ex_i[123];
  assign ex_o[122] = ex_i[122];
  assign ex_o[121] = ex_i[121];
  assign ex_o[120] = ex_i[120];
  assign ex_o[119] = ex_i[119];
  assign ex_o[118] = ex_i[118];
  assign ex_o[117] = ex_i[117];
  assign ex_o[116] = ex_i[116];
  assign ex_o[115] = ex_i[115];
  assign ex_o[114] = ex_i[114];
  assign ex_o[113] = ex_i[113];
  assign ex_o[112] = ex_i[112];
  assign ex_o[111] = ex_i[111];
  assign ex_o[110] = ex_i[110];
  assign ex_o[109] = ex_i[109];
  assign ex_o[108] = ex_i[108];
  assign ex_o[107] = ex_i[107];
  assign ex_o[106] = ex_i[106];
  assign ex_o[105] = ex_i[105];
  assign ex_o[104] = ex_i[104];
  assign ex_o[103] = ex_i[103];
  assign ex_o[102] = ex_i[102];
  assign ex_o[101] = ex_i[101];
  assign ex_o[100] = ex_i[100];
  assign ex_o[99] = ex_i[99];
  assign ex_o[98] = ex_i[98];
  assign ex_o[97] = ex_i[97];
  assign ex_o[96] = ex_i[96];
  assign ex_o[95] = ex_i[95];
  assign ex_o[94] = ex_i[94];
  assign ex_o[93] = ex_i[93];
  assign ex_o[92] = ex_i[92];
  assign ex_o[91] = ex_i[91];
  assign ex_o[90] = ex_i[90];
  assign ex_o[89] = ex_i[89];
  assign ex_o[88] = ex_i[88];
  assign ex_o[87] = ex_i[87];
  assign ex_o[86] = ex_i[86];
  assign ex_o[85] = ex_i[85];
  assign ex_o[84] = ex_i[84];
  assign ex_o[83] = ex_i[83];
  assign ex_o[82] = ex_i[82];
  assign ex_o[81] = ex_i[81];
  assign ex_o[80] = ex_i[80];
  assign ex_o[79] = ex_i[79];
  assign ex_o[78] = ex_i[78];
  assign ex_o[77] = ex_i[77];
  assign ex_o[76] = ex_i[76];
  assign ex_o[75] = ex_i[75];
  assign ex_o[74] = ex_i[74];
  assign ex_o[73] = ex_i[73];
  assign ex_o[72] = ex_i[72];
  assign ex_o[71] = ex_i[71];
  assign ex_o[70] = ex_i[70];
  assign ex_o[69] = ex_i[69];
  assign ex_o[68] = ex_i[68];
  assign ex_o[67] = ex_i[67];
  assign ex_o[66] = ex_i[66];
  assign ex_o[65] = ex_i[65];
  assign ex_o[64] = ex_i[64];
  assign ex_o[63] = ex_i[63];
  assign ex_o[62] = ex_i[62];
  assign ex_o[61] = ex_i[61];
  assign ex_o[60] = ex_i[60];
  assign ex_o[59] = ex_i[59];
  assign ex_o[58] = ex_i[58];
  assign ex_o[57] = ex_i[57];
  assign ex_o[56] = ex_i[56];
  assign ex_o[55] = ex_i[55];
  assign ex_o[54] = ex_i[54];
  assign ex_o[53] = ex_i[53];
  assign ex_o[52] = ex_i[52];
  assign ex_o[51] = ex_i[51];
  assign ex_o[50] = ex_i[50];
  assign ex_o[49] = ex_i[49];
  assign ex_o[48] = ex_i[48];
  assign ex_o[47] = ex_i[47];
  assign ex_o[46] = ex_i[46];
  assign ex_o[45] = ex_i[45];
  assign ex_o[44] = ex_i[44];
  assign ex_o[43] = ex_i[43];
  assign ex_o[42] = ex_i[42];
  assign ex_o[41] = ex_i[41];
  assign ex_o[40] = ex_i[40];
  assign ex_o[39] = ex_i[39];
  assign ex_o[38] = ex_i[38];
  assign ex_o[37] = ex_i[37];
  assign ex_o[36] = ex_i[36];
  assign ex_o[35] = ex_i[35];
  assign ex_o[34] = ex_i[34];
  assign ex_o[33] = ex_i[33];
  assign ex_o[32] = ex_i[32];
  assign ex_o[31] = ex_i[31];
  assign ex_o[30] = ex_i[30];
  assign ex_o[29] = ex_i[29];
  assign ex_o[28] = ex_i[28];
  assign ex_o[27] = ex_i[27];
  assign ex_o[26] = ex_i[26];
  assign ex_o[25] = ex_i[25];
  assign ex_o[24] = ex_i[24];
  assign ex_o[23] = ex_i[23];
  assign ex_o[22] = ex_i[22];
  assign ex_o[21] = ex_i[21];
  assign ex_o[20] = ex_i[20];
  assign ex_o[19] = ex_i[19];
  assign ex_o[18] = ex_i[18];
  assign ex_o[17] = ex_i[17];
  assign ex_o[16] = ex_i[16];
  assign ex_o[15] = ex_i[15];
  assign ex_o[14] = ex_i[14];
  assign ex_o[13] = ex_i[13];
  assign ex_o[12] = ex_i[12];
  assign ex_o[11] = ex_i[11];
  assign ex_o[10] = ex_i[10];
  assign ex_o[9] = ex_i[9];
  assign ex_o[8] = ex_i[8];
  assign ex_o[7] = ex_i[7];
  assign ex_o[6] = ex_i[6];
  assign ex_o[5] = ex_i[5];
  assign ex_o[4] = ex_i[4];
  assign ex_o[3] = ex_i[3];
  assign ex_o[2] = ex_i[2];
  assign ex_o[1] = ex_i[1];
  assign ex_o[0] = ex_i[0];
  assign req_port_o[121] = paddr_i[55];
  assign req_port_o[120] = paddr_i[54];
  assign req_port_o[119] = paddr_i[53];
  assign req_port_o[118] = paddr_i[52];
  assign req_port_o[117] = paddr_i[51];
  assign req_port_o[116] = paddr_i[50];
  assign req_port_o[115] = paddr_i[49];
  assign req_port_o[114] = paddr_i[48];
  assign req_port_o[113] = paddr_i[47];
  assign req_port_o[112] = paddr_i[46];
  assign req_port_o[111] = paddr_i[45];
  assign req_port_o[110] = paddr_i[44];
  assign req_port_o[109] = paddr_i[43];
  assign req_port_o[108] = paddr_i[42];
  assign req_port_o[107] = paddr_i[41];
  assign req_port_o[106] = paddr_i[40];
  assign req_port_o[105] = paddr_i[39];
  assign req_port_o[104] = paddr_i[38];
  assign req_port_o[103] = paddr_i[37];
  assign req_port_o[102] = paddr_i[36];
  assign req_port_o[101] = paddr_i[35];
  assign req_port_o[100] = paddr_i[34];
  assign req_port_o[99] = paddr_i[33];
  assign req_port_o[98] = paddr_i[32];
  assign req_port_o[97] = paddr_i[31];
  assign req_port_o[96] = paddr_i[30];
  assign req_port_o[95] = paddr_i[29];
  assign req_port_o[94] = paddr_i[28];
  assign req_port_o[93] = paddr_i[27];
  assign req_port_o[92] = paddr_i[26];
  assign req_port_o[91] = paddr_i[25];
  assign req_port_o[90] = paddr_i[24];
  assign req_port_o[89] = paddr_i[23];
  assign req_port_o[88] = paddr_i[22];
  assign req_port_o[87] = paddr_i[21];
  assign req_port_o[86] = paddr_i[20];
  assign req_port_o[85] = paddr_i[19];
  assign req_port_o[84] = paddr_i[18];
  assign req_port_o[83] = paddr_i[17];
  assign req_port_o[82] = paddr_i[16];
  assign req_port_o[81] = paddr_i[15];
  assign req_port_o[80] = paddr_i[14];
  assign req_port_o[79] = paddr_i[13];
  assign req_port_o[78] = paddr_i[12];
  assign N41 = lsu_ctrl_i[9] | N122;
  assign N42 = lsu_ctrl_i[7] | lsu_ctrl_i[6];
  assign N43 = lsu_ctrl_i[5] | N127;
  assign N44 = N41 | N42;
  assign N45 = N43 | lsu_ctrl_i[3];
  assign N46 = N44 | N45;
  assign N48 = N43 | N47;
  assign N49 = N44 | N48;
  assign N50 = N125 | lsu_ctrl_i[8];
  assign N51 = N113 | lsu_ctrl_i[6];
  assign N52 = lsu_ctrl_i[5] | lsu_ctrl_i[4];
  assign N53 = N50 | N51;
  assign N54 = N52 | lsu_ctrl_i[3];
  assign N55 = N53 | N54;
  assign N57 = N56 | lsu_ctrl_i[4];
  assign N58 = N57 | lsu_ctrl_i[3];
  assign N59 = N53 | N58;
  assign N61 = lsu_ctrl_i[7] | N60;
  assign N62 = N56 | N127;
  assign N63 = N41 | N61;
  assign N64 = N62 | lsu_ctrl_i[3];
  assign N65 = N63 | N64;
  assign N66 = N41 | N51;
  assign N67 = N66 | N54;
  assign N68 = N113 | N60;
  assign N69 = N41 | N68;
  assign N70 = N69 | N45;
  assign N71 = N69 | N48;
  assign N72 = N69 | N58;
  assign N73 = N57 | N47;
  assign N74 = N69 | N73;
  assign N75 = N69 | N64;
  assign N76 = N62 | N47;
  assign N77 = N69 | N76;
  assign N78 = N50 | N42;
  assign N79 = N78 | N54;
  assign N80 = N52 | N47;
  assign N81 = N78 | N80;
  assign N82 = N78 | N45;
  assign N84 = N44 | N58;
  assign N85 = N44 | N73;
  assign N86 = N44 | N64;
  assign N87 = N53 | N80;
  assign N88 = N53 | N73;
  assign N89 = N63 | N73;
  assign N90 = N63 | N76;
  assign N91 = N66 | N80;
  assign N92 = N66 | N45;
  assign N93 = N66 | N48;
  assign N94 = N66 | N58;
  assign N95 = N66 | N73;
  assign N96 = N66 | N64;
  assign N97 = N66 | N76;
  assign N98 = N69 | N54;
  assign N99 = N69 | N80;
  assign N101 = N44 | N76;
  assign N102 = N63 | N54;
  assign N103 = N63 | N80;
  assign N104 = N53 | N45;
  assign N105 = N53 | N64;
  assign N107 = N63 | N45;
  assign N108 = N63 | N58;
  assign N109 = N63 | N48;
  assign N110 = N53 | N48;
  assign N111 = N53 | N76;
  assign N114 = lsu_ctrl_i[9] & N113;
  assign N115 = lsu_ctrl_i[4] & lsu_ctrl_i[3];
  assign N116 = N114 & N115;
  assign N117 = N122 & N113;
  assign N118 = N117 & N115;
  assign N119 = N114 & lsu_ctrl_i[5];
  assign N120 = N117 & lsu_ctrl_i[5];
  assign N121 = lsu_ctrl_i[9] & lsu_ctrl_i[6];
  assign N123 = N122 & lsu_ctrl_i[6];
  assign N124 = lsu_ctrl_i[9] & lsu_ctrl_i[8];
  assign N126 = N125 & N122;
  assign N128 = N125 & N113;
  assign N129 = N60 & N56;
  assign N130 = N128 & N129;
  assign N131 = N130 & N127;
  assign N132 = lsu_ctrl_i[8] & N113;
  assign N133 = N132 & N129;
  assign N134 = N133 & N127;
  assign N136 = N372 & N377;
  assign N137 = N136 & N373;
  assign N138 = state_q[2] | N377;
  assign N139 = N138 | N373;
  assign N141 = N372 | state_q[1];
  assign N142 = N141 | state_q[0];
  assign N144 = N372 | state_q[1];
  assign N145 = N144 | N373;
  assign N147 = state_q[2] | state_q[1];
  assign N148 = N147 | N373;
  assign N150 = state_q[2] | N377;
  assign N151 = N150 | state_q[0];
  assign N153 = N372 | N377;
  assign N154 = N153 | state_q[0];

  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[12] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[12] <= load_data_d[12];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[11] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[11] <= load_data_d[11];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[10] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[10] <= load_data_d[10];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[9] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[9] <= load_data_d[9];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[8] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[8] <= load_data_d[8];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[7] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[7] <= load_data_d[7];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[6] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[6] <= load_data_d[6];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[5] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[5] <= load_data_d[5];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[4] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[4] <= load_data_d[4];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[3] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[3] <= load_data_d[3];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[2] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[2] <= load_data_d[2];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[1] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[1] <= load_data_d[1];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      load_data_q[0] <= 1'b0;
    end else if(1'b1) begin
      load_data_q[0] <= load_data_d[0];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      state_q[2] <= 1'b0;
    end else if(N371) begin
      state_q[2] <= state_d[2];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      state_q[1] <= 1'b0;
    end else if(N371) begin
      state_q[1] <= state_d[1];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      state_q[0] <= 1'b0;
    end else if(N371) begin
      state_q[0] <= state_d[0];
    end 
  end

  assign { shifted_data, result_o[7:0] } = req_port_i[63:0] >> { load_data_q[9:7], 1'b0, 1'b0, 1'b0 };
  assign N212 = load_data_d[6] | N211;
  assign N213 = N212 | load_data_d[4];
  assign N216 = load_data_d[3] | N215;
  assign N217 = load_data_d[1] | load_data_d[0];
  assign N218 = N216 | N217;
  assign N221 = load_data_d[3] | N215;
  assign N222 = N219 | N220;
  assign N223 = N221 | N222;
  assign N225 = N224 | load_data_d[2];
  assign N226 = N219 | load_data_d[0];
  assign N227 = N225 | N226;
  assign N231 = N229 | load_data_d[5];
  assign N232 = N230 | load_data_d[3];
  assign N233 = N231 | N232;
  assign N234 = N233 | load_data_d[2];
  assign N236 = load_data_d[1] | N220;
  assign N237 = N219 | load_data_d[0];
  assign N238 = load_data_d[1] & load_data_d[0];
  assign N240 = N224 & N219;
  assign N241 = load_data_d[6] | N211;
  assign N242 = load_data_d[4] | N215;
  assign N243 = N241 | N242;
  assign N244 = N243 | load_data_d[0];
  assign N245 = N229 | load_data_d[5];
  assign N246 = N230 | load_data_d[2];
  assign N247 = N245 | N246;
  assign N248 = N247 | N220;
  assign N253 = N224 & load_data_d[1];
  assign N254 = load_data_d[6] | N211;
  assign N255 = load_data_d[4] | N215;
  assign N256 = N254 | N255;
  assign N257 = N256 | N220;
  assign N258 = N229 | load_data_d[5];
  assign N259 = N230 | load_data_d[2];
  assign N260 = N258 | N259;
  assign N261 = N260 | load_data_d[0];

  always @(N264 or N252) begin
    if(N252) begin
      n__tmp493 <= N264;
    end 
  end

  assign N291 = (N283)? req_port_i[7] : 
                (N285)? req_port_i[15] : 
                (N287)? req_port_i[23] : 
                (N289)? req_port_i[31] : 
                (N284)? req_port_i[39] : 
                (N286)? req_port_i[47] : 
                (N288)? req_port_i[55] : 
                (N290)? req_port_i[63] : 1'b0;
  assign N294 = load_data_q[6] | N292;
  assign N295 = load_data_q[4] | load_data_q[3];
  assign N296 = N293 | load_data_q[1];
  assign N297 = N294 | N295;
  assign N298 = N296 | load_data_q[0];
  assign N299 = N297 | N298;
  assign N301 = load_data_q[6] | N292;
  assign N302 = load_data_q[4] | load_data_q[3];
  assign N303 = N293 | load_data_q[1];
  assign N304 = N301 | N302;
  assign N305 = N303 | N300;
  assign N306 = N304 | N305;
  assign N309 = N307 | load_data_q[5];
  assign N310 = N308 | load_data_q[3];
  assign N311 = load_data_q[2] | load_data_q[1];
  assign N312 = N309 | N310;
  assign N313 = N311 | N300;
  assign N314 = N312 | N313;
  assign N317 = load_data_q[6] | N292;
  assign N318 = load_data_q[4] | load_data_q[3];
  assign N319 = N293 | N316;
  assign N320 = N317 | N318;
  assign N321 = N319 | N300;
  assign N322 = N320 | N321;
  assign N324 = load_data_q[6] | N292;
  assign N325 = load_data_q[4] | N323;
  assign N326 = load_data_q[2] | load_data_q[1];
  assign N327 = N324 | N325;
  assign N328 = N326 | load_data_q[0];
  assign N329 = N327 | N328;
  assign N330 = N307 | load_data_q[5];
  assign N331 = N308 | load_data_q[3];
  assign N332 = load_data_q[2] | N316;
  assign N333 = N330 | N331;
  assign N334 = N332 | load_data_q[0];
  assign N335 = N333 | N334;
  assign N337 = load_data_q[6] | N292;
  assign N338 = load_data_q[4] | N323;
  assign N339 = load_data_q[2] | N316;
  assign N340 = N337 | N338;
  assign N341 = N339 | load_data_q[0];
  assign N342 = N340 | N341;
  assign N343 = load_data_q[6] | N292;
  assign N344 = load_data_q[4] | N323;
  assign N345 = N293 | load_data_q[1];
  assign N346 = N343 | N344;
  assign N347 = N345 | load_data_q[0];
  assign N348 = N346 | N347;
  assign N349 = N307 | load_data_q[5];
  assign N350 = N308 | load_data_q[3];
  assign N351 = load_data_q[2] | N316;
  assign N352 = N349 | N350;
  assign N353 = N351 | N300;
  assign N354 = N352 | N353;

  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      signed_q <= 1'b0;
    end else if(1'b1) begin
      signed_q <= signed_d;
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      fp_sign_q <= 1'b0;
    end else if(1'b1) begin
      fp_sign_q <= fp_sign_d;
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      idx_q[2] <= 1'b0;
    end else if(1'b1) begin
      idx_q[2] <= idx_d[2];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      idx_q[1] <= 1'b0;
    end else if(1'b1) begin
      idx_q[1] <= idx_d[1];
    end 
  end


  always @(posedge clk_i or posedge N210) begin
    if(N210) begin
      idx_q[0] <= 1'b0;
    end else if(1'b1) begin
      idx_q[0] <= idx_d[0];
    end 
  end

  assign N372 = ~state_q[2];
  assign N373 = ~state_q[0];
  assign N374 = state_q[1] | N372;
  assign N375 = N373 | N374;
  assign N376 = ~N375;
  assign N377 = ~state_q[1];
  assign N378 = N377 | N372;
  assign N379 = state_q[0] | N378;
  assign { N269, N268, N267 } = load_data_d[9:7] + { 1'b1, 1'b1 };
  assign { N273, N272, N271 } = load_data_d[9:7] + 1'b1;
  assign req_port_o[3:2] = (N0)? { 1'b1, 1'b1 } : 
                           (N1)? { 1'b1, 1'b0 } : 
                           (N2)? { 1'b0, 1'b1 } : 
                           (N3)? { 1'b0, 1'b0 } : 
                           (N4)? { 1'b1, 1'b1 } : 1'b0;
  assign N0 = N83;
  assign N1 = N100;
  assign N2 = N106;
  assign N3 = N112;
  assign N4 = N135;
  assign { N160, N159, N158 } = (N5)? { 1'b0, 1'b0, 1'b1 } : 
                                (N170)? { 1'b0, 1'b1, 1'b0 } : 
                                (N6)? { 1'b1, 1'b0, 1'b0 } : 1'b0;
  assign N5 = N39;
  assign N6 = N171;
  assign N161 = (N7)? N159 : 
                (N8)? 1'b0 : 1'b0;
  assign N7 = N40;
  assign N8 = page_offset_matches_i;
  assign { N164, N163, N162 } = (N7)? { N160, N159, N158 } : 
                                (N8)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign N165 = (N9)? N40 : 
                (N10)? 1'b0 : 1'b0;
  assign N9 = valid_i;
  assign N10 = N156;
  assign N166 = (N9)? N161 : 
                (N10)? 1'b0 : 1'b0;
  assign N169 = (N11)? dtlb_hit_i : 
                (N168)? 1'b0 : 1'b0;
  assign N11 = req_port_i[65];
  assign N171 = ~N157;
  assign { N174, N173, N172 } = (N7)? { N171, N170, N39 } : 
                                (N8)? { 1'b0, 1'b1, 1'b1 } : 1'b0;
  assign { N177, N176, N175 } = (N9)? { N174, N173, N172 } : 
                                (N10)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N185 = (N12)? N166 : 
                (N13)? 1'b0 : 
                (N14)? 1'b0 : 
                (N15)? 1'b0 : 
                (N16)? N169 : 
                (N17)? N166 : 
                (N18)? 1'b0 : 
                (N184)? 1'b0 : 1'b0;
  assign N12 = N137;
  assign N13 = N140;
  assign N14 = N143;
  assign N15 = N146;
  assign N16 = N149;
  assign N17 = N152;
  assign N18 = N155;
  assign translation_req_o = (N12)? valid_i : 
                             (N13)? 1'b0 : 
                             (N14)? 1'b0 : 
                             (N15)? 1'b1 : 
                             (N16)? 1'b1 : 
                             (N17)? valid_i : 
                             (N18)? 1'b0 : 
                             (N184)? 1'b0 : 1'b0;
  assign { N188, N187, N186 } = (N12)? { N164, N163, N162 } : 
                                (N13)? { 1'b0, 1'b0, 1'b1 } : 
                                (N14)? { 1'b1, 1'b0, 1'b1 } : 
                                (N15)? { 1'b0, 1'b0, 1'b1 } : 
                                (N16)? { N167, dtlb_hit_i, 1'b0 } : 
                                (N17)? { N177, N176, N175 } : 
                                (N18)? { 1'b0, 1'b0, 1'b0 } : 
                                (N184)? state_q : 1'b0;
  assign { req_port_o[13:13], req_port_o[1:0] } = (N12)? { N165, 1'b0, 1'b0 } : 
                                                  (N13)? { 1'b0, 1'b0, 1'b0 } : 
                                                  (N14)? { 1'b0, 1'b1, 1'b1 } : 
                                                  (N15)? { 1'b0, 1'b0, 1'b0 } : 
                                                  (N16)? { 1'b1, 1'b0, 1'b0 } : 
                                                  (N17)? { N165, ex_i[0:0], 1'b1 } : 
                                                  (N18)? { 1'b0, 1'b1, 1'b1 } : 
                                                  (N184)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N192 = (N19)? 1'b1 : 
                (N20)? N185 : 1'b0;
  assign N19 = N191;
  assign N20 = req_port_i[64];
  assign { N195, N194, N193 } = (N21)? { 1'b0, 1'b0, 1'b0 } : 
                                (N190)? { N188, N187, N186 } : 1'b0;
  assign N21 = N189;
  assign pop_ld_o = (N21)? N192 : 
                    (N190)? N185 : 1'b0;
  assign load_data_d = (N22)? { lsu_ctrl_i[2:0], lsu_ctrl_i[88:86], lsu_ctrl_i[9:3] } : 
                       (N197)? load_data_q : 1'b0;
  assign N22 = N196;
  assign state_d = (N23)? { 1'b1, 1'b1, 1'b0 } : 
                   (N24)? { N195, N194, N193 } : 1'b0;
  assign N23 = flush_i;
  assign N24 = N198;
  assign N203 = (N25)? 1'b1 : 
                (N202)? N201 : 1'b0;
  assign N25 = ex_i[0];
  assign N204 = (N26)? N203 : 
                (N200)? 1'b0 : 1'b0;
  assign N26 = N199;
  assign valid_o = (N27)? 1'b1 : 
                   (N209)? 1'b0 : 
                   (N207)? N204 : 1'b0;
  assign N27 = N205;
  assign trans_id_o = (N27)? lsu_ctrl_i[2:0] : 
                      (N208)? load_data_q[12:10] : 
                      (N28)? load_data_q[12:10] : 1'b0;
  assign N28 = 1'b0;
  assign signed_d = (N29)? N228 : 
                    (N30)? 1'b0 : 1'b0;
  assign N29 = N214;
  assign N30 = N213;
  assign fp_sign_d = (N31)? N239 : 
                     (N32)? 1'b0 : 1'b0;
  assign N31 = N235;
  assign N32 = N234;
  assign N251 = (N33)? N249 : 
                (N250)? 1'b0 : 1'b0;
  assign N33 = N240;
  assign N264 = (N34)? N262 : 
                (N263)? 1'b0 : 1'b0;
  assign N34 = N253;
  assign idx_d = (N35)? { N269, N268, N267 } : 
                 (N275)? { N273, N272, N271 } : 
                 (N266)? load_data_d[9:7] : 1'b0;
  assign N35 = N251;
  assign result_o[63:8] = (N36)? { sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, shifted_data[31:8] } : 
                          (N37)? { sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, shifted_data[15:8] } : 
                          (N38)? { sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit, sign_bit } : 
                          (N358)? shifted_data : 1'b0;
  assign N36 = N315;
  assign N37 = N336;
  assign N38 = N355;
  assign N39 = ~req_port_i[65];
  assign N40 = ~page_offset_matches_i;
  assign N47 = ~lsu_ctrl_i[3];
  assign N56 = ~lsu_ctrl_i[5];
  assign N60 = ~lsu_ctrl_i[6];
  assign N83 = N406 | N407;
  assign N406 = N404 | N405;
  assign N404 = N402 | N403;
  assign N402 = N400 | N401;
  assign N400 = N398 | N399;
  assign N398 = N396 | N397;
  assign N396 = N394 | N395;
  assign N394 = N392 | N393;
  assign N392 = N390 | N391;
  assign N390 = N388 | N389;
  assign N388 = N386 | N387;
  assign N386 = N384 | N385;
  assign N384 = N382 | N383;
  assign N382 = N380 | N381;
  assign N380 = ~N46;
  assign N381 = ~N49;
  assign N383 = ~N55;
  assign N385 = ~N59;
  assign N387 = ~N65;
  assign N389 = ~N67;
  assign N391 = ~N70;
  assign N393 = ~N71;
  assign N395 = ~N72;
  assign N397 = ~N74;
  assign N399 = ~N75;
  assign N401 = ~N77;
  assign N403 = ~N79;
  assign N405 = ~N81;
  assign N407 = ~N82;
  assign N100 = N436 | N437;
  assign N436 = N434 | N435;
  assign N434 = N432 | N433;
  assign N432 = N430 | N431;
  assign N430 = N428 | N429;
  assign N428 = N426 | N427;
  assign N426 = N424 | N425;
  assign N424 = N422 | N423;
  assign N422 = N420 | N421;
  assign N420 = N418 | N419;
  assign N418 = N416 | N417;
  assign N416 = N414 | N415;
  assign N414 = N412 | N413;
  assign N412 = N410 | N411;
  assign N410 = N408 | N409;
  assign N408 = ~N84;
  assign N409 = ~N85;
  assign N411 = ~N86;
  assign N413 = ~N87;
  assign N415 = ~N88;
  assign N417 = ~N89;
  assign N419 = ~N90;
  assign N421 = ~N91;
  assign N423 = ~N92;
  assign N425 = ~N93;
  assign N427 = ~N94;
  assign N429 = ~N95;
  assign N431 = ~N96;
  assign N433 = ~N97;
  assign N435 = ~N98;
  assign N437 = ~N99;
  assign N106 = N444 | N445;
  assign N444 = N442 | N443;
  assign N442 = N440 | N441;
  assign N440 = N438 | N439;
  assign N438 = ~N101;
  assign N439 = ~N102;
  assign N441 = ~N103;
  assign N443 = ~N104;
  assign N445 = ~N105;
  assign N112 = N452 | N453;
  assign N452 = N450 | N451;
  assign N450 = N448 | N449;
  assign N448 = N446 | N447;
  assign N446 = ~N107;
  assign N447 = ~N108;
  assign N449 = ~N109;
  assign N451 = ~N110;
  assign N453 = ~N111;
  assign N113 = ~lsu_ctrl_i[7];
  assign N122 = ~lsu_ctrl_i[8];
  assign N125 = ~lsu_ctrl_i[9];
  assign N127 = ~lsu_ctrl_i[4];
  assign N135 = N116 | N461;
  assign N461 = N118 | N460;
  assign N460 = N119 | N459;
  assign N459 = N120 | N458;
  assign N458 = N121 | N457;
  assign N457 = N123 | N456;
  assign N456 = N124 | N455;
  assign N455 = N126 | N454;
  assign N454 = N131 | N134;
  assign N140 = ~N139;
  assign N143 = ~N142;
  assign N146 = ~N145;
  assign N149 = ~N148;
  assign N152 = ~N151;
  assign N155 = ~N154;
  assign N156 = ~valid_i;
  assign N157 = dtlb_hit_i | N39;
  assign N167 = ~dtlb_hit_i;
  assign N168 = ~req_port_i[65];
  assign N178 = N140 | N137;
  assign N179 = N143 | N178;
  assign N180 = N146 | N179;
  assign N181 = N149 | N180;
  assign N182 = N152 | N181;
  assign N183 = N155 | N182;
  assign N184 = ~N183;
  assign N189 = ex_i[0] & valid_i;
  assign N190 = ~N189;
  assign N191 = ~req_port_i[64];
  assign N196 = pop_ld_o & N462;
  assign N462 = ~ex_i[0];
  assign N197 = ~N196;
  assign N198 = ~flush_i;
  assign N170 = dtlb_hit_i & req_port_i[65];
  assign N199 = req_port_i[64] & N379;
  assign N200 = ~N199;
  assign N201 = ~req_port_o[1];
  assign N202 = ~ex_i[0];
  assign N205 = N463 & N191;
  assign N463 = valid_i & ex_i[0];
  assign N206 = N376 | N205;
  assign N207 = ~N206;
  assign N208 = ~N205;
  assign N209 = N376 & N208;
  assign N210 = ~rst_ni;
  assign N211 = ~load_data_d[5];
  assign N214 = ~N213;
  assign N215 = ~load_data_d[2];
  assign N219 = ~load_data_d[1];
  assign N220 = ~load_data_d[0];
  assign N224 = ~load_data_d[3];
  assign N228 = N466 | N467;
  assign N466 = N464 | N465;
  assign N464 = ~N218;
  assign N465 = ~N223;
  assign N467 = ~N227;
  assign N229 = ~load_data_d[6];
  assign N230 = ~load_data_d[4];
  assign N235 = ~N234;
  assign N239 = N470 | N238;
  assign N470 = N468 | N469;
  assign N468 = ~N236;
  assign N469 = ~N237;
  assign N249 = N471 | N472;
  assign N471 = ~N244;
  assign N472 = ~N248;
  assign N250 = ~N240;
  assign N252 = ~N251;
  assign N262 = N473 | N474;
  assign N473 = ~N257;
  assign N474 = ~N261;
  assign N263 = ~N253;
  assign N265 = n__tmp493 | N251;
  assign N266 = ~N265;
  assign N270 = N275;
  assign N274 = ~N251;
  assign N275 = n__tmp493 & N274;
  assign N276 = ~idx_q[0];
  assign N277 = ~idx_q[1];
  assign N278 = N276 & N277;
  assign N279 = N276 & idx_q[1];
  assign N280 = idx_q[0] & N277;
  assign N281 = idx_q[0] & idx_q[1];
  assign N282 = ~idx_q[2];
  assign N283 = N278 & N282;
  assign N284 = N278 & idx_q[2];
  assign N285 = N280 & N282;
  assign N286 = N280 & idx_q[2];
  assign N287 = N279 & N282;
  assign N288 = N279 & idx_q[2];
  assign N289 = N281 & N282;
  assign N290 = N281 & idx_q[2];
  assign sign_bit = N475 | fp_sign_q;
  assign N475 = signed_q & N291;
  assign N292 = ~load_data_q[5];
  assign N293 = ~load_data_q[2];
  assign N300 = ~load_data_q[0];
  assign N307 = ~load_data_q[6];
  assign N308 = ~load_data_q[4];
  assign N315 = N478 | N479;
  assign N478 = N476 | N477;
  assign N476 = ~N299;
  assign N477 = ~N306;
  assign N479 = ~N314;
  assign N316 = ~load_data_q[1];
  assign N323 = ~load_data_q[3];
  assign N336 = N482 | N483;
  assign N482 = N480 | N481;
  assign N480 = ~N322;
  assign N481 = ~N329;
  assign N483 = ~N335;
  assign N355 = N486 | N487;
  assign N486 = N484 | N485;
  assign N484 = ~N342;
  assign N485 = ~N348;
  assign N487 = ~N354;
  assign N356 = N336 | N315;
  assign N357 = N355 | N356;
  assign N358 = ~N357;
  assign N359 = N190 & N198;
  assign N360 = N137 & N359;
  assign N361 = N156 & N360;
  assign N362 = N140 & N359;
  assign N363 = page_offset_matches_i & N362;
  assign N364 = N361 | N363;
  assign N365 = N146 & N359;
  assign N366 = N167 & N365;
  assign N367 = N364 | N366;
  assign N368 = N149 & N359;
  assign N369 = N168 & N368;
  assign N370 = N367 | N369;
  assign N371 = ~N370;

endmodule