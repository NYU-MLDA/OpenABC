module MulAddRecFN_postMul_1
(
  io_fromPreMul_highExpA,
  io_fromPreMul_isNaN_isQuietNaNA,
  io_fromPreMul_highExpB,
  io_fromPreMul_isNaN_isQuietNaNB,
  io_fromPreMul_signProd,
  io_fromPreMul_isZeroProd,
  io_fromPreMul_opSignC,
  io_fromPreMul_highExpC,
  io_fromPreMul_isNaN_isQuietNaNC,
  io_fromPreMul_isCDominant,
  io_fromPreMul_CAlignDist_0,
  io_fromPreMul_CAlignDist,
  io_fromPreMul_bit0AlignedNegSigC,
  io_fromPreMul_highAlignedNegSigC,
  io_fromPreMul_sExpSum,
  io_fromPreMul_roundingMode,
  io_mulAddResult,
  io_out,
  io_exceptionFlags
);

  input [2:0] io_fromPreMul_highExpA;
  input [2:0] io_fromPreMul_highExpB;
  input [2:0] io_fromPreMul_highExpC;
  input [7:0] io_fromPreMul_CAlignDist;
  input [54:0] io_fromPreMul_highAlignedNegSigC;
  input [13:0] io_fromPreMul_sExpSum;
  input [1:0] io_fromPreMul_roundingMode;
  input [106:0] io_mulAddResult;
  output [64:0] io_out;
  output [4:0] io_exceptionFlags;
  input io_fromPreMul_isNaN_isQuietNaNA;
  input io_fromPreMul_isNaN_isQuietNaNB;
  input io_fromPreMul_signProd;
  input io_fromPreMul_isZeroProd;
  input io_fromPreMul_opSignC;
  input io_fromPreMul_isNaN_isQuietNaNC;
  input io_fromPreMul_isCDominant;
  input io_fromPreMul_CAlignDist_0;
  input io_fromPreMul_bit0AlignedNegSigC;
  wire [64:0] io_out,T261;
  wire [4:0] io_exceptionFlags,T525,T526,T527,T528,T529,T530,T531,T532,T533,T534,T535,T536,
  T537,T538,T539,T540,normTo2ShiftDist;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,T3,commonCase,inexactY,doIncrSig,N250,T287,anyRound,
  sigX3_56,T104_0,T9_0,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,
  N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
  N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,
  N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,
  N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,
  N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
  N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,T36,N358,
  T49_13,T49_11,T49_9,T49_7,T49_5,T49_3,T49_1,T50_12,T50_10,T50_8,T50_6,T50_4,T50_2,
  T53_11,T53_10,T53_7,T53_6,T53_3,T53_2,T54_9,T54_8,T54_5,T54_4,T57_7,T57_6,T57_5,
  T57_4,T74_29,T74_27,T74_25,T74_23,T74_21,T74_19,T74_17,T74_15,T74_13,T74_11,
  T74_9,T74_7,T74_5,T74_3,T74_1,T75_28,T75_26,T75_24,T75_22,T75_20,T75_18,T75_16,
  T75_14,T75_12,T75_10,T75_8,T75_6,T75_4,T75_2,T78_27,T78_26,T78_23,T78_22,T78_19,
  T78_18,T78_15,T78_14,T78_11,T78_10,T78_7,T78_6,T78_3,T78_2,T79_25,T79_24,T79_21,
  T79_20,T79_17,T79_16,T79_13,T79_12,T79_9,T79_8,T79_5,T79_4,T82_23,T82_22,T82_21,
  T82_20,T82_15,T82_14,T82_13,T82_12,T82_7,T82_6,T82_5,T82_4,T83_19,T83_18,T83_17,
  T83_16,T83_11,T83_10,T83_9,T83_8,T86_15,T86_14,T86_13,T86_12,T86_11,T86_10,T86_9,
  T86_8,absSigSumExtraMask_1,T136_5,T136_3,T136_1,T137_4,T137_2,T140_3,T140_2,T155_13,
  T155_11,T155_9,T155_7,T155_5,T155_3,T155_1,T156_12,T156_10,T156_8,T156_6,T156_4,
  T156_2,T159_11,T159_10,T159_7,T159_6,T159_3,T159_2,T160_9,T160_8,T160_5,T160_4,
  T163_7,T163_6,T163_5,T163_4,N359,N360,N361,T182_0,N362,T186_0,N363,T196,T213_0,
  T224,T233,T235,T243,T246,T252,T256,T254,T261_87,T261_86,allRound,T291,T293,T292,
  T295,T294,notSpecial_addZeros,addSpecial,mulSpecial,underflowY,T299,T300,
  sigX3Shift1,N364,roundEven,N365,T319,T316,T318,T317,T320,T321,T324,N366,T331,T325,
  roundDirectUp,signY,N367,isZeroY,N368,T327,doNegSignSum,N369,T328,T329,T334,T332,T333,
  T336,T335,T340,T337,T338,T339,T341,T342,T343,T348,N370,T351,T350,N371,N372,T377,
  notSigNaN_invalid,T374,T359,T360,T363,isInfC,T361,T369,T364,isInfA,isInfB,T365,
  T367,T372,T370,isNaNB,isNaNA,T376,T375,T380,isSigNaNC,isNaNC,T378,isSigNaNA,
  isSigNaNB,T381,T382,T385_0,T386,overflowY_roundMagUp,roundMagUp,T389,T387,T388,T392,
  T393,T397,N373,T398,totalUnderflowY,T403,T399,T400,notNaN_isInfOut,T408,T407,T409,
  pegMinFiniteMagOut,T414,notSpecial_isZeroOut,T427,T429,T428,T444,
  uncommonCaseSignOut,T434,T430,T431,T432,T433,T438,T435,T436,T437,T442,T439,T440,T441,T443,N374,
  N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,
  N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,
  N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,
  N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,
  N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,
  N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,
  N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,
  N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,
  N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,
  N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,
  N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,
  N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,
  N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,
  N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,
  N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,
  N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,
  N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,
  N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,
  N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,
  N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,
  N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,
  N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,
  N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
  N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,
  N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,
  N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,
  N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,
  N807,N808,N809,N810,N811,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,
  SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,
  SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11,SV2V_UNCONNECTED_12,
  SV2V_UNCONNECTED_13,SV2V_UNCONNECTED_14,SV2V_UNCONNECTED_15,SV2V_UNCONNECTED_16,
  SV2V_UNCONNECTED_17,SV2V_UNCONNECTED_18,SV2V_UNCONNECTED_19,
  SV2V_UNCONNECTED_20,SV2V_UNCONNECTED_21,SV2V_UNCONNECTED_22,
  SV2V_UNCONNECTED_23,SV2V_UNCONNECTED_24,SV2V_UNCONNECTED_25,SV2V_UNCONNECTED_26,
  SV2V_UNCONNECTED_27,SV2V_UNCONNECTED_28,SV2V_UNCONNECTED_29,
  SV2V_UNCONNECTED_30,SV2V_UNCONNECTED_31,SV2V_UNCONNECTED_32,
  SV2V_UNCONNECTED_33,SV2V_UNCONNECTED_34,SV2V_UNCONNECTED_35,SV2V_UNCONNECTED_36,
  SV2V_UNCONNECTED_37,SV2V_UNCONNECTED_38,SV2V_UNCONNECTED_39,
  SV2V_UNCONNECTED_40,SV2V_UNCONNECTED_41,SV2V_UNCONNECTED_42,
  SV2V_UNCONNECTED_43,SV2V_UNCONNECTED_44,SV2V_UNCONNECTED_45,SV2V_UNCONNECTED_46,
  SV2V_UNCONNECTED_47,SV2V_UNCONNECTED_48,SV2V_UNCONNECTED_49,
  SV2V_UNCONNECTED_50,SV2V_UNCONNECTED_51,SV2V_UNCONNECTED_52,
  SV2V_UNCONNECTED_53,SV2V_UNCONNECTED_54,SV2V_UNCONNECTED_55,SV2V_UNCONNECTED_56,
  SV2V_UNCONNECTED_57,SV2V_UNCONNECTED_58,SV2V_UNCONNECTED_59,
  SV2V_UNCONNECTED_60,SV2V_UNCONNECTED_61,SV2V_UNCONNECTED_62,
  SV2V_UNCONNECTED_63,SV2V_UNCONNECTED_64,SV2V_UNCONNECTED_65,SV2V_UNCONNECTED_66,
  SV2V_UNCONNECTED_67,SV2V_UNCONNECTED_68,SV2V_UNCONNECTED_69,
  SV2V_UNCONNECTED_70,SV2V_UNCONNECTED_71,SV2V_UNCONNECTED_72,
  SV2V_UNCONNECTED_73,SV2V_UNCONNECTED_74,SV2V_UNCONNECTED_75,SV2V_UNCONNECTED_76,
  SV2V_UNCONNECTED_77,SV2V_UNCONNECTED_78,SV2V_UNCONNECTED_79,
  SV2V_UNCONNECTED_80,SV2V_UNCONNECTED_81,SV2V_UNCONNECTED_82,
  SV2V_UNCONNECTED_83,SV2V_UNCONNECTED_84,SV2V_UNCONNECTED_85,SV2V_UNCONNECTED_86,
  SV2V_UNCONNECTED_87,SV2V_UNCONNECTED_88,SV2V_UNCONNECTED_89,
  SV2V_UNCONNECTED_90,SV2V_UNCONNECTED_91,SV2V_UNCONNECTED_92,
  SV2V_UNCONNECTED_93,SV2V_UNCONNECTED_94,SV2V_UNCONNECTED_95,SV2V_UNCONNECTED_96,
  SV2V_UNCONNECTED_97,SV2V_UNCONNECTED_98,SV2V_UNCONNECTED_99,
  SV2V_UNCONNECTED_100,SV2V_UNCONNECTED_101,SV2V_UNCONNECTED_102,
  SV2V_UNCONNECTED_103,SV2V_UNCONNECTED_104,SV2V_UNCONNECTED_105,
  SV2V_UNCONNECTED_106,SV2V_UNCONNECTED_107,SV2V_UNCONNECTED_108,
  SV2V_UNCONNECTED_109,SV2V_UNCONNECTED_110,SV2V_UNCONNECTED_111,SV2V_UNCONNECTED_112,
  SV2V_UNCONNECTED_113,SV2V_UNCONNECTED_114,SV2V_UNCONNECTED_115,
  SV2V_UNCONNECTED_116,SV2V_UNCONNECTED_117,SV2V_UNCONNECTED_118,
  SV2V_UNCONNECTED_119,SV2V_UNCONNECTED_120,SV2V_UNCONNECTED_121,
  SV2V_UNCONNECTED_122,SV2V_UNCONNECTED_123,SV2V_UNCONNECTED_124,
  SV2V_UNCONNECTED_125,SV2V_UNCONNECTED_126,SV2V_UNCONNECTED_127,SV2V_UNCONNECTED_128,
  SV2V_UNCONNECTED_129,SV2V_UNCONNECTED_130,SV2V_UNCONNECTED_131,
  SV2V_UNCONNECTED_132,SV2V_UNCONNECTED_133,SV2V_UNCONNECTED_134,
  SV2V_UNCONNECTED_135,SV2V_UNCONNECTED_136,SV2V_UNCONNECTED_137,
  SV2V_UNCONNECTED_138,SV2V_UNCONNECTED_139,SV2V_UNCONNECTED_140,
  SV2V_UNCONNECTED_141,SV2V_UNCONNECTED_142,SV2V_UNCONNECTED_143,SV2V_UNCONNECTED_144,
  SV2V_UNCONNECTED_145,SV2V_UNCONNECTED_146,SV2V_UNCONNECTED_147,
  SV2V_UNCONNECTED_148,SV2V_UNCONNECTED_149,SV2V_UNCONNECTED_150,
  SV2V_UNCONNECTED_151,SV2V_UNCONNECTED_152,SV2V_UNCONNECTED_153,
  SV2V_UNCONNECTED_154,SV2V_UNCONNECTED_155,SV2V_UNCONNECTED_156,
  SV2V_UNCONNECTED_157,SV2V_UNCONNECTED_158,SV2V_UNCONNECTED_159,SV2V_UNCONNECTED_160,
  SV2V_UNCONNECTED_161,SV2V_UNCONNECTED_162,SV2V_UNCONNECTED_163,
  SV2V_UNCONNECTED_164,SV2V_UNCONNECTED_165,SV2V_UNCONNECTED_166,
  SV2V_UNCONNECTED_167,SV2V_UNCONNECTED_168,SV2V_UNCONNECTED_169,
  SV2V_UNCONNECTED_170,SV2V_UNCONNECTED_171,SV2V_UNCONNECTED_172,
  SV2V_UNCONNECTED_173,SV2V_UNCONNECTED_174,SV2V_UNCONNECTED_175,SV2V_UNCONNECTED_176,
  SV2V_UNCONNECTED_177,SV2V_UNCONNECTED_178,SV2V_UNCONNECTED_179,
  SV2V_UNCONNECTED_180,SV2V_UNCONNECTED_181,SV2V_UNCONNECTED_182,
  SV2V_UNCONNECTED_183,SV2V_UNCONNECTED_184,SV2V_UNCONNECTED_185,
  SV2V_UNCONNECTED_186,SV2V_UNCONNECTED_187,SV2V_UNCONNECTED_188,
  SV2V_UNCONNECTED_189,SV2V_UNCONNECTED_190,SV2V_UNCONNECTED_191,SV2V_UNCONNECTED_192,
  SV2V_UNCONNECTED_193,SV2V_UNCONNECTED_194,SV2V_UNCONNECTED_195,
  SV2V_UNCONNECTED_196,SV2V_UNCONNECTED_197,SV2V_UNCONNECTED_198,
  SV2V_UNCONNECTED_199,SV2V_UNCONNECTED_200,SV2V_UNCONNECTED_201,
  SV2V_UNCONNECTED_202,SV2V_UNCONNECTED_203,SV2V_UNCONNECTED_204,
  SV2V_UNCONNECTED_205,SV2V_UNCONNECTED_206,SV2V_UNCONNECTED_207,SV2V_UNCONNECTED_208,
  SV2V_UNCONNECTED_209,SV2V_UNCONNECTED_210,SV2V_UNCONNECTED_211,
  SV2V_UNCONNECTED_212,SV2V_UNCONNECTED_213,SV2V_UNCONNECTED_214,
  SV2V_UNCONNECTED_215,SV2V_UNCONNECTED_216,SV2V_UNCONNECTED_217,
  SV2V_UNCONNECTED_218,SV2V_UNCONNECTED_219,SV2V_UNCONNECTED_220,
  SV2V_UNCONNECTED_221,SV2V_UNCONNECTED_222,SV2V_UNCONNECTED_223,SV2V_UNCONNECTED_224,
  SV2V_UNCONNECTED_225,SV2V_UNCONNECTED_226,SV2V_UNCONNECTED_227,
  SV2V_UNCONNECTED_228,SV2V_UNCONNECTED_229,SV2V_UNCONNECTED_230,
  SV2V_UNCONNECTED_231,SV2V_UNCONNECTED_232,SV2V_UNCONNECTED_233,
  SV2V_UNCONNECTED_234,SV2V_UNCONNECTED_235,SV2V_UNCONNECTED_236,
  SV2V_UNCONNECTED_237,SV2V_UNCONNECTED_238,SV2V_UNCONNECTED_239,SV2V_UNCONNECTED_240,
  SV2V_UNCONNECTED_241,SV2V_UNCONNECTED_242,SV2V_UNCONNECTED_243,
  SV2V_UNCONNECTED_244,SV2V_UNCONNECTED_245,SV2V_UNCONNECTED_246,
  SV2V_UNCONNECTED_247,SV2V_UNCONNECTED_248,SV2V_UNCONNECTED_249,
  SV2V_UNCONNECTED_250,SV2V_UNCONNECTED_251,SV2V_UNCONNECTED_252,
  SV2V_UNCONNECTED_253,SV2V_UNCONNECTED_254,SV2V_UNCONNECTED_255,SV2V_UNCONNECTED_256,
  SV2V_UNCONNECTED_257,SV2V_UNCONNECTED_258,SV2V_UNCONNECTED_259,
  SV2V_UNCONNECTED_260,SV2V_UNCONNECTED_261,SV2V_UNCONNECTED_262,
  SV2V_UNCONNECTED_263,SV2V_UNCONNECTED_264,SV2V_UNCONNECTED_265,
  SV2V_UNCONNECTED_266,SV2V_UNCONNECTED_267,SV2V_UNCONNECTED_268,
  SV2V_UNCONNECTED_269,SV2V_UNCONNECTED_270,SV2V_UNCONNECTED_271,SV2V_UNCONNECTED_272,
  SV2V_UNCONNECTED_273,SV2V_UNCONNECTED_274,SV2V_UNCONNECTED_275,
  SV2V_UNCONNECTED_276,SV2V_UNCONNECTED_277,SV2V_UNCONNECTED_278,
  SV2V_UNCONNECTED_279,SV2V_UNCONNECTED_280,SV2V_UNCONNECTED_281,
  SV2V_UNCONNECTED_282,SV2V_UNCONNECTED_283,SV2V_UNCONNECTED_284,
  SV2V_UNCONNECTED_285,SV2V_UNCONNECTED_286,SV2V_UNCONNECTED_287,SV2V_UNCONNECTED_288,
  SV2V_UNCONNECTED_289,SV2V_UNCONNECTED_290,SV2V_UNCONNECTED_291,
  SV2V_UNCONNECTED_292,SV2V_UNCONNECTED_293,SV2V_UNCONNECTED_294,
  SV2V_UNCONNECTED_295,SV2V_UNCONNECTED_296,SV2V_UNCONNECTED_297,
  SV2V_UNCONNECTED_298,SV2V_UNCONNECTED_299,SV2V_UNCONNECTED_300,
  SV2V_UNCONNECTED_301,SV2V_UNCONNECTED_302,SV2V_UNCONNECTED_303,SV2V_UNCONNECTED_304,
  SV2V_UNCONNECTED_305,SV2V_UNCONNECTED_306,SV2V_UNCONNECTED_307,
  SV2V_UNCONNECTED_308,SV2V_UNCONNECTED_309,SV2V_UNCONNECTED_310,
  SV2V_UNCONNECTED_311,SV2V_UNCONNECTED_312,SV2V_UNCONNECTED_313,
  SV2V_UNCONNECTED_314,SV2V_UNCONNECTED_315,SV2V_UNCONNECTED_316,
  SV2V_UNCONNECTED_317,SV2V_UNCONNECTED_318,SV2V_UNCONNECTED_319,SV2V_UNCONNECTED_320,
  SV2V_UNCONNECTED_321,SV2V_UNCONNECTED_322,SV2V_UNCONNECTED_323,
  SV2V_UNCONNECTED_324,SV2V_UNCONNECTED_325,SV2V_UNCONNECTED_326,
  SV2V_UNCONNECTED_327,SV2V_UNCONNECTED_328,SV2V_UNCONNECTED_329,
  SV2V_UNCONNECTED_330,SV2V_UNCONNECTED_331,SV2V_UNCONNECTED_332,
  SV2V_UNCONNECTED_333,SV2V_UNCONNECTED_334,SV2V_UNCONNECTED_335,SV2V_UNCONNECTED_336,
  SV2V_UNCONNECTED_337,SV2V_UNCONNECTED_338,SV2V_UNCONNECTED_339,
  SV2V_UNCONNECTED_340,SV2V_UNCONNECTED_341,SV2V_UNCONNECTED_342,
  SV2V_UNCONNECTED_343,SV2V_UNCONNECTED_344,SV2V_UNCONNECTED_345,
  SV2V_UNCONNECTED_346,SV2V_UNCONNECTED_347,SV2V_UNCONNECTED_348,
  SV2V_UNCONNECTED_349,SV2V_UNCONNECTED_350,SV2V_UNCONNECTED_351,SV2V_UNCONNECTED_352,
  SV2V_UNCONNECTED_353,SV2V_UNCONNECTED_354,SV2V_UNCONNECTED_355,
  SV2V_UNCONNECTED_356,SV2V_UNCONNECTED_357,SV2V_UNCONNECTED_358,
  SV2V_UNCONNECTED_359,SV2V_UNCONNECTED_360,SV2V_UNCONNECTED_361,
  SV2V_UNCONNECTED_362,SV2V_UNCONNECTED_363,SV2V_UNCONNECTED_364,
  SV2V_UNCONNECTED_365,SV2V_UNCONNECTED_366,SV2V_UNCONNECTED_367,SV2V_UNCONNECTED_368,
  SV2V_UNCONNECTED_369,SV2V_UNCONNECTED_370,SV2V_UNCONNECTED_371,
  SV2V_UNCONNECTED_372,SV2V_UNCONNECTED_373,SV2V_UNCONNECTED_374,
  SV2V_UNCONNECTED_375,SV2V_UNCONNECTED_376,SV2V_UNCONNECTED_377,
  SV2V_UNCONNECTED_378,SV2V_UNCONNECTED_379,SV2V_UNCONNECTED_380,
  SV2V_UNCONNECTED_381,SV2V_UNCONNECTED_382,SV2V_UNCONNECTED_383,SV2V_UNCONNECTED_384,
  SV2V_UNCONNECTED_385,SV2V_UNCONNECTED_386,SV2V_UNCONNECTED_387,
  SV2V_UNCONNECTED_388,SV2V_UNCONNECTED_389,SV2V_UNCONNECTED_390,
  SV2V_UNCONNECTED_391,SV2V_UNCONNECTED_392,SV2V_UNCONNECTED_393,
  SV2V_UNCONNECTED_394,SV2V_UNCONNECTED_395,SV2V_UNCONNECTED_396,
  SV2V_UNCONNECTED_397,SV2V_UNCONNECTED_398,SV2V_UNCONNECTED_399,SV2V_UNCONNECTED_400,
  SV2V_UNCONNECTED_401,SV2V_UNCONNECTED_402,SV2V_UNCONNECTED_403,
  SV2V_UNCONNECTED_404,SV2V_UNCONNECTED_405,SV2V_UNCONNECTED_406,
  SV2V_UNCONNECTED_407,SV2V_UNCONNECTED_408,SV2V_UNCONNECTED_409,
  SV2V_UNCONNECTED_410,SV2V_UNCONNECTED_411,SV2V_UNCONNECTED_412,
  SV2V_UNCONNECTED_413,SV2V_UNCONNECTED_414,SV2V_UNCONNECTED_415,SV2V_UNCONNECTED_416,
  SV2V_UNCONNECTED_417,SV2V_UNCONNECTED_418,SV2V_UNCONNECTED_419,
  SV2V_UNCONNECTED_420,SV2V_UNCONNECTED_421,SV2V_UNCONNECTED_422,
  SV2V_UNCONNECTED_423,SV2V_UNCONNECTED_424,SV2V_UNCONNECTED_425,
  SV2V_UNCONNECTED_426,SV2V_UNCONNECTED_427,SV2V_UNCONNECTED_428,
  SV2V_UNCONNECTED_429,SV2V_UNCONNECTED_430,SV2V_UNCONNECTED_431,SV2V_UNCONNECTED_432,
  SV2V_UNCONNECTED_433,SV2V_UNCONNECTED_434,SV2V_UNCONNECTED_435,
  SV2V_UNCONNECTED_436,SV2V_UNCONNECTED_437,SV2V_UNCONNECTED_438,
  SV2V_UNCONNECTED_439,SV2V_UNCONNECTED_440,SV2V_UNCONNECTED_441,
  SV2V_UNCONNECTED_442,SV2V_UNCONNECTED_443,SV2V_UNCONNECTED_444,
  SV2V_UNCONNECTED_445,SV2V_UNCONNECTED_446,SV2V_UNCONNECTED_447,SV2V_UNCONNECTED_448,
  SV2V_UNCONNECTED_449,SV2V_UNCONNECTED_450,SV2V_UNCONNECTED_451,
  SV2V_UNCONNECTED_452,SV2V_UNCONNECTED_453,SV2V_UNCONNECTED_454,
  SV2V_UNCONNECTED_455,SV2V_UNCONNECTED_456,SV2V_UNCONNECTED_457,
  SV2V_UNCONNECTED_458,SV2V_UNCONNECTED_459,SV2V_UNCONNECTED_460,
  SV2V_UNCONNECTED_461,SV2V_UNCONNECTED_462,SV2V_UNCONNECTED_463,SV2V_UNCONNECTED_464,
  SV2V_UNCONNECTED_465,SV2V_UNCONNECTED_466,SV2V_UNCONNECTED_467,
  SV2V_UNCONNECTED_468,SV2V_UNCONNECTED_469,SV2V_UNCONNECTED_470,
  SV2V_UNCONNECTED_471,SV2V_UNCONNECTED_472,SV2V_UNCONNECTED_473,
  SV2V_UNCONNECTED_474,SV2V_UNCONNECTED_475,SV2V_UNCONNECTED_476,
  SV2V_UNCONNECTED_477,SV2V_UNCONNECTED_478,SV2V_UNCONNECTED_479,SV2V_UNCONNECTED_480,
  SV2V_UNCONNECTED_481,SV2V_UNCONNECTED_482,SV2V_UNCONNECTED_483,
  SV2V_UNCONNECTED_484,SV2V_UNCONNECTED_485,SV2V_UNCONNECTED_486,
  SV2V_UNCONNECTED_487,SV2V_UNCONNECTED_488,SV2V_UNCONNECTED_489,
  SV2V_UNCONNECTED_490,SV2V_UNCONNECTED_491,SV2V_UNCONNECTED_492,
  SV2V_UNCONNECTED_493,SV2V_UNCONNECTED_494,SV2V_UNCONNECTED_495,SV2V_UNCONNECTED_496,
  SV2V_UNCONNECTED_497,SV2V_UNCONNECTED_498,SV2V_UNCONNECTED_499,
  SV2V_UNCONNECTED_500,SV2V_UNCONNECTED_501,SV2V_UNCONNECTED_502,
  SV2V_UNCONNECTED_503,SV2V_UNCONNECTED_504,SV2V_UNCONNECTED_505,
  SV2V_UNCONNECTED_506,SV2V_UNCONNECTED_507,SV2V_UNCONNECTED_508,
  SV2V_UNCONNECTED_509,SV2V_UNCONNECTED_510,SV2V_UNCONNECTED_511,SV2V_UNCONNECTED_512,
  SV2V_UNCONNECTED_513,SV2V_UNCONNECTED_514,SV2V_UNCONNECTED_515,
  SV2V_UNCONNECTED_516,SV2V_UNCONNECTED_517,SV2V_UNCONNECTED_518,
  SV2V_UNCONNECTED_519,SV2V_UNCONNECTED_520,SV2V_UNCONNECTED_521,
  SV2V_UNCONNECTED_522,SV2V_UNCONNECTED_523,SV2V_UNCONNECTED_524,
  SV2V_UNCONNECTED_525,SV2V_UNCONNECTED_526,SV2V_UNCONNECTED_527,SV2V_UNCONNECTED_528,
  SV2V_UNCONNECTED_529,SV2V_UNCONNECTED_530,SV2V_UNCONNECTED_531,
  SV2V_UNCONNECTED_532,SV2V_UNCONNECTED_533,SV2V_UNCONNECTED_534,
  SV2V_UNCONNECTED_535,SV2V_UNCONNECTED_536,SV2V_UNCONNECTED_537,
  SV2V_UNCONNECTED_538,SV2V_UNCONNECTED_539,SV2V_UNCONNECTED_540,
  SV2V_UNCONNECTED_541,SV2V_UNCONNECTED_542,SV2V_UNCONNECTED_543,SV2V_UNCONNECTED_544,
  SV2V_UNCONNECTED_545,SV2V_UNCONNECTED_546,SV2V_UNCONNECTED_547,
  SV2V_UNCONNECTED_548,SV2V_UNCONNECTED_549,SV2V_UNCONNECTED_550,
  SV2V_UNCONNECTED_551,SV2V_UNCONNECTED_552,SV2V_UNCONNECTED_553,
  SV2V_UNCONNECTED_554,SV2V_UNCONNECTED_555,SV2V_UNCONNECTED_556,
  SV2V_UNCONNECTED_557,SV2V_UNCONNECTED_558,SV2V_UNCONNECTED_559,SV2V_UNCONNECTED_560,
  SV2V_UNCONNECTED_561,SV2V_UNCONNECTED_562,SV2V_UNCONNECTED_563,
  SV2V_UNCONNECTED_564,SV2V_UNCONNECTED_565,SV2V_UNCONNECTED_566,
  SV2V_UNCONNECTED_567,SV2V_UNCONNECTED_568,SV2V_UNCONNECTED_569,
  SV2V_UNCONNECTED_570,SV2V_UNCONNECTED_571,SV2V_UNCONNECTED_572,
  SV2V_UNCONNECTED_573,SV2V_UNCONNECTED_574,SV2V_UNCONNECTED_575,SV2V_UNCONNECTED_576,
  SV2V_UNCONNECTED_577,SV2V_UNCONNECTED_578,SV2V_UNCONNECTED_579,
  SV2V_UNCONNECTED_580,SV2V_UNCONNECTED_581,SV2V_UNCONNECTED_582,
  SV2V_UNCONNECTED_583,SV2V_UNCONNECTED_584,SV2V_UNCONNECTED_585,
  SV2V_UNCONNECTED_586,SV2V_UNCONNECTED_587,SV2V_UNCONNECTED_588,
  SV2V_UNCONNECTED_589,SV2V_UNCONNECTED_590,SV2V_UNCONNECTED_591,SV2V_UNCONNECTED_592,
  SV2V_UNCONNECTED_593,SV2V_UNCONNECTED_594,SV2V_UNCONNECTED_595,
  SV2V_UNCONNECTED_596,SV2V_UNCONNECTED_597,SV2V_UNCONNECTED_598,
  SV2V_UNCONNECTED_599,SV2V_UNCONNECTED_600,SV2V_UNCONNECTED_601,
  SV2V_UNCONNECTED_602,SV2V_UNCONNECTED_603,SV2V_UNCONNECTED_604,
  SV2V_UNCONNECTED_605,SV2V_UNCONNECTED_606,SV2V_UNCONNECTED_607,SV2V_UNCONNECTED_608,
  SV2V_UNCONNECTED_609,SV2V_UNCONNECTED_610,SV2V_UNCONNECTED_611,
  SV2V_UNCONNECTED_612,SV2V_UNCONNECTED_613,SV2V_UNCONNECTED_614,
  SV2V_UNCONNECTED_615,SV2V_UNCONNECTED_616,SV2V_UNCONNECTED_617,
  SV2V_UNCONNECTED_618,SV2V_UNCONNECTED_619,SV2V_UNCONNECTED_620,
  SV2V_UNCONNECTED_621,SV2V_UNCONNECTED_622,SV2V_UNCONNECTED_623,SV2V_UNCONNECTED_624,
  SV2V_UNCONNECTED_625,SV2V_UNCONNECTED_626,SV2V_UNCONNECTED_627,
  SV2V_UNCONNECTED_628,SV2V_UNCONNECTED_629,SV2V_UNCONNECTED_630,
  SV2V_UNCONNECTED_631,SV2V_UNCONNECTED_632,SV2V_UNCONNECTED_633,
  SV2V_UNCONNECTED_634,SV2V_UNCONNECTED_635,SV2V_UNCONNECTED_636,
  SV2V_UNCONNECTED_637,SV2V_UNCONNECTED_638,SV2V_UNCONNECTED_639,SV2V_UNCONNECTED_640,
  SV2V_UNCONNECTED_641,SV2V_UNCONNECTED_642,SV2V_UNCONNECTED_643,
  SV2V_UNCONNECTED_644,SV2V_UNCONNECTED_645,SV2V_UNCONNECTED_646,
  SV2V_UNCONNECTED_647,SV2V_UNCONNECTED_648,SV2V_UNCONNECTED_649,
  SV2V_UNCONNECTED_650,SV2V_UNCONNECTED_651,SV2V_UNCONNECTED_652,
  SV2V_UNCONNECTED_653,SV2V_UNCONNECTED_654,SV2V_UNCONNECTED_655,SV2V_UNCONNECTED_656,
  SV2V_UNCONNECTED_657,SV2V_UNCONNECTED_658,SV2V_UNCONNECTED_659,
  SV2V_UNCONNECTED_660,SV2V_UNCONNECTED_661,SV2V_UNCONNECTED_662,
  SV2V_UNCONNECTED_663,SV2V_UNCONNECTED_664,SV2V_UNCONNECTED_665,
  SV2V_UNCONNECTED_666,SV2V_UNCONNECTED_667,SV2V_UNCONNECTED_668,
  SV2V_UNCONNECTED_669,SV2V_UNCONNECTED_670,SV2V_UNCONNECTED_671,SV2V_UNCONNECTED_672,
  SV2V_UNCONNECTED_673,SV2V_UNCONNECTED_674,SV2V_UNCONNECTED_675,
  SV2V_UNCONNECTED_676,SV2V_UNCONNECTED_677,SV2V_UNCONNECTED_678,
  SV2V_UNCONNECTED_679,SV2V_UNCONNECTED_680,SV2V_UNCONNECTED_681,
  SV2V_UNCONNECTED_682,SV2V_UNCONNECTED_683,SV2V_UNCONNECTED_684,
  SV2V_UNCONNECTED_685,SV2V_UNCONNECTED_686,SV2V_UNCONNECTED_687,SV2V_UNCONNECTED_688,
  SV2V_UNCONNECTED_689,SV2V_UNCONNECTED_690,SV2V_UNCONNECTED_691,
  SV2V_UNCONNECTED_692,SV2V_UNCONNECTED_693,SV2V_UNCONNECTED_694,
  SV2V_UNCONNECTED_695,SV2V_UNCONNECTED_696,SV2V_UNCONNECTED_697,
  SV2V_UNCONNECTED_698,SV2V_UNCONNECTED_699,SV2V_UNCONNECTED_700,
  SV2V_UNCONNECTED_701,SV2V_UNCONNECTED_702,SV2V_UNCONNECTED_703,SV2V_UNCONNECTED_704,
  SV2V_UNCONNECTED_705,SV2V_UNCONNECTED_706,SV2V_UNCONNECTED_707,
  SV2V_UNCONNECTED_708,SV2V_UNCONNECTED_709,SV2V_UNCONNECTED_710,
  SV2V_UNCONNECTED_711,SV2V_UNCONNECTED_712,SV2V_UNCONNECTED_713,
  SV2V_UNCONNECTED_714,SV2V_UNCONNECTED_715,SV2V_UNCONNECTED_716,
  SV2V_UNCONNECTED_717,SV2V_UNCONNECTED_718,SV2V_UNCONNECTED_719,SV2V_UNCONNECTED_720,
  SV2V_UNCONNECTED_721,SV2V_UNCONNECTED_722,SV2V_UNCONNECTED_723,
  SV2V_UNCONNECTED_724,SV2V_UNCONNECTED_725,SV2V_UNCONNECTED_726,
  SV2V_UNCONNECTED_727,SV2V_UNCONNECTED_728,SV2V_UNCONNECTED_729,
  SV2V_UNCONNECTED_730,SV2V_UNCONNECTED_731,SV2V_UNCONNECTED_732,
  SV2V_UNCONNECTED_733,SV2V_UNCONNECTED_734,SV2V_UNCONNECTED_735,SV2V_UNCONNECTED_736,
  SV2V_UNCONNECTED_737,SV2V_UNCONNECTED_738,SV2V_UNCONNECTED_739,
  SV2V_UNCONNECTED_740,SV2V_UNCONNECTED_741,SV2V_UNCONNECTED_742,
  SV2V_UNCONNECTED_743,SV2V_UNCONNECTED_744,SV2V_UNCONNECTED_745,
  SV2V_UNCONNECTED_746,SV2V_UNCONNECTED_747,SV2V_UNCONNECTED_748,
  SV2V_UNCONNECTED_749,SV2V_UNCONNECTED_750,SV2V_UNCONNECTED_751,SV2V_UNCONNECTED_752,
  SV2V_UNCONNECTED_753,SV2V_UNCONNECTED_754,SV2V_UNCONNECTED_755,
  SV2V_UNCONNECTED_756,SV2V_UNCONNECTED_757,SV2V_UNCONNECTED_758,
  SV2V_UNCONNECTED_759,SV2V_UNCONNECTED_760,SV2V_UNCONNECTED_761,
  SV2V_UNCONNECTED_762,SV2V_UNCONNECTED_763,SV2V_UNCONNECTED_764,
  SV2V_UNCONNECTED_765,SV2V_UNCONNECTED_766,SV2V_UNCONNECTED_767,SV2V_UNCONNECTED_768,
  SV2V_UNCONNECTED_769,SV2V_UNCONNECTED_770,SV2V_UNCONNECTED_771,
  SV2V_UNCONNECTED_772,SV2V_UNCONNECTED_773,SV2V_UNCONNECTED_774,
  SV2V_UNCONNECTED_775,SV2V_UNCONNECTED_776,SV2V_UNCONNECTED_777,
  SV2V_UNCONNECTED_778,SV2V_UNCONNECTED_779,SV2V_UNCONNECTED_780,
  SV2V_UNCONNECTED_781,SV2V_UNCONNECTED_782,SV2V_UNCONNECTED_783,SV2V_UNCONNECTED_784,
  SV2V_UNCONNECTED_785,SV2V_UNCONNECTED_786,SV2V_UNCONNECTED_787,
  SV2V_UNCONNECTED_788,SV2V_UNCONNECTED_789,SV2V_UNCONNECTED_790,
  SV2V_UNCONNECTED_791,SV2V_UNCONNECTED_792,SV2V_UNCONNECTED_793,
  SV2V_UNCONNECTED_794,SV2V_UNCONNECTED_795,SV2V_UNCONNECTED_796,
  SV2V_UNCONNECTED_797,SV2V_UNCONNECTED_798,SV2V_UNCONNECTED_799,SV2V_UNCONNECTED_800,
  SV2V_UNCONNECTED_801,SV2V_UNCONNECTED_802,SV2V_UNCONNECTED_803,
  SV2V_UNCONNECTED_804,SV2V_UNCONNECTED_805,SV2V_UNCONNECTED_806,
  SV2V_UNCONNECTED_807,SV2V_UNCONNECTED_808,SV2V_UNCONNECTED_809,
  SV2V_UNCONNECTED_810,SV2V_UNCONNECTED_811,SV2V_UNCONNECTED_812,
  SV2V_UNCONNECTED_813,SV2V_UNCONNECTED_814,SV2V_UNCONNECTED_815,SV2V_UNCONNECTED_816,
  SV2V_UNCONNECTED_817,SV2V_UNCONNECTED_818,SV2V_UNCONNECTED_819,
  SV2V_UNCONNECTED_820,SV2V_UNCONNECTED_821,SV2V_UNCONNECTED_822,
  SV2V_UNCONNECTED_823,SV2V_UNCONNECTED_824,SV2V_UNCONNECTED_825,
  SV2V_UNCONNECTED_826,SV2V_UNCONNECTED_827,SV2V_UNCONNECTED_828,
  SV2V_UNCONNECTED_829,SV2V_UNCONNECTED_830,SV2V_UNCONNECTED_831,SV2V_UNCONNECTED_832,
  SV2V_UNCONNECTED_833,SV2V_UNCONNECTED_834,SV2V_UNCONNECTED_835,
  SV2V_UNCONNECTED_836,SV2V_UNCONNECTED_837,SV2V_UNCONNECTED_838,
  SV2V_UNCONNECTED_839,SV2V_UNCONNECTED_840,SV2V_UNCONNECTED_841,
  SV2V_UNCONNECTED_842,SV2V_UNCONNECTED_843,SV2V_UNCONNECTED_844,
  SV2V_UNCONNECTED_845,SV2V_UNCONNECTED_846,SV2V_UNCONNECTED_847,SV2V_UNCONNECTED_848,
  SV2V_UNCONNECTED_849,SV2V_UNCONNECTED_850,SV2V_UNCONNECTED_851,
  SV2V_UNCONNECTED_852,SV2V_UNCONNECTED_853,SV2V_UNCONNECTED_854,
  SV2V_UNCONNECTED_855,SV2V_UNCONNECTED_856,SV2V_UNCONNECTED_857,
  SV2V_UNCONNECTED_858,SV2V_UNCONNECTED_859,SV2V_UNCONNECTED_860,
  SV2V_UNCONNECTED_861,SV2V_UNCONNECTED_862,SV2V_UNCONNECTED_863,SV2V_UNCONNECTED_864,
  SV2V_UNCONNECTED_865,SV2V_UNCONNECTED_866,SV2V_UNCONNECTED_867,
  SV2V_UNCONNECTED_868,SV2V_UNCONNECTED_869,SV2V_UNCONNECTED_870,
  SV2V_UNCONNECTED_871,SV2V_UNCONNECTED_872,SV2V_UNCONNECTED_873,
  SV2V_UNCONNECTED_874,SV2V_UNCONNECTED_875,SV2V_UNCONNECTED_876,
  SV2V_UNCONNECTED_877,SV2V_UNCONNECTED_878,SV2V_UNCONNECTED_879,SV2V_UNCONNECTED_880,
  SV2V_UNCONNECTED_881,SV2V_UNCONNECTED_882,SV2V_UNCONNECTED_883,
  SV2V_UNCONNECTED_884,SV2V_UNCONNECTED_885,SV2V_UNCONNECTED_886,
  SV2V_UNCONNECTED_887,SV2V_UNCONNECTED_888,SV2V_UNCONNECTED_889,
  SV2V_UNCONNECTED_890,SV2V_UNCONNECTED_891,SV2V_UNCONNECTED_892,
  SV2V_UNCONNECTED_893,SV2V_UNCONNECTED_894,SV2V_UNCONNECTED_895,SV2V_UNCONNECTED_896,
  SV2V_UNCONNECTED_897,SV2V_UNCONNECTED_898,SV2V_UNCONNECTED_899,
  SV2V_UNCONNECTED_900,SV2V_UNCONNECTED_901,SV2V_UNCONNECTED_902,
  SV2V_UNCONNECTED_903,SV2V_UNCONNECTED_904,SV2V_UNCONNECTED_905,
  SV2V_UNCONNECTED_906,SV2V_UNCONNECTED_907,SV2V_UNCONNECTED_908,
  SV2V_UNCONNECTED_909,SV2V_UNCONNECTED_910,SV2V_UNCONNECTED_911,SV2V_UNCONNECTED_912,
  SV2V_UNCONNECTED_913,SV2V_UNCONNECTED_914,SV2V_UNCONNECTED_915,
  SV2V_UNCONNECTED_916,SV2V_UNCONNECTED_917,SV2V_UNCONNECTED_918,
  SV2V_UNCONNECTED_919,SV2V_UNCONNECTED_920,SV2V_UNCONNECTED_921,
  SV2V_UNCONNECTED_922,SV2V_UNCONNECTED_923,SV2V_UNCONNECTED_924,
  SV2V_UNCONNECTED_925,SV2V_UNCONNECTED_926,SV2V_UNCONNECTED_927,SV2V_UNCONNECTED_928,
  SV2V_UNCONNECTED_929,SV2V_UNCONNECTED_930,SV2V_UNCONNECTED_931,
  SV2V_UNCONNECTED_932,SV2V_UNCONNECTED_933,SV2V_UNCONNECTED_934,
  SV2V_UNCONNECTED_935,SV2V_UNCONNECTED_936,SV2V_UNCONNECTED_937,
  SV2V_UNCONNECTED_938,SV2V_UNCONNECTED_939,SV2V_UNCONNECTED_940,
  SV2V_UNCONNECTED_941,SV2V_UNCONNECTED_942,SV2V_UNCONNECTED_943,SV2V_UNCONNECTED_944,
  SV2V_UNCONNECTED_945,SV2V_UNCONNECTED_946,SV2V_UNCONNECTED_947,
  SV2V_UNCONNECTED_948,SV2V_UNCONNECTED_949,SV2V_UNCONNECTED_950,
  SV2V_UNCONNECTED_951,SV2V_UNCONNECTED_952,SV2V_UNCONNECTED_953,
  SV2V_UNCONNECTED_954,SV2V_UNCONNECTED_955,SV2V_UNCONNECTED_956,
  SV2V_UNCONNECTED_957,SV2V_UNCONNECTED_958,SV2V_UNCONNECTED_959,SV2V_UNCONNECTED_960,
  SV2V_UNCONNECTED_961,SV2V_UNCONNECTED_962,SV2V_UNCONNECTED_963,
  SV2V_UNCONNECTED_964,SV2V_UNCONNECTED_965,SV2V_UNCONNECTED_966,
  SV2V_UNCONNECTED_967,SV2V_UNCONNECTED_968,SV2V_UNCONNECTED_969,
  SV2V_UNCONNECTED_970,SV2V_UNCONNECTED_971,SV2V_UNCONNECTED_972,
  SV2V_UNCONNECTED_973,SV2V_UNCONNECTED_974,SV2V_UNCONNECTED_975,SV2V_UNCONNECTED_976,
  SV2V_UNCONNECTED_977,SV2V_UNCONNECTED_978,SV2V_UNCONNECTED_979,
  SV2V_UNCONNECTED_980,SV2V_UNCONNECTED_981,SV2V_UNCONNECTED_982,
  SV2V_UNCONNECTED_983,SV2V_UNCONNECTED_984,SV2V_UNCONNECTED_985,
  SV2V_UNCONNECTED_986,SV2V_UNCONNECTED_987,SV2V_UNCONNECTED_988,
  SV2V_UNCONNECTED_989,SV2V_UNCONNECTED_990,SV2V_UNCONNECTED_991,SV2V_UNCONNECTED_992,
  SV2V_UNCONNECTED_993,SV2V_UNCONNECTED_994,SV2V_UNCONNECTED_995,
  SV2V_UNCONNECTED_996,SV2V_UNCONNECTED_997,SV2V_UNCONNECTED_998,
  SV2V_UNCONNECTED_999,SV2V_UNCONNECTED_1000,SV2V_UNCONNECTED_1001,
  SV2V_UNCONNECTED_1002,SV2V_UNCONNECTED_1003,SV2V_UNCONNECTED_1004,
  SV2V_UNCONNECTED_1005,SV2V_UNCONNECTED_1006,SV2V_UNCONNECTED_1007,
  SV2V_UNCONNECTED_1008,SV2V_UNCONNECTED_1009,SV2V_UNCONNECTED_1010,
  SV2V_UNCONNECTED_1011,SV2V_UNCONNECTED_1012,SV2V_UNCONNECTED_1013,
  SV2V_UNCONNECTED_1014,SV2V_UNCONNECTED_1015,SV2V_UNCONNECTED_1016,SV2V_UNCONNECTED_1017,
  SV2V_UNCONNECTED_1018,SV2V_UNCONNECTED_1019,SV2V_UNCONNECTED_1020,
  SV2V_UNCONNECTED_1021,SV2V_UNCONNECTED_1022,SV2V_UNCONNECTED_1023,
  SV2V_UNCONNECTED_1024,SV2V_UNCONNECTED_1025,SV2V_UNCONNECTED_1026,
  SV2V_UNCONNECTED_1027,SV2V_UNCONNECTED_1028,SV2V_UNCONNECTED_1029,
  SV2V_UNCONNECTED_1030,SV2V_UNCONNECTED_1031,SV2V_UNCONNECTED_1032,
  SV2V_UNCONNECTED_1033,SV2V_UNCONNECTED_1034,SV2V_UNCONNECTED_1035,
  SV2V_UNCONNECTED_1036,SV2V_UNCONNECTED_1037,SV2V_UNCONNECTED_1038,
  SV2V_UNCONNECTED_1039,SV2V_UNCONNECTED_1040,SV2V_UNCONNECTED_1041,
  SV2V_UNCONNECTED_1042,SV2V_UNCONNECTED_1043,SV2V_UNCONNECTED_1044,
  SV2V_UNCONNECTED_1045,SV2V_UNCONNECTED_1046,SV2V_UNCONNECTED_1047,
  SV2V_UNCONNECTED_1048,SV2V_UNCONNECTED_1049,SV2V_UNCONNECTED_1050,
  SV2V_UNCONNECTED_1051,SV2V_UNCONNECTED_1052,SV2V_UNCONNECTED_1053,
  SV2V_UNCONNECTED_1054,SV2V_UNCONNECTED_1055,SV2V_UNCONNECTED_1056,SV2V_UNCONNECTED_1057,
  SV2V_UNCONNECTED_1058,SV2V_UNCONNECTED_1059,SV2V_UNCONNECTED_1060,
  SV2V_UNCONNECTED_1061,SV2V_UNCONNECTED_1062,SV2V_UNCONNECTED_1063,
  SV2V_UNCONNECTED_1064,SV2V_UNCONNECTED_1065,SV2V_UNCONNECTED_1066,
  SV2V_UNCONNECTED_1067,SV2V_UNCONNECTED_1068,SV2V_UNCONNECTED_1069,
  SV2V_UNCONNECTED_1070,SV2V_UNCONNECTED_1071,SV2V_UNCONNECTED_1072,
  SV2V_UNCONNECTED_1073,SV2V_UNCONNECTED_1074,SV2V_UNCONNECTED_1075,
  SV2V_UNCONNECTED_1076,SV2V_UNCONNECTED_1077,SV2V_UNCONNECTED_1078,
  SV2V_UNCONNECTED_1079,SV2V_UNCONNECTED_1080,SV2V_UNCONNECTED_1081,
  SV2V_UNCONNECTED_1082,SV2V_UNCONNECTED_1083,SV2V_UNCONNECTED_1084,
  SV2V_UNCONNECTED_1085,SV2V_UNCONNECTED_1086,SV2V_UNCONNECTED_1087,
  SV2V_UNCONNECTED_1088,SV2V_UNCONNECTED_1089,SV2V_UNCONNECTED_1090,
  SV2V_UNCONNECTED_1091,SV2V_UNCONNECTED_1092,SV2V_UNCONNECTED_1093,
  SV2V_UNCONNECTED_1094,SV2V_UNCONNECTED_1095,SV2V_UNCONNECTED_1096,SV2V_UNCONNECTED_1097,
  SV2V_UNCONNECTED_1098,SV2V_UNCONNECTED_1099,SV2V_UNCONNECTED_1100,
  SV2V_UNCONNECTED_1101,SV2V_UNCONNECTED_1102,SV2V_UNCONNECTED_1103,
  SV2V_UNCONNECTED_1104,SV2V_UNCONNECTED_1105,SV2V_UNCONNECTED_1106,
  SV2V_UNCONNECTED_1107,SV2V_UNCONNECTED_1108,SV2V_UNCONNECTED_1109,
  SV2V_UNCONNECTED_1110,SV2V_UNCONNECTED_1111,SV2V_UNCONNECTED_1112,
  SV2V_UNCONNECTED_1113,SV2V_UNCONNECTED_1114,SV2V_UNCONNECTED_1115,
  SV2V_UNCONNECTED_1116,SV2V_UNCONNECTED_1117,SV2V_UNCONNECTED_1118,
  SV2V_UNCONNECTED_1119,SV2V_UNCONNECTED_1120,SV2V_UNCONNECTED_1121,
  SV2V_UNCONNECTED_1122,SV2V_UNCONNECTED_1123,SV2V_UNCONNECTED_1124,
  SV2V_UNCONNECTED_1125,SV2V_UNCONNECTED_1126,SV2V_UNCONNECTED_1127,
  SV2V_UNCONNECTED_1128,SV2V_UNCONNECTED_1129,SV2V_UNCONNECTED_1130,
  SV2V_UNCONNECTED_1131,SV2V_UNCONNECTED_1132,SV2V_UNCONNECTED_1133,
  SV2V_UNCONNECTED_1134,SV2V_UNCONNECTED_1135,SV2V_UNCONNECTED_1136,SV2V_UNCONNECTED_1137,
  SV2V_UNCONNECTED_1138,SV2V_UNCONNECTED_1139,SV2V_UNCONNECTED_1140,
  SV2V_UNCONNECTED_1141,SV2V_UNCONNECTED_1142,SV2V_UNCONNECTED_1143,
  SV2V_UNCONNECTED_1144,SV2V_UNCONNECTED_1145,SV2V_UNCONNECTED_1146,
  SV2V_UNCONNECTED_1147,SV2V_UNCONNECTED_1148,SV2V_UNCONNECTED_1149,
  SV2V_UNCONNECTED_1150,SV2V_UNCONNECTED_1151,SV2V_UNCONNECTED_1152,
  SV2V_UNCONNECTED_1153,SV2V_UNCONNECTED_1154,SV2V_UNCONNECTED_1155,
  SV2V_UNCONNECTED_1156,SV2V_UNCONNECTED_1157,SV2V_UNCONNECTED_1158,
  SV2V_UNCONNECTED_1159,SV2V_UNCONNECTED_1160,SV2V_UNCONNECTED_1161,
  SV2V_UNCONNECTED_1162,SV2V_UNCONNECTED_1163,SV2V_UNCONNECTED_1164,
  SV2V_UNCONNECTED_1165,SV2V_UNCONNECTED_1166,SV2V_UNCONNECTED_1167,
  SV2V_UNCONNECTED_1168,SV2V_UNCONNECTED_1169,SV2V_UNCONNECTED_1170,
  SV2V_UNCONNECTED_1171,SV2V_UNCONNECTED_1172,SV2V_UNCONNECTED_1173,
  SV2V_UNCONNECTED_1174,SV2V_UNCONNECTED_1175,SV2V_UNCONNECTED_1176,SV2V_UNCONNECTED_1177,
  SV2V_UNCONNECTED_1178,SV2V_UNCONNECTED_1179,SV2V_UNCONNECTED_1180,
  SV2V_UNCONNECTED_1181,SV2V_UNCONNECTED_1182,SV2V_UNCONNECTED_1183,
  SV2V_UNCONNECTED_1184,SV2V_UNCONNECTED_1185,SV2V_UNCONNECTED_1186,
  SV2V_UNCONNECTED_1187,SV2V_UNCONNECTED_1188,SV2V_UNCONNECTED_1189,
  SV2V_UNCONNECTED_1190,SV2V_UNCONNECTED_1191,SV2V_UNCONNECTED_1192,
  SV2V_UNCONNECTED_1193,SV2V_UNCONNECTED_1194,SV2V_UNCONNECTED_1195,
  SV2V_UNCONNECTED_1196,SV2V_UNCONNECTED_1197,SV2V_UNCONNECTED_1198,
  SV2V_UNCONNECTED_1199,SV2V_UNCONNECTED_1200,SV2V_UNCONNECTED_1201,
  SV2V_UNCONNECTED_1202,SV2V_UNCONNECTED_1203,SV2V_UNCONNECTED_1204,
  SV2V_UNCONNECTED_1205,SV2V_UNCONNECTED_1206,SV2V_UNCONNECTED_1207,
  SV2V_UNCONNECTED_1208,SV2V_UNCONNECTED_1209,SV2V_UNCONNECTED_1210,
  SV2V_UNCONNECTED_1211,SV2V_UNCONNECTED_1212,SV2V_UNCONNECTED_1213,
  SV2V_UNCONNECTED_1214,SV2V_UNCONNECTED_1215,SV2V_UNCONNECTED_1216,SV2V_UNCONNECTED_1217,
  SV2V_UNCONNECTED_1218,SV2V_UNCONNECTED_1219,SV2V_UNCONNECTED_1220,
  SV2V_UNCONNECTED_1221,SV2V_UNCONNECTED_1222,SV2V_UNCONNECTED_1223,
  SV2V_UNCONNECTED_1224,SV2V_UNCONNECTED_1225,SV2V_UNCONNECTED_1226,
  SV2V_UNCONNECTED_1227,SV2V_UNCONNECTED_1228,SV2V_UNCONNECTED_1229,
  SV2V_UNCONNECTED_1230,SV2V_UNCONNECTED_1231,SV2V_UNCONNECTED_1232,
  SV2V_UNCONNECTED_1233,SV2V_UNCONNECTED_1234,SV2V_UNCONNECTED_1235,
  SV2V_UNCONNECTED_1236,SV2V_UNCONNECTED_1237,SV2V_UNCONNECTED_1238,
  SV2V_UNCONNECTED_1239,SV2V_UNCONNECTED_1240,SV2V_UNCONNECTED_1241,
  SV2V_UNCONNECTED_1242,SV2V_UNCONNECTED_1243,SV2V_UNCONNECTED_1244,
  SV2V_UNCONNECTED_1245,SV2V_UNCONNECTED_1246,SV2V_UNCONNECTED_1247,
  SV2V_UNCONNECTED_1248,SV2V_UNCONNECTED_1249,SV2V_UNCONNECTED_1250,
  SV2V_UNCONNECTED_1251,SV2V_UNCONNECTED_1252,SV2V_UNCONNECTED_1253,
  SV2V_UNCONNECTED_1254,SV2V_UNCONNECTED_1255,SV2V_UNCONNECTED_1256,SV2V_UNCONNECTED_1257,
  SV2V_UNCONNECTED_1258,SV2V_UNCONNECTED_1259,SV2V_UNCONNECTED_1260,
  SV2V_UNCONNECTED_1261,SV2V_UNCONNECTED_1262,SV2V_UNCONNECTED_1263,
  SV2V_UNCONNECTED_1264,SV2V_UNCONNECTED_1265,SV2V_UNCONNECTED_1266,
  SV2V_UNCONNECTED_1267,SV2V_UNCONNECTED_1268,SV2V_UNCONNECTED_1269,
  SV2V_UNCONNECTED_1270,SV2V_UNCONNECTED_1271,SV2V_UNCONNECTED_1272,
  SV2V_UNCONNECTED_1273,SV2V_UNCONNECTED_1274,SV2V_UNCONNECTED_1275,
  SV2V_UNCONNECTED_1276,SV2V_UNCONNECTED_1277,SV2V_UNCONNECTED_1278,
  SV2V_UNCONNECTED_1279,SV2V_UNCONNECTED_1280,SV2V_UNCONNECTED_1281,
  SV2V_UNCONNECTED_1282,SV2V_UNCONNECTED_1283,SV2V_UNCONNECTED_1284,
  SV2V_UNCONNECTED_1285,SV2V_UNCONNECTED_1286,SV2V_UNCONNECTED_1287,
  SV2V_UNCONNECTED_1288,SV2V_UNCONNECTED_1289,SV2V_UNCONNECTED_1290,
  SV2V_UNCONNECTED_1291,SV2V_UNCONNECTED_1292,SV2V_UNCONNECTED_1293,
  SV2V_UNCONNECTED_1294,SV2V_UNCONNECTED_1295,SV2V_UNCONNECTED_1296,SV2V_UNCONNECTED_1297,
  SV2V_UNCONNECTED_1298,SV2V_UNCONNECTED_1299,SV2V_UNCONNECTED_1300,
  SV2V_UNCONNECTED_1301,SV2V_UNCONNECTED_1302,SV2V_UNCONNECTED_1303,
  SV2V_UNCONNECTED_1304,SV2V_UNCONNECTED_1305,SV2V_UNCONNECTED_1306,
  SV2V_UNCONNECTED_1307,SV2V_UNCONNECTED_1308,SV2V_UNCONNECTED_1309,
  SV2V_UNCONNECTED_1310,SV2V_UNCONNECTED_1311,SV2V_UNCONNECTED_1312,
  SV2V_UNCONNECTED_1313,SV2V_UNCONNECTED_1314,SV2V_UNCONNECTED_1315,
  SV2V_UNCONNECTED_1316,SV2V_UNCONNECTED_1317,SV2V_UNCONNECTED_1318,
  SV2V_UNCONNECTED_1319,SV2V_UNCONNECTED_1320,SV2V_UNCONNECTED_1321,
  SV2V_UNCONNECTED_1322,SV2V_UNCONNECTED_1323,SV2V_UNCONNECTED_1324,
  SV2V_UNCONNECTED_1325,SV2V_UNCONNECTED_1326,SV2V_UNCONNECTED_1327,
  SV2V_UNCONNECTED_1328,SV2V_UNCONNECTED_1329,SV2V_UNCONNECTED_1330,
  SV2V_UNCONNECTED_1331,SV2V_UNCONNECTED_1332,SV2V_UNCONNECTED_1333,
  SV2V_UNCONNECTED_1334,SV2V_UNCONNECTED_1335,SV2V_UNCONNECTED_1336,SV2V_UNCONNECTED_1337,
  SV2V_UNCONNECTED_1338,SV2V_UNCONNECTED_1339,SV2V_UNCONNECTED_1340,
  SV2V_UNCONNECTED_1341,SV2V_UNCONNECTED_1342,SV2V_UNCONNECTED_1343,
  SV2V_UNCONNECTED_1344,SV2V_UNCONNECTED_1345,SV2V_UNCONNECTED_1346,
  SV2V_UNCONNECTED_1347,SV2V_UNCONNECTED_1348,SV2V_UNCONNECTED_1349,
  SV2V_UNCONNECTED_1350,SV2V_UNCONNECTED_1351,SV2V_UNCONNECTED_1352,
  SV2V_UNCONNECTED_1353,SV2V_UNCONNECTED_1354,SV2V_UNCONNECTED_1355,
  SV2V_UNCONNECTED_1356,SV2V_UNCONNECTED_1357,SV2V_UNCONNECTED_1358,
  SV2V_UNCONNECTED_1359,SV2V_UNCONNECTED_1360,SV2V_UNCONNECTED_1361,
  SV2V_UNCONNECTED_1362,SV2V_UNCONNECTED_1363,SV2V_UNCONNECTED_1364,
  SV2V_UNCONNECTED_1365,SV2V_UNCONNECTED_1366,SV2V_UNCONNECTED_1367,
  SV2V_UNCONNECTED_1368,SV2V_UNCONNECTED_1369,SV2V_UNCONNECTED_1370,
  SV2V_UNCONNECTED_1371,SV2V_UNCONNECTED_1372,SV2V_UNCONNECTED_1373,
  SV2V_UNCONNECTED_1374,SV2V_UNCONNECTED_1375,SV2V_UNCONNECTED_1376,SV2V_UNCONNECTED_1377,
  SV2V_UNCONNECTED_1378,SV2V_UNCONNECTED_1379,SV2V_UNCONNECTED_1380,
  SV2V_UNCONNECTED_1381,SV2V_UNCONNECTED_1382,SV2V_UNCONNECTED_1383,
  SV2V_UNCONNECTED_1384,SV2V_UNCONNECTED_1385,SV2V_UNCONNECTED_1386,
  SV2V_UNCONNECTED_1387,SV2V_UNCONNECTED_1388,SV2V_UNCONNECTED_1389,
  SV2V_UNCONNECTED_1390,SV2V_UNCONNECTED_1391,SV2V_UNCONNECTED_1392,
  SV2V_UNCONNECTED_1393,SV2V_UNCONNECTED_1394,SV2V_UNCONNECTED_1395,
  SV2V_UNCONNECTED_1396,SV2V_UNCONNECTED_1397,SV2V_UNCONNECTED_1398,
  SV2V_UNCONNECTED_1399,SV2V_UNCONNECTED_1400,SV2V_UNCONNECTED_1401,
  SV2V_UNCONNECTED_1402,SV2V_UNCONNECTED_1403,SV2V_UNCONNECTED_1404,
  SV2V_UNCONNECTED_1405,SV2V_UNCONNECTED_1406,SV2V_UNCONNECTED_1407,
  SV2V_UNCONNECTED_1408,SV2V_UNCONNECTED_1409,SV2V_UNCONNECTED_1410,
  SV2V_UNCONNECTED_1411,SV2V_UNCONNECTED_1412,SV2V_UNCONNECTED_1413,
  SV2V_UNCONNECTED_1414,SV2V_UNCONNECTED_1415,SV2V_UNCONNECTED_1416,SV2V_UNCONNECTED_1417,
  SV2V_UNCONNECTED_1418,SV2V_UNCONNECTED_1419,SV2V_UNCONNECTED_1420,
  SV2V_UNCONNECTED_1421,SV2V_UNCONNECTED_1422,SV2V_UNCONNECTED_1423,
  SV2V_UNCONNECTED_1424,SV2V_UNCONNECTED_1425,SV2V_UNCONNECTED_1426,
  SV2V_UNCONNECTED_1427,SV2V_UNCONNECTED_1428,SV2V_UNCONNECTED_1429,
  SV2V_UNCONNECTED_1430,SV2V_UNCONNECTED_1431,SV2V_UNCONNECTED_1432,
  SV2V_UNCONNECTED_1433,SV2V_UNCONNECTED_1434,SV2V_UNCONNECTED_1435,
  SV2V_UNCONNECTED_1436,SV2V_UNCONNECTED_1437,SV2V_UNCONNECTED_1438,
  SV2V_UNCONNECTED_1439,SV2V_UNCONNECTED_1440,SV2V_UNCONNECTED_1441,
  SV2V_UNCONNECTED_1442,SV2V_UNCONNECTED_1443,SV2V_UNCONNECTED_1444,
  SV2V_UNCONNECTED_1445,SV2V_UNCONNECTED_1446,SV2V_UNCONNECTED_1447,
  SV2V_UNCONNECTED_1448,SV2V_UNCONNECTED_1449,SV2V_UNCONNECTED_1450,
  SV2V_UNCONNECTED_1451,SV2V_UNCONNECTED_1452,SV2V_UNCONNECTED_1453,
  SV2V_UNCONNECTED_1454,SV2V_UNCONNECTED_1455,SV2V_UNCONNECTED_1456,SV2V_UNCONNECTED_1457,
  SV2V_UNCONNECTED_1458,SV2V_UNCONNECTED_1459,SV2V_UNCONNECTED_1460,
  SV2V_UNCONNECTED_1461,SV2V_UNCONNECTED_1462,SV2V_UNCONNECTED_1463,
  SV2V_UNCONNECTED_1464,SV2V_UNCONNECTED_1465,SV2V_UNCONNECTED_1466,
  SV2V_UNCONNECTED_1467,SV2V_UNCONNECTED_1468,SV2V_UNCONNECTED_1469,
  SV2V_UNCONNECTED_1470,SV2V_UNCONNECTED_1471,SV2V_UNCONNECTED_1472,
  SV2V_UNCONNECTED_1473,SV2V_UNCONNECTED_1474,SV2V_UNCONNECTED_1475,
  SV2V_UNCONNECTED_1476,SV2V_UNCONNECTED_1477,SV2V_UNCONNECTED_1478,
  SV2V_UNCONNECTED_1479,SV2V_UNCONNECTED_1480,SV2V_UNCONNECTED_1481,
  SV2V_UNCONNECTED_1482,SV2V_UNCONNECTED_1483,SV2V_UNCONNECTED_1484,
  SV2V_UNCONNECTED_1485,SV2V_UNCONNECTED_1486,SV2V_UNCONNECTED_1487,
  SV2V_UNCONNECTED_1488,SV2V_UNCONNECTED_1489,SV2V_UNCONNECTED_1490,
  SV2V_UNCONNECTED_1491,SV2V_UNCONNECTED_1492,SV2V_UNCONNECTED_1493,
  SV2V_UNCONNECTED_1494,SV2V_UNCONNECTED_1495,SV2V_UNCONNECTED_1496,SV2V_UNCONNECTED_1497,
  SV2V_UNCONNECTED_1498,SV2V_UNCONNECTED_1499,SV2V_UNCONNECTED_1500,
  SV2V_UNCONNECTED_1501,SV2V_UNCONNECTED_1502,SV2V_UNCONNECTED_1503,
  SV2V_UNCONNECTED_1504,SV2V_UNCONNECTED_1505,SV2V_UNCONNECTED_1506,
  SV2V_UNCONNECTED_1507,SV2V_UNCONNECTED_1508,SV2V_UNCONNECTED_1509,
  SV2V_UNCONNECTED_1510,SV2V_UNCONNECTED_1511,SV2V_UNCONNECTED_1512,
  SV2V_UNCONNECTED_1513,SV2V_UNCONNECTED_1514,SV2V_UNCONNECTED_1515,
  SV2V_UNCONNECTED_1516,SV2V_UNCONNECTED_1517,SV2V_UNCONNECTED_1518,
  SV2V_UNCONNECTED_1519,SV2V_UNCONNECTED_1520,SV2V_UNCONNECTED_1521,
  SV2V_UNCONNECTED_1522,SV2V_UNCONNECTED_1523,SV2V_UNCONNECTED_1524,
  SV2V_UNCONNECTED_1525,SV2V_UNCONNECTED_1526,SV2V_UNCONNECTED_1527,
  SV2V_UNCONNECTED_1528,SV2V_UNCONNECTED_1529,SV2V_UNCONNECTED_1530,
  SV2V_UNCONNECTED_1531,SV2V_UNCONNECTED_1532,SV2V_UNCONNECTED_1533,
  SV2V_UNCONNECTED_1534,SV2V_UNCONNECTED_1535,SV2V_UNCONNECTED_1536,SV2V_UNCONNECTED_1537,
  SV2V_UNCONNECTED_1538,SV2V_UNCONNECTED_1539,SV2V_UNCONNECTED_1540,
  SV2V_UNCONNECTED_1541,SV2V_UNCONNECTED_1542,SV2V_UNCONNECTED_1543,
  SV2V_UNCONNECTED_1544,SV2V_UNCONNECTED_1545,SV2V_UNCONNECTED_1546,
  SV2V_UNCONNECTED_1547,SV2V_UNCONNECTED_1548,SV2V_UNCONNECTED_1549,
  SV2V_UNCONNECTED_1550,SV2V_UNCONNECTED_1551,SV2V_UNCONNECTED_1552,
  SV2V_UNCONNECTED_1553,SV2V_UNCONNECTED_1554,SV2V_UNCONNECTED_1555,
  SV2V_UNCONNECTED_1556,SV2V_UNCONNECTED_1557,SV2V_UNCONNECTED_1558,
  SV2V_UNCONNECTED_1559,SV2V_UNCONNECTED_1560,SV2V_UNCONNECTED_1561,
  SV2V_UNCONNECTED_1562,SV2V_UNCONNECTED_1563,SV2V_UNCONNECTED_1564,
  SV2V_UNCONNECTED_1565,SV2V_UNCONNECTED_1566,SV2V_UNCONNECTED_1567,
  SV2V_UNCONNECTED_1568,SV2V_UNCONNECTED_1569,SV2V_UNCONNECTED_1570,
  SV2V_UNCONNECTED_1571,SV2V_UNCONNECTED_1572,SV2V_UNCONNECTED_1573,
  SV2V_UNCONNECTED_1574,SV2V_UNCONNECTED_1575,SV2V_UNCONNECTED_1576,SV2V_UNCONNECTED_1577,
  SV2V_UNCONNECTED_1578,SV2V_UNCONNECTED_1579,SV2V_UNCONNECTED_1580,
  SV2V_UNCONNECTED_1581,SV2V_UNCONNECTED_1582,SV2V_UNCONNECTED_1583,
  SV2V_UNCONNECTED_1584,SV2V_UNCONNECTED_1585,SV2V_UNCONNECTED_1586,
  SV2V_UNCONNECTED_1587,SV2V_UNCONNECTED_1588,SV2V_UNCONNECTED_1589,
  SV2V_UNCONNECTED_1590,SV2V_UNCONNECTED_1591,SV2V_UNCONNECTED_1592,
  SV2V_UNCONNECTED_1593,SV2V_UNCONNECTED_1594,SV2V_UNCONNECTED_1595,
  SV2V_UNCONNECTED_1596,SV2V_UNCONNECTED_1597,SV2V_UNCONNECTED_1598,
  SV2V_UNCONNECTED_1599,SV2V_UNCONNECTED_1600,SV2V_UNCONNECTED_1601,
  SV2V_UNCONNECTED_1602,SV2V_UNCONNECTED_1603,SV2V_UNCONNECTED_1604,
  SV2V_UNCONNECTED_1605,SV2V_UNCONNECTED_1606,SV2V_UNCONNECTED_1607,
  SV2V_UNCONNECTED_1608,SV2V_UNCONNECTED_1609,SV2V_UNCONNECTED_1610,
  SV2V_UNCONNECTED_1611,SV2V_UNCONNECTED_1612,SV2V_UNCONNECTED_1613,
  SV2V_UNCONNECTED_1614,SV2V_UNCONNECTED_1615,SV2V_UNCONNECTED_1616,SV2V_UNCONNECTED_1617,
  SV2V_UNCONNECTED_1618,SV2V_UNCONNECTED_1619,SV2V_UNCONNECTED_1620,
  SV2V_UNCONNECTED_1621,SV2V_UNCONNECTED_1622,SV2V_UNCONNECTED_1623,
  SV2V_UNCONNECTED_1624,SV2V_UNCONNECTED_1625,SV2V_UNCONNECTED_1626,
  SV2V_UNCONNECTED_1627,SV2V_UNCONNECTED_1628,SV2V_UNCONNECTED_1629,
  SV2V_UNCONNECTED_1630,SV2V_UNCONNECTED_1631,SV2V_UNCONNECTED_1632,
  SV2V_UNCONNECTED_1633,SV2V_UNCONNECTED_1634,SV2V_UNCONNECTED_1635,
  SV2V_UNCONNECTED_1636,SV2V_UNCONNECTED_1637,SV2V_UNCONNECTED_1638,
  SV2V_UNCONNECTED_1639,SV2V_UNCONNECTED_1640,SV2V_UNCONNECTED_1641,
  SV2V_UNCONNECTED_1642,SV2V_UNCONNECTED_1643,SV2V_UNCONNECTED_1644,
  SV2V_UNCONNECTED_1645,SV2V_UNCONNECTED_1646,SV2V_UNCONNECTED_1647,
  SV2V_UNCONNECTED_1648,SV2V_UNCONNECTED_1649,SV2V_UNCONNECTED_1650,
  SV2V_UNCONNECTED_1651,SV2V_UNCONNECTED_1652,SV2V_UNCONNECTED_1653,
  SV2V_UNCONNECTED_1654,SV2V_UNCONNECTED_1655,SV2V_UNCONNECTED_1656,SV2V_UNCONNECTED_1657,
  SV2V_UNCONNECTED_1658,SV2V_UNCONNECTED_1659,SV2V_UNCONNECTED_1660,
  SV2V_UNCONNECTED_1661,SV2V_UNCONNECTED_1662,SV2V_UNCONNECTED_1663,
  SV2V_UNCONNECTED_1664,SV2V_UNCONNECTED_1665,SV2V_UNCONNECTED_1666,
  SV2V_UNCONNECTED_1667,SV2V_UNCONNECTED_1668,SV2V_UNCONNECTED_1669,
  SV2V_UNCONNECTED_1670,SV2V_UNCONNECTED_1671,SV2V_UNCONNECTED_1672,
  SV2V_UNCONNECTED_1673,SV2V_UNCONNECTED_1674,SV2V_UNCONNECTED_1675,
  SV2V_UNCONNECTED_1676,SV2V_UNCONNECTED_1677,SV2V_UNCONNECTED_1678,
  SV2V_UNCONNECTED_1679,SV2V_UNCONNECTED_1680,SV2V_UNCONNECTED_1681,
  SV2V_UNCONNECTED_1682,SV2V_UNCONNECTED_1683,SV2V_UNCONNECTED_1684,
  SV2V_UNCONNECTED_1685,SV2V_UNCONNECTED_1686,SV2V_UNCONNECTED_1687,
  SV2V_UNCONNECTED_1688,SV2V_UNCONNECTED_1689,SV2V_UNCONNECTED_1690,
  SV2V_UNCONNECTED_1691,SV2V_UNCONNECTED_1692,SV2V_UNCONNECTED_1693,
  SV2V_UNCONNECTED_1694,SV2V_UNCONNECTED_1695,SV2V_UNCONNECTED_1696,SV2V_UNCONNECTED_1697,
  SV2V_UNCONNECTED_1698,SV2V_UNCONNECTED_1699,SV2V_UNCONNECTED_1700,
  SV2V_UNCONNECTED_1701,SV2V_UNCONNECTED_1702,SV2V_UNCONNECTED_1703,
  SV2V_UNCONNECTED_1704,SV2V_UNCONNECTED_1705,SV2V_UNCONNECTED_1706,
  SV2V_UNCONNECTED_1707,SV2V_UNCONNECTED_1708,SV2V_UNCONNECTED_1709,
  SV2V_UNCONNECTED_1710,SV2V_UNCONNECTED_1711,SV2V_UNCONNECTED_1712,
  SV2V_UNCONNECTED_1713,SV2V_UNCONNECTED_1714,SV2V_UNCONNECTED_1715,
  SV2V_UNCONNECTED_1716,SV2V_UNCONNECTED_1717,SV2V_UNCONNECTED_1718,
  SV2V_UNCONNECTED_1719,SV2V_UNCONNECTED_1720,SV2V_UNCONNECTED_1721,
  SV2V_UNCONNECTED_1722,SV2V_UNCONNECTED_1723,SV2V_UNCONNECTED_1724,
  SV2V_UNCONNECTED_1725,SV2V_UNCONNECTED_1726,SV2V_UNCONNECTED_1727,
  SV2V_UNCONNECTED_1728,SV2V_UNCONNECTED_1729,SV2V_UNCONNECTED_1730,
  SV2V_UNCONNECTED_1731,SV2V_UNCONNECTED_1732,SV2V_UNCONNECTED_1733,
  SV2V_UNCONNECTED_1734,SV2V_UNCONNECTED_1735,SV2V_UNCONNECTED_1736,SV2V_UNCONNECTED_1737,
  SV2V_UNCONNECTED_1738,SV2V_UNCONNECTED_1739,SV2V_UNCONNECTED_1740,
  SV2V_UNCONNECTED_1741,SV2V_UNCONNECTED_1742,SV2V_UNCONNECTED_1743,
  SV2V_UNCONNECTED_1744,SV2V_UNCONNECTED_1745,SV2V_UNCONNECTED_1746,
  SV2V_UNCONNECTED_1747,SV2V_UNCONNECTED_1748,SV2V_UNCONNECTED_1749,
  SV2V_UNCONNECTED_1750,SV2V_UNCONNECTED_1751,SV2V_UNCONNECTED_1752,
  SV2V_UNCONNECTED_1753,SV2V_UNCONNECTED_1754,SV2V_UNCONNECTED_1755,
  SV2V_UNCONNECTED_1756,SV2V_UNCONNECTED_1757,SV2V_UNCONNECTED_1758,
  SV2V_UNCONNECTED_1759,SV2V_UNCONNECTED_1760,SV2V_UNCONNECTED_1761,
  SV2V_UNCONNECTED_1762,SV2V_UNCONNECTED_1763,SV2V_UNCONNECTED_1764,
  SV2V_UNCONNECTED_1765,SV2V_UNCONNECTED_1766,SV2V_UNCONNECTED_1767,
  SV2V_UNCONNECTED_1768,SV2V_UNCONNECTED_1769,SV2V_UNCONNECTED_1770,
  SV2V_UNCONNECTED_1771,SV2V_UNCONNECTED_1772,SV2V_UNCONNECTED_1773,
  SV2V_UNCONNECTED_1774,SV2V_UNCONNECTED_1775,SV2V_UNCONNECTED_1776,SV2V_UNCONNECTED_1777,
  SV2V_UNCONNECTED_1778,SV2V_UNCONNECTED_1779,SV2V_UNCONNECTED_1780,
  SV2V_UNCONNECTED_1781,SV2V_UNCONNECTED_1782,SV2V_UNCONNECTED_1783,
  SV2V_UNCONNECTED_1784,SV2V_UNCONNECTED_1785,SV2V_UNCONNECTED_1786,
  SV2V_UNCONNECTED_1787,SV2V_UNCONNECTED_1788,SV2V_UNCONNECTED_1789,
  SV2V_UNCONNECTED_1790,SV2V_UNCONNECTED_1791,SV2V_UNCONNECTED_1792,
  SV2V_UNCONNECTED_1793,SV2V_UNCONNECTED_1794,SV2V_UNCONNECTED_1795,
  SV2V_UNCONNECTED_1796,SV2V_UNCONNECTED_1797,SV2V_UNCONNECTED_1798,
  SV2V_UNCONNECTED_1799,SV2V_UNCONNECTED_1800,SV2V_UNCONNECTED_1801,
  SV2V_UNCONNECTED_1802,SV2V_UNCONNECTED_1803,SV2V_UNCONNECTED_1804,
  SV2V_UNCONNECTED_1805,SV2V_UNCONNECTED_1806,SV2V_UNCONNECTED_1807,
  SV2V_UNCONNECTED_1808,SV2V_UNCONNECTED_1809,SV2V_UNCONNECTED_1810,
  SV2V_UNCONNECTED_1811,SV2V_UNCONNECTED_1812,SV2V_UNCONNECTED_1813,
  SV2V_UNCONNECTED_1814,SV2V_UNCONNECTED_1815,SV2V_UNCONNECTED_1816,SV2V_UNCONNECTED_1817,
  SV2V_UNCONNECTED_1818,SV2V_UNCONNECTED_1819,SV2V_UNCONNECTED_1820,
  SV2V_UNCONNECTED_1821,SV2V_UNCONNECTED_1822,SV2V_UNCONNECTED_1823,
  SV2V_UNCONNECTED_1824,SV2V_UNCONNECTED_1825,SV2V_UNCONNECTED_1826,
  SV2V_UNCONNECTED_1827,SV2V_UNCONNECTED_1828,SV2V_UNCONNECTED_1829,
  SV2V_UNCONNECTED_1830,SV2V_UNCONNECTED_1831,SV2V_UNCONNECTED_1832,
  SV2V_UNCONNECTED_1833,SV2V_UNCONNECTED_1834,SV2V_UNCONNECTED_1835,
  SV2V_UNCONNECTED_1836,SV2V_UNCONNECTED_1837,SV2V_UNCONNECTED_1838,
  SV2V_UNCONNECTED_1839,SV2V_UNCONNECTED_1840,SV2V_UNCONNECTED_1841,
  SV2V_UNCONNECTED_1842,SV2V_UNCONNECTED_1843,SV2V_UNCONNECTED_1844,
  SV2V_UNCONNECTED_1845,SV2V_UNCONNECTED_1846,SV2V_UNCONNECTED_1847,
  SV2V_UNCONNECTED_1848,SV2V_UNCONNECTED_1849,SV2V_UNCONNECTED_1850,
  SV2V_UNCONNECTED_1851,SV2V_UNCONNECTED_1852,SV2V_UNCONNECTED_1853,
  SV2V_UNCONNECTED_1854,SV2V_UNCONNECTED_1855,SV2V_UNCONNECTED_1856,SV2V_UNCONNECTED_1857,
  SV2V_UNCONNECTED_1858,SV2V_UNCONNECTED_1859,SV2V_UNCONNECTED_1860,
  SV2V_UNCONNECTED_1861,SV2V_UNCONNECTED_1862,SV2V_UNCONNECTED_1863,
  SV2V_UNCONNECTED_1864,SV2V_UNCONNECTED_1865,SV2V_UNCONNECTED_1866,
  SV2V_UNCONNECTED_1867,SV2V_UNCONNECTED_1868,SV2V_UNCONNECTED_1869,
  SV2V_UNCONNECTED_1870,SV2V_UNCONNECTED_1871,SV2V_UNCONNECTED_1872,
  SV2V_UNCONNECTED_1873,SV2V_UNCONNECTED_1874,SV2V_UNCONNECTED_1875,
  SV2V_UNCONNECTED_1876,SV2V_UNCONNECTED_1877,SV2V_UNCONNECTED_1878,
  SV2V_UNCONNECTED_1879,SV2V_UNCONNECTED_1880,SV2V_UNCONNECTED_1881,
  SV2V_UNCONNECTED_1882,SV2V_UNCONNECTED_1883,SV2V_UNCONNECTED_1884,
  SV2V_UNCONNECTED_1885,SV2V_UNCONNECTED_1886,SV2V_UNCONNECTED_1887,
  SV2V_UNCONNECTED_1888,SV2V_UNCONNECTED_1889,SV2V_UNCONNECTED_1890,
  SV2V_UNCONNECTED_1891,SV2V_UNCONNECTED_1892,SV2V_UNCONNECTED_1893,
  SV2V_UNCONNECTED_1894,SV2V_UNCONNECTED_1895,SV2V_UNCONNECTED_1896,SV2V_UNCONNECTED_1897,
  SV2V_UNCONNECTED_1898,SV2V_UNCONNECTED_1899,SV2V_UNCONNECTED_1900,
  SV2V_UNCONNECTED_1901,SV2V_UNCONNECTED_1902,SV2V_UNCONNECTED_1903,
  SV2V_UNCONNECTED_1904,SV2V_UNCONNECTED_1905,SV2V_UNCONNECTED_1906,
  SV2V_UNCONNECTED_1907,SV2V_UNCONNECTED_1908,SV2V_UNCONNECTED_1909,
  SV2V_UNCONNECTED_1910,SV2V_UNCONNECTED_1911,SV2V_UNCONNECTED_1912,
  SV2V_UNCONNECTED_1913,SV2V_UNCONNECTED_1914,SV2V_UNCONNECTED_1915,
  SV2V_UNCONNECTED_1916,SV2V_UNCONNECTED_1917,SV2V_UNCONNECTED_1918,
  SV2V_UNCONNECTED_1919,SV2V_UNCONNECTED_1920,SV2V_UNCONNECTED_1921,
  SV2V_UNCONNECTED_1922,SV2V_UNCONNECTED_1923,SV2V_UNCONNECTED_1924,
  SV2V_UNCONNECTED_1925,SV2V_UNCONNECTED_1926,SV2V_UNCONNECTED_1927,
  SV2V_UNCONNECTED_1928,SV2V_UNCONNECTED_1929,SV2V_UNCONNECTED_1930,
  SV2V_UNCONNECTED_1931,SV2V_UNCONNECTED_1932,SV2V_UNCONNECTED_1933,
  SV2V_UNCONNECTED_1934,SV2V_UNCONNECTED_1935,SV2V_UNCONNECTED_1936,SV2V_UNCONNECTED_1937,
  SV2V_UNCONNECTED_1938,SV2V_UNCONNECTED_1939,SV2V_UNCONNECTED_1940,
  SV2V_UNCONNECTED_1941,SV2V_UNCONNECTED_1942,SV2V_UNCONNECTED_1943,
  SV2V_UNCONNECTED_1944,SV2V_UNCONNECTED_1945,SV2V_UNCONNECTED_1946,
  SV2V_UNCONNECTED_1947,SV2V_UNCONNECTED_1948,SV2V_UNCONNECTED_1949,
  SV2V_UNCONNECTED_1950,SV2V_UNCONNECTED_1951,SV2V_UNCONNECTED_1952,
  SV2V_UNCONNECTED_1953,SV2V_UNCONNECTED_1954,SV2V_UNCONNECTED_1955,
  SV2V_UNCONNECTED_1956,SV2V_UNCONNECTED_1957,SV2V_UNCONNECTED_1958,
  SV2V_UNCONNECTED_1959,SV2V_UNCONNECTED_1960,SV2V_UNCONNECTED_1961,
  SV2V_UNCONNECTED_1962,SV2V_UNCONNECTED_1963,SV2V_UNCONNECTED_1964,
  SV2V_UNCONNECTED_1965,SV2V_UNCONNECTED_1966,SV2V_UNCONNECTED_1967,
  SV2V_UNCONNECTED_1968,SV2V_UNCONNECTED_1969,SV2V_UNCONNECTED_1970,
  SV2V_UNCONNECTED_1971,SV2V_UNCONNECTED_1972,SV2V_UNCONNECTED_1973,
  SV2V_UNCONNECTED_1974,SV2V_UNCONNECTED_1975,SV2V_UNCONNECTED_1976,SV2V_UNCONNECTED_1977,
  SV2V_UNCONNECTED_1978,SV2V_UNCONNECTED_1979,SV2V_UNCONNECTED_1980,
  SV2V_UNCONNECTED_1981,SV2V_UNCONNECTED_1982,SV2V_UNCONNECTED_1983,
  SV2V_UNCONNECTED_1984,SV2V_UNCONNECTED_1985,SV2V_UNCONNECTED_1986,
  SV2V_UNCONNECTED_1987,SV2V_UNCONNECTED_1988,SV2V_UNCONNECTED_1989,
  SV2V_UNCONNECTED_1990,SV2V_UNCONNECTED_1991,SV2V_UNCONNECTED_1992,
  SV2V_UNCONNECTED_1993,SV2V_UNCONNECTED_1994,SV2V_UNCONNECTED_1995,
  SV2V_UNCONNECTED_1996,SV2V_UNCONNECTED_1997,SV2V_UNCONNECTED_1998,
  SV2V_UNCONNECTED_1999,SV2V_UNCONNECTED_2000,SV2V_UNCONNECTED_2001,
  SV2V_UNCONNECTED_2002,SV2V_UNCONNECTED_2003,SV2V_UNCONNECTED_2004,
  SV2V_UNCONNECTED_2005,SV2V_UNCONNECTED_2006,SV2V_UNCONNECTED_2007,
  SV2V_UNCONNECTED_2008,SV2V_UNCONNECTED_2009,SV2V_UNCONNECTED_2010,
  SV2V_UNCONNECTED_2011,SV2V_UNCONNECTED_2012,SV2V_UNCONNECTED_2013,
  SV2V_UNCONNECTED_2014,SV2V_UNCONNECTED_2015,SV2V_UNCONNECTED_2016,SV2V_UNCONNECTED_2017,
  SV2V_UNCONNECTED_2018,SV2V_UNCONNECTED_2019,SV2V_UNCONNECTED_2020,
  SV2V_UNCONNECTED_2021,SV2V_UNCONNECTED_2022,SV2V_UNCONNECTED_2023,
  SV2V_UNCONNECTED_2024,SV2V_UNCONNECTED_2025,SV2V_UNCONNECTED_2026,
  SV2V_UNCONNECTED_2027,SV2V_UNCONNECTED_2028,SV2V_UNCONNECTED_2029,
  SV2V_UNCONNECTED_2030,SV2V_UNCONNECTED_2031,SV2V_UNCONNECTED_2032,
  SV2V_UNCONNECTED_2033,SV2V_UNCONNECTED_2034,SV2V_UNCONNECTED_2035,
  SV2V_UNCONNECTED_2036,SV2V_UNCONNECTED_2037,SV2V_UNCONNECTED_2038,
  SV2V_UNCONNECTED_2039,SV2V_UNCONNECTED_2040,SV2V_UNCONNECTED_2041,
  SV2V_UNCONNECTED_2042,SV2V_UNCONNECTED_2043,SV2V_UNCONNECTED_2044,
  SV2V_UNCONNECTED_2045,SV2V_UNCONNECTED_2046,SV2V_UNCONNECTED_2047,
  SV2V_UNCONNECTED_2048,SV2V_UNCONNECTED_2049,SV2V_UNCONNECTED_2050,
  SV2V_UNCONNECTED_2051,SV2V_UNCONNECTED_2052,SV2V_UNCONNECTED_2053,
  SV2V_UNCONNECTED_2054,SV2V_UNCONNECTED_2055,SV2V_UNCONNECTED_2056,SV2V_UNCONNECTED_2057,
  SV2V_UNCONNECTED_2058,SV2V_UNCONNECTED_2059,SV2V_UNCONNECTED_2060,
  SV2V_UNCONNECTED_2061,SV2V_UNCONNECTED_2062,SV2V_UNCONNECTED_2063,
  SV2V_UNCONNECTED_2064,SV2V_UNCONNECTED_2065,SV2V_UNCONNECTED_2066,
  SV2V_UNCONNECTED_2067,SV2V_UNCONNECTED_2068,SV2V_UNCONNECTED_2069,
  SV2V_UNCONNECTED_2070,SV2V_UNCONNECTED_2071,SV2V_UNCONNECTED_2072,
  SV2V_UNCONNECTED_2073,SV2V_UNCONNECTED_2074,SV2V_UNCONNECTED_2075,
  SV2V_UNCONNECTED_2076,SV2V_UNCONNECTED_2077,SV2V_UNCONNECTED_2078,
  SV2V_UNCONNECTED_2079,SV2V_UNCONNECTED_2080,SV2V_UNCONNECTED_2081,
  SV2V_UNCONNECTED_2082,SV2V_UNCONNECTED_2083,SV2V_UNCONNECTED_2084,
  SV2V_UNCONNECTED_2085,SV2V_UNCONNECTED_2086,SV2V_UNCONNECTED_2087,
  SV2V_UNCONNECTED_2088,SV2V_UNCONNECTED_2089,SV2V_UNCONNECTED_2090,
  SV2V_UNCONNECTED_2091,SV2V_UNCONNECTED_2092,SV2V_UNCONNECTED_2093,
  SV2V_UNCONNECTED_2094,SV2V_UNCONNECTED_2095,SV2V_UNCONNECTED_2096,SV2V_UNCONNECTED_2097,
  SV2V_UNCONNECTED_2098,SV2V_UNCONNECTED_2099,SV2V_UNCONNECTED_2100,
  SV2V_UNCONNECTED_2101,SV2V_UNCONNECTED_2102,SV2V_UNCONNECTED_2103,
  SV2V_UNCONNECTED_2104,SV2V_UNCONNECTED_2105,SV2V_UNCONNECTED_2106,
  SV2V_UNCONNECTED_2107,SV2V_UNCONNECTED_2108,SV2V_UNCONNECTED_2109,
  SV2V_UNCONNECTED_2110,SV2V_UNCONNECTED_2111,SV2V_UNCONNECTED_2112,
  SV2V_UNCONNECTED_2113,SV2V_UNCONNECTED_2114,SV2V_UNCONNECTED_2115,
  SV2V_UNCONNECTED_2116,SV2V_UNCONNECTED_2117,SV2V_UNCONNECTED_2118,
  SV2V_UNCONNECTED_2119,SV2V_UNCONNECTED_2120,SV2V_UNCONNECTED_2121,
  SV2V_UNCONNECTED_2122,SV2V_UNCONNECTED_2123,SV2V_UNCONNECTED_2124,
  SV2V_UNCONNECTED_2125,SV2V_UNCONNECTED_2126,SV2V_UNCONNECTED_2127,
  SV2V_UNCONNECTED_2128,SV2V_UNCONNECTED_2129,SV2V_UNCONNECTED_2130,
  SV2V_UNCONNECTED_2131,SV2V_UNCONNECTED_2132,SV2V_UNCONNECTED_2133,
  SV2V_UNCONNECTED_2134,SV2V_UNCONNECTED_2135,SV2V_UNCONNECTED_2136,SV2V_UNCONNECTED_2137,
  SV2V_UNCONNECTED_2138,SV2V_UNCONNECTED_2139,SV2V_UNCONNECTED_2140,
  SV2V_UNCONNECTED_2141,SV2V_UNCONNECTED_2142,SV2V_UNCONNECTED_2143,
  SV2V_UNCONNECTED_2144,SV2V_UNCONNECTED_2145,SV2V_UNCONNECTED_2146,
  SV2V_UNCONNECTED_2147,SV2V_UNCONNECTED_2148,SV2V_UNCONNECTED_2149,
  SV2V_UNCONNECTED_2150,SV2V_UNCONNECTED_2151,SV2V_UNCONNECTED_2152,
  SV2V_UNCONNECTED_2153,SV2V_UNCONNECTED_2154,SV2V_UNCONNECTED_2155,
  SV2V_UNCONNECTED_2156,SV2V_UNCONNECTED_2157,SV2V_UNCONNECTED_2158,
  SV2V_UNCONNECTED_2159,SV2V_UNCONNECTED_2160,SV2V_UNCONNECTED_2161,
  SV2V_UNCONNECTED_2162,SV2V_UNCONNECTED_2163,SV2V_UNCONNECTED_2164,
  SV2V_UNCONNECTED_2165,SV2V_UNCONNECTED_2166,SV2V_UNCONNECTED_2167,
  SV2V_UNCONNECTED_2168,SV2V_UNCONNECTED_2169,SV2V_UNCONNECTED_2170,
  SV2V_UNCONNECTED_2171,SV2V_UNCONNECTED_2172,SV2V_UNCONNECTED_2173,
  SV2V_UNCONNECTED_2174,SV2V_UNCONNECTED_2175,SV2V_UNCONNECTED_2176,SV2V_UNCONNECTED_2177,
  SV2V_UNCONNECTED_2178,SV2V_UNCONNECTED_2179,SV2V_UNCONNECTED_2180,
  SV2V_UNCONNECTED_2181,SV2V_UNCONNECTED_2182,SV2V_UNCONNECTED_2183,
  SV2V_UNCONNECTED_2184,SV2V_UNCONNECTED_2185,SV2V_UNCONNECTED_2186,
  SV2V_UNCONNECTED_2187,SV2V_UNCONNECTED_2188,SV2V_UNCONNECTED_2189,
  SV2V_UNCONNECTED_2190,SV2V_UNCONNECTED_2191,SV2V_UNCONNECTED_2192,
  SV2V_UNCONNECTED_2193,SV2V_UNCONNECTED_2194,SV2V_UNCONNECTED_2195,
  SV2V_UNCONNECTED_2196,SV2V_UNCONNECTED_2197,SV2V_UNCONNECTED_2198,
  SV2V_UNCONNECTED_2199,SV2V_UNCONNECTED_2200,SV2V_UNCONNECTED_2201,
  SV2V_UNCONNECTED_2202,SV2V_UNCONNECTED_2203,SV2V_UNCONNECTED_2204,
  SV2V_UNCONNECTED_2205,SV2V_UNCONNECTED_2206,SV2V_UNCONNECTED_2207,
  SV2V_UNCONNECTED_2208,SV2V_UNCONNECTED_2209,SV2V_UNCONNECTED_2210,
  SV2V_UNCONNECTED_2211,SV2V_UNCONNECTED_2212,SV2V_UNCONNECTED_2213,
  SV2V_UNCONNECTED_2214,SV2V_UNCONNECTED_2215,SV2V_UNCONNECTED_2216,SV2V_UNCONNECTED_2217,
  SV2V_UNCONNECTED_2218,SV2V_UNCONNECTED_2219,SV2V_UNCONNECTED_2220,
  SV2V_UNCONNECTED_2221,SV2V_UNCONNECTED_2222,SV2V_UNCONNECTED_2223,
  SV2V_UNCONNECTED_2224,SV2V_UNCONNECTED_2225,SV2V_UNCONNECTED_2226,
  SV2V_UNCONNECTED_2227,SV2V_UNCONNECTED_2228,SV2V_UNCONNECTED_2229,
  SV2V_UNCONNECTED_2230,SV2V_UNCONNECTED_2231,SV2V_UNCONNECTED_2232,
  SV2V_UNCONNECTED_2233,SV2V_UNCONNECTED_2234,SV2V_UNCONNECTED_2235,
  SV2V_UNCONNECTED_2236,SV2V_UNCONNECTED_2237,SV2V_UNCONNECTED_2238,
  SV2V_UNCONNECTED_2239,SV2V_UNCONNECTED_2240,SV2V_UNCONNECTED_2241,
  SV2V_UNCONNECTED_2242,SV2V_UNCONNECTED_2243,SV2V_UNCONNECTED_2244,
  SV2V_UNCONNECTED_2245,SV2V_UNCONNECTED_2246,SV2V_UNCONNECTED_2247,
  SV2V_UNCONNECTED_2248,SV2V_UNCONNECTED_2249,SV2V_UNCONNECTED_2250,
  SV2V_UNCONNECTED_2251,SV2V_UNCONNECTED_2252,SV2V_UNCONNECTED_2253,
  SV2V_UNCONNECTED_2254,SV2V_UNCONNECTED_2255,SV2V_UNCONNECTED_2256,SV2V_UNCONNECTED_2257,
  SV2V_UNCONNECTED_2258,SV2V_UNCONNECTED_2259,SV2V_UNCONNECTED_2260,
  SV2V_UNCONNECTED_2261,SV2V_UNCONNECTED_2262,SV2V_UNCONNECTED_2263,
  SV2V_UNCONNECTED_2264,SV2V_UNCONNECTED_2265,SV2V_UNCONNECTED_2266,
  SV2V_UNCONNECTED_2267,SV2V_UNCONNECTED_2268,SV2V_UNCONNECTED_2269,
  SV2V_UNCONNECTED_2270,SV2V_UNCONNECTED_2271,SV2V_UNCONNECTED_2272,
  SV2V_UNCONNECTED_2273,SV2V_UNCONNECTED_2274,SV2V_UNCONNECTED_2275,
  SV2V_UNCONNECTED_2276,SV2V_UNCONNECTED_2277,SV2V_UNCONNECTED_2278,
  SV2V_UNCONNECTED_2279,SV2V_UNCONNECTED_2280,SV2V_UNCONNECTED_2281,
  SV2V_UNCONNECTED_2282,SV2V_UNCONNECTED_2283,SV2V_UNCONNECTED_2284,
  SV2V_UNCONNECTED_2285,SV2V_UNCONNECTED_2286,SV2V_UNCONNECTED_2287,
  SV2V_UNCONNECTED_2288,SV2V_UNCONNECTED_2289,SV2V_UNCONNECTED_2290,
  SV2V_UNCONNECTED_2291,SV2V_UNCONNECTED_2292,SV2V_UNCONNECTED_2293,
  SV2V_UNCONNECTED_2294,SV2V_UNCONNECTED_2295,SV2V_UNCONNECTED_2296,SV2V_UNCONNECTED_2297,
  SV2V_UNCONNECTED_2298,SV2V_UNCONNECTED_2299,SV2V_UNCONNECTED_2300,
  SV2V_UNCONNECTED_2301,SV2V_UNCONNECTED_2302,SV2V_UNCONNECTED_2303,
  SV2V_UNCONNECTED_2304,SV2V_UNCONNECTED_2305,SV2V_UNCONNECTED_2306,
  SV2V_UNCONNECTED_2307,SV2V_UNCONNECTED_2308,SV2V_UNCONNECTED_2309,
  SV2V_UNCONNECTED_2310,SV2V_UNCONNECTED_2311,SV2V_UNCONNECTED_2312,
  SV2V_UNCONNECTED_2313,SV2V_UNCONNECTED_2314,SV2V_UNCONNECTED_2315,
  SV2V_UNCONNECTED_2316,SV2V_UNCONNECTED_2317,SV2V_UNCONNECTED_2318,
  SV2V_UNCONNECTED_2319,SV2V_UNCONNECTED_2320,SV2V_UNCONNECTED_2321,
  SV2V_UNCONNECTED_2322,SV2V_UNCONNECTED_2323,SV2V_UNCONNECTED_2324,
  SV2V_UNCONNECTED_2325,SV2V_UNCONNECTED_2326,SV2V_UNCONNECTED_2327,
  SV2V_UNCONNECTED_2328,SV2V_UNCONNECTED_2329,SV2V_UNCONNECTED_2330,
  SV2V_UNCONNECTED_2331,SV2V_UNCONNECTED_2332,SV2V_UNCONNECTED_2333,
  SV2V_UNCONNECTED_2334,SV2V_UNCONNECTED_2335,SV2V_UNCONNECTED_2336,SV2V_UNCONNECTED_2337,
  SV2V_UNCONNECTED_2338,SV2V_UNCONNECTED_2339,SV2V_UNCONNECTED_2340,
  SV2V_UNCONNECTED_2341,SV2V_UNCONNECTED_2342,SV2V_UNCONNECTED_2343,
  SV2V_UNCONNECTED_2344,SV2V_UNCONNECTED_2345,SV2V_UNCONNECTED_2346,
  SV2V_UNCONNECTED_2347,SV2V_UNCONNECTED_2348,SV2V_UNCONNECTED_2349,
  SV2V_UNCONNECTED_2350,SV2V_UNCONNECTED_2351,SV2V_UNCONNECTED_2352,
  SV2V_UNCONNECTED_2353,SV2V_UNCONNECTED_2354,SV2V_UNCONNECTED_2355,
  SV2V_UNCONNECTED_2356,SV2V_UNCONNECTED_2357,SV2V_UNCONNECTED_2358,
  SV2V_UNCONNECTED_2359,SV2V_UNCONNECTED_2360,SV2V_UNCONNECTED_2361,
  SV2V_UNCONNECTED_2362,SV2V_UNCONNECTED_2363,SV2V_UNCONNECTED_2364,
  SV2V_UNCONNECTED_2365,SV2V_UNCONNECTED_2366,SV2V_UNCONNECTED_2367,
  SV2V_UNCONNECTED_2368,SV2V_UNCONNECTED_2369,SV2V_UNCONNECTED_2370,
  SV2V_UNCONNECTED_2371,SV2V_UNCONNECTED_2372,SV2V_UNCONNECTED_2373,
  SV2V_UNCONNECTED_2374,SV2V_UNCONNECTED_2375,SV2V_UNCONNECTED_2376,SV2V_UNCONNECTED_2377,
  SV2V_UNCONNECTED_2378,SV2V_UNCONNECTED_2379,SV2V_UNCONNECTED_2380,
  SV2V_UNCONNECTED_2381,SV2V_UNCONNECTED_2382,SV2V_UNCONNECTED_2383,
  SV2V_UNCONNECTED_2384,SV2V_UNCONNECTED_2385,SV2V_UNCONNECTED_2386,
  SV2V_UNCONNECTED_2387,SV2V_UNCONNECTED_2388,SV2V_UNCONNECTED_2389,
  SV2V_UNCONNECTED_2390,SV2V_UNCONNECTED_2391,SV2V_UNCONNECTED_2392,
  SV2V_UNCONNECTED_2393,SV2V_UNCONNECTED_2394,SV2V_UNCONNECTED_2395,
  SV2V_UNCONNECTED_2396,SV2V_UNCONNECTED_2397,SV2V_UNCONNECTED_2398,
  SV2V_UNCONNECTED_2399,SV2V_UNCONNECTED_2400,SV2V_UNCONNECTED_2401,
  SV2V_UNCONNECTED_2402,SV2V_UNCONNECTED_2403,SV2V_UNCONNECTED_2404,
  SV2V_UNCONNECTED_2405,SV2V_UNCONNECTED_2406,SV2V_UNCONNECTED_2407,
  SV2V_UNCONNECTED_2408,SV2V_UNCONNECTED_2409,SV2V_UNCONNECTED_2410,
  SV2V_UNCONNECTED_2411,SV2V_UNCONNECTED_2412,SV2V_UNCONNECTED_2413,
  SV2V_UNCONNECTED_2414,SV2V_UNCONNECTED_2415,SV2V_UNCONNECTED_2416,SV2V_UNCONNECTED_2417,
  SV2V_UNCONNECTED_2418,SV2V_UNCONNECTED_2419,SV2V_UNCONNECTED_2420,
  SV2V_UNCONNECTED_2421,SV2V_UNCONNECTED_2422,SV2V_UNCONNECTED_2423,
  SV2V_UNCONNECTED_2424,SV2V_UNCONNECTED_2425,SV2V_UNCONNECTED_2426,
  SV2V_UNCONNECTED_2427,SV2V_UNCONNECTED_2428,SV2V_UNCONNECTED_2429,
  SV2V_UNCONNECTED_2430,SV2V_UNCONNECTED_2431,SV2V_UNCONNECTED_2432,
  SV2V_UNCONNECTED_2433,SV2V_UNCONNECTED_2434,SV2V_UNCONNECTED_2435,
  SV2V_UNCONNECTED_2436,SV2V_UNCONNECTED_2437,SV2V_UNCONNECTED_2438,
  SV2V_UNCONNECTED_2439,SV2V_UNCONNECTED_2440,SV2V_UNCONNECTED_2441,
  SV2V_UNCONNECTED_2442,SV2V_UNCONNECTED_2443,SV2V_UNCONNECTED_2444,
  SV2V_UNCONNECTED_2445,SV2V_UNCONNECTED_2446,SV2V_UNCONNECTED_2447,
  SV2V_UNCONNECTED_2448,SV2V_UNCONNECTED_2449,SV2V_UNCONNECTED_2450,
  SV2V_UNCONNECTED_2451,SV2V_UNCONNECTED_2452,SV2V_UNCONNECTED_2453,
  SV2V_UNCONNECTED_2454,SV2V_UNCONNECTED_2455,SV2V_UNCONNECTED_2456,SV2V_UNCONNECTED_2457,
  SV2V_UNCONNECTED_2458,SV2V_UNCONNECTED_2459,SV2V_UNCONNECTED_2460,
  SV2V_UNCONNECTED_2461,SV2V_UNCONNECTED_2462,SV2V_UNCONNECTED_2463,
  SV2V_UNCONNECTED_2464,SV2V_UNCONNECTED_2465,SV2V_UNCONNECTED_2466,
  SV2V_UNCONNECTED_2467,SV2V_UNCONNECTED_2468,SV2V_UNCONNECTED_2469,
  SV2V_UNCONNECTED_2470,SV2V_UNCONNECTED_2471,SV2V_UNCONNECTED_2472,
  SV2V_UNCONNECTED_2473,SV2V_UNCONNECTED_2474,SV2V_UNCONNECTED_2475,
  SV2V_UNCONNECTED_2476,SV2V_UNCONNECTED_2477,SV2V_UNCONNECTED_2478,
  SV2V_UNCONNECTED_2479,SV2V_UNCONNECTED_2480,SV2V_UNCONNECTED_2481,
  SV2V_UNCONNECTED_2482,SV2V_UNCONNECTED_2483,SV2V_UNCONNECTED_2484,
  SV2V_UNCONNECTED_2485,SV2V_UNCONNECTED_2486,SV2V_UNCONNECTED_2487,
  SV2V_UNCONNECTED_2488,SV2V_UNCONNECTED_2489,SV2V_UNCONNECTED_2490,
  SV2V_UNCONNECTED_2491,SV2V_UNCONNECTED_2492,SV2V_UNCONNECTED_2493,
  SV2V_UNCONNECTED_2494,SV2V_UNCONNECTED_2495,SV2V_UNCONNECTED_2496,SV2V_UNCONNECTED_2497,
  SV2V_UNCONNECTED_2498,SV2V_UNCONNECTED_2499,SV2V_UNCONNECTED_2500,
  SV2V_UNCONNECTED_2501,SV2V_UNCONNECTED_2502,SV2V_UNCONNECTED_2503,
  SV2V_UNCONNECTED_2504,SV2V_UNCONNECTED_2505,SV2V_UNCONNECTED_2506,
  SV2V_UNCONNECTED_2507,SV2V_UNCONNECTED_2508,SV2V_UNCONNECTED_2509,
  SV2V_UNCONNECTED_2510,SV2V_UNCONNECTED_2511,SV2V_UNCONNECTED_2512,
  SV2V_UNCONNECTED_2513,SV2V_UNCONNECTED_2514,SV2V_UNCONNECTED_2515,
  SV2V_UNCONNECTED_2516,SV2V_UNCONNECTED_2517,SV2V_UNCONNECTED_2518,
  SV2V_UNCONNECTED_2519,SV2V_UNCONNECTED_2520,SV2V_UNCONNECTED_2521,
  SV2V_UNCONNECTED_2522,SV2V_UNCONNECTED_2523,SV2V_UNCONNECTED_2524,
  SV2V_UNCONNECTED_2525,SV2V_UNCONNECTED_2526,SV2V_UNCONNECTED_2527,
  SV2V_UNCONNECTED_2528,SV2V_UNCONNECTED_2529,SV2V_UNCONNECTED_2530,
  SV2V_UNCONNECTED_2531,SV2V_UNCONNECTED_2532,SV2V_UNCONNECTED_2533,
  SV2V_UNCONNECTED_2534,SV2V_UNCONNECTED_2535,SV2V_UNCONNECTED_2536,SV2V_UNCONNECTED_2537,
  SV2V_UNCONNECTED_2538,SV2V_UNCONNECTED_2539,SV2V_UNCONNECTED_2540,
  SV2V_UNCONNECTED_2541,SV2V_UNCONNECTED_2542,SV2V_UNCONNECTED_2543,
  SV2V_UNCONNECTED_2544,SV2V_UNCONNECTED_2545,SV2V_UNCONNECTED_2546,
  SV2V_UNCONNECTED_2547,SV2V_UNCONNECTED_2548,SV2V_UNCONNECTED_2549,
  SV2V_UNCONNECTED_2550,SV2V_UNCONNECTED_2551,SV2V_UNCONNECTED_2552,
  SV2V_UNCONNECTED_2553,SV2V_UNCONNECTED_2554,SV2V_UNCONNECTED_2555,
  SV2V_UNCONNECTED_2556,SV2V_UNCONNECTED_2557,SV2V_UNCONNECTED_2558,
  SV2V_UNCONNECTED_2559,SV2V_UNCONNECTED_2560,SV2V_UNCONNECTED_2561,
  SV2V_UNCONNECTED_2562,SV2V_UNCONNECTED_2563,SV2V_UNCONNECTED_2564,
  SV2V_UNCONNECTED_2565,SV2V_UNCONNECTED_2566,SV2V_UNCONNECTED_2567,
  SV2V_UNCONNECTED_2568,SV2V_UNCONNECTED_2569,SV2V_UNCONNECTED_2570,
  SV2V_UNCONNECTED_2571,SV2V_UNCONNECTED_2572,SV2V_UNCONNECTED_2573,
  SV2V_UNCONNECTED_2574,SV2V_UNCONNECTED_2575,SV2V_UNCONNECTED_2576,SV2V_UNCONNECTED_2577,
  SV2V_UNCONNECTED_2578,SV2V_UNCONNECTED_2579,SV2V_UNCONNECTED_2580,
  SV2V_UNCONNECTED_2581,SV2V_UNCONNECTED_2582,SV2V_UNCONNECTED_2583,
  SV2V_UNCONNECTED_2584,SV2V_UNCONNECTED_2585,SV2V_UNCONNECTED_2586,
  SV2V_UNCONNECTED_2587,SV2V_UNCONNECTED_2588,SV2V_UNCONNECTED_2589,
  SV2V_UNCONNECTED_2590,SV2V_UNCONNECTED_2591,SV2V_UNCONNECTED_2592,
  SV2V_UNCONNECTED_2593,SV2V_UNCONNECTED_2594,SV2V_UNCONNECTED_2595,
  SV2V_UNCONNECTED_2596,SV2V_UNCONNECTED_2597,SV2V_UNCONNECTED_2598,
  SV2V_UNCONNECTED_2599,SV2V_UNCONNECTED_2600,SV2V_UNCONNECTED_2601,
  SV2V_UNCONNECTED_2602,SV2V_UNCONNECTED_2603,SV2V_UNCONNECTED_2604,
  SV2V_UNCONNECTED_2605,SV2V_UNCONNECTED_2606,SV2V_UNCONNECTED_2607,
  SV2V_UNCONNECTED_2608,SV2V_UNCONNECTED_2609,SV2V_UNCONNECTED_2610,
  SV2V_UNCONNECTED_2611,SV2V_UNCONNECTED_2612,SV2V_UNCONNECTED_2613,
  SV2V_UNCONNECTED_2614,SV2V_UNCONNECTED_2615,SV2V_UNCONNECTED_2616,SV2V_UNCONNECTED_2617,
  SV2V_UNCONNECTED_2618,SV2V_UNCONNECTED_2619,SV2V_UNCONNECTED_2620,
  SV2V_UNCONNECTED_2621,SV2V_UNCONNECTED_2622,SV2V_UNCONNECTED_2623,
  SV2V_UNCONNECTED_2624,SV2V_UNCONNECTED_2625,SV2V_UNCONNECTED_2626,
  SV2V_UNCONNECTED_2627,SV2V_UNCONNECTED_2628,SV2V_UNCONNECTED_2629,
  SV2V_UNCONNECTED_2630,SV2V_UNCONNECTED_2631,SV2V_UNCONNECTED_2632,
  SV2V_UNCONNECTED_2633,SV2V_UNCONNECTED_2634,SV2V_UNCONNECTED_2635,
  SV2V_UNCONNECTED_2636,SV2V_UNCONNECTED_2637,SV2V_UNCONNECTED_2638,
  SV2V_UNCONNECTED_2639,SV2V_UNCONNECTED_2640,SV2V_UNCONNECTED_2641,
  SV2V_UNCONNECTED_2642,SV2V_UNCONNECTED_2643,SV2V_UNCONNECTED_2644,
  SV2V_UNCONNECTED_2645,SV2V_UNCONNECTED_2646,SV2V_UNCONNECTED_2647,
  SV2V_UNCONNECTED_2648,SV2V_UNCONNECTED_2649,SV2V_UNCONNECTED_2650,
  SV2V_UNCONNECTED_2651,SV2V_UNCONNECTED_2652,SV2V_UNCONNECTED_2653,
  SV2V_UNCONNECTED_2654,SV2V_UNCONNECTED_2655,SV2V_UNCONNECTED_2656,SV2V_UNCONNECTED_2657,
  SV2V_UNCONNECTED_2658,SV2V_UNCONNECTED_2659,SV2V_UNCONNECTED_2660,
  SV2V_UNCONNECTED_2661,SV2V_UNCONNECTED_2662,SV2V_UNCONNECTED_2663,
  SV2V_UNCONNECTED_2664,SV2V_UNCONNECTED_2665,SV2V_UNCONNECTED_2666,
  SV2V_UNCONNECTED_2667,SV2V_UNCONNECTED_2668,SV2V_UNCONNECTED_2669,
  SV2V_UNCONNECTED_2670,SV2V_UNCONNECTED_2671,SV2V_UNCONNECTED_2672,
  SV2V_UNCONNECTED_2673,SV2V_UNCONNECTED_2674,SV2V_UNCONNECTED_2675,
  SV2V_UNCONNECTED_2676,SV2V_UNCONNECTED_2677,SV2V_UNCONNECTED_2678,
  SV2V_UNCONNECTED_2679,SV2V_UNCONNECTED_2680,SV2V_UNCONNECTED_2681,
  SV2V_UNCONNECTED_2682,SV2V_UNCONNECTED_2683,SV2V_UNCONNECTED_2684,
  SV2V_UNCONNECTED_2685,SV2V_UNCONNECTED_2686,SV2V_UNCONNECTED_2687,
  SV2V_UNCONNECTED_2688,SV2V_UNCONNECTED_2689,SV2V_UNCONNECTED_2690,
  SV2V_UNCONNECTED_2691,SV2V_UNCONNECTED_2692,SV2V_UNCONNECTED_2693,
  SV2V_UNCONNECTED_2694,SV2V_UNCONNECTED_2695,SV2V_UNCONNECTED_2696,SV2V_UNCONNECTED_2697,
  SV2V_UNCONNECTED_2698,SV2V_UNCONNECTED_2699,SV2V_UNCONNECTED_2700,
  SV2V_UNCONNECTED_2701,SV2V_UNCONNECTED_2702,SV2V_UNCONNECTED_2703,
  SV2V_UNCONNECTED_2704,SV2V_UNCONNECTED_2705,SV2V_UNCONNECTED_2706,
  SV2V_UNCONNECTED_2707,SV2V_UNCONNECTED_2708,SV2V_UNCONNECTED_2709,
  SV2V_UNCONNECTED_2710,SV2V_UNCONNECTED_2711,SV2V_UNCONNECTED_2712,
  SV2V_UNCONNECTED_2713,SV2V_UNCONNECTED_2714,SV2V_UNCONNECTED_2715,
  SV2V_UNCONNECTED_2716,SV2V_UNCONNECTED_2717,SV2V_UNCONNECTED_2718,
  SV2V_UNCONNECTED_2719,SV2V_UNCONNECTED_2720,SV2V_UNCONNECTED_2721,
  SV2V_UNCONNECTED_2722,SV2V_UNCONNECTED_2723,SV2V_UNCONNECTED_2724,
  SV2V_UNCONNECTED_2725,SV2V_UNCONNECTED_2726,SV2V_UNCONNECTED_2727,
  SV2V_UNCONNECTED_2728,SV2V_UNCONNECTED_2729,SV2V_UNCONNECTED_2730,
  SV2V_UNCONNECTED_2731,SV2V_UNCONNECTED_2732,SV2V_UNCONNECTED_2733,
  SV2V_UNCONNECTED_2734,SV2V_UNCONNECTED_2735,SV2V_UNCONNECTED_2736,SV2V_UNCONNECTED_2737,
  SV2V_UNCONNECTED_2738,SV2V_UNCONNECTED_2739,SV2V_UNCONNECTED_2740,
  SV2V_UNCONNECTED_2741,SV2V_UNCONNECTED_2742,SV2V_UNCONNECTED_2743,
  SV2V_UNCONNECTED_2744,SV2V_UNCONNECTED_2745,SV2V_UNCONNECTED_2746,
  SV2V_UNCONNECTED_2747,SV2V_UNCONNECTED_2748,SV2V_UNCONNECTED_2749,
  SV2V_UNCONNECTED_2750,SV2V_UNCONNECTED_2751,SV2V_UNCONNECTED_2752,
  SV2V_UNCONNECTED_2753,SV2V_UNCONNECTED_2754,SV2V_UNCONNECTED_2755,
  SV2V_UNCONNECTED_2756,SV2V_UNCONNECTED_2757,SV2V_UNCONNECTED_2758,
  SV2V_UNCONNECTED_2759,SV2V_UNCONNECTED_2760,SV2V_UNCONNECTED_2761,
  SV2V_UNCONNECTED_2762,SV2V_UNCONNECTED_2763,SV2V_UNCONNECTED_2764,
  SV2V_UNCONNECTED_2765,SV2V_UNCONNECTED_2766,SV2V_UNCONNECTED_2767,
  SV2V_UNCONNECTED_2768,SV2V_UNCONNECTED_2769,SV2V_UNCONNECTED_2770,
  SV2V_UNCONNECTED_2771,SV2V_UNCONNECTED_2772,SV2V_UNCONNECTED_2773,
  SV2V_UNCONNECTED_2774,SV2V_UNCONNECTED_2775,SV2V_UNCONNECTED_2776,SV2V_UNCONNECTED_2777,
  SV2V_UNCONNECTED_2778,SV2V_UNCONNECTED_2779,SV2V_UNCONNECTED_2780,
  SV2V_UNCONNECTED_2781,SV2V_UNCONNECTED_2782,SV2V_UNCONNECTED_2783,
  SV2V_UNCONNECTED_2784,SV2V_UNCONNECTED_2785,SV2V_UNCONNECTED_2786,
  SV2V_UNCONNECTED_2787,SV2V_UNCONNECTED_2788,SV2V_UNCONNECTED_2789,
  SV2V_UNCONNECTED_2790,SV2V_UNCONNECTED_2791,SV2V_UNCONNECTED_2792,
  SV2V_UNCONNECTED_2793,SV2V_UNCONNECTED_2794,SV2V_UNCONNECTED_2795,
  SV2V_UNCONNECTED_2796,SV2V_UNCONNECTED_2797,SV2V_UNCONNECTED_2798,
  SV2V_UNCONNECTED_2799,SV2V_UNCONNECTED_2800,SV2V_UNCONNECTED_2801,
  SV2V_UNCONNECTED_2802,SV2V_UNCONNECTED_2803,SV2V_UNCONNECTED_2804,
  SV2V_UNCONNECTED_2805,SV2V_UNCONNECTED_2806,SV2V_UNCONNECTED_2807,
  SV2V_UNCONNECTED_2808,SV2V_UNCONNECTED_2809,SV2V_UNCONNECTED_2810,
  SV2V_UNCONNECTED_2811,SV2V_UNCONNECTED_2812,SV2V_UNCONNECTED_2813,
  SV2V_UNCONNECTED_2814,SV2V_UNCONNECTED_2815,SV2V_UNCONNECTED_2816,SV2V_UNCONNECTED_2817,
  SV2V_UNCONNECTED_2818,SV2V_UNCONNECTED_2819,SV2V_UNCONNECTED_2820,
  SV2V_UNCONNECTED_2821,SV2V_UNCONNECTED_2822,SV2V_UNCONNECTED_2823,
  SV2V_UNCONNECTED_2824,SV2V_UNCONNECTED_2825,SV2V_UNCONNECTED_2826,
  SV2V_UNCONNECTED_2827,SV2V_UNCONNECTED_2828,SV2V_UNCONNECTED_2829,
  SV2V_UNCONNECTED_2830,SV2V_UNCONNECTED_2831,SV2V_UNCONNECTED_2832,
  SV2V_UNCONNECTED_2833,SV2V_UNCONNECTED_2834,SV2V_UNCONNECTED_2835,
  SV2V_UNCONNECTED_2836,SV2V_UNCONNECTED_2837,SV2V_UNCONNECTED_2838,
  SV2V_UNCONNECTED_2839,SV2V_UNCONNECTED_2840,SV2V_UNCONNECTED_2841,
  SV2V_UNCONNECTED_2842,SV2V_UNCONNECTED_2843,SV2V_UNCONNECTED_2844,
  SV2V_UNCONNECTED_2845,SV2V_UNCONNECTED_2846,SV2V_UNCONNECTED_2847,
  SV2V_UNCONNECTED_2848,SV2V_UNCONNECTED_2849,SV2V_UNCONNECTED_2850,
  SV2V_UNCONNECTED_2851,SV2V_UNCONNECTED_2852,SV2V_UNCONNECTED_2853,
  SV2V_UNCONNECTED_2854,SV2V_UNCONNECTED_2855,SV2V_UNCONNECTED_2856,SV2V_UNCONNECTED_2857,
  SV2V_UNCONNECTED_2858,SV2V_UNCONNECTED_2859,SV2V_UNCONNECTED_2860,
  SV2V_UNCONNECTED_2861,SV2V_UNCONNECTED_2862,SV2V_UNCONNECTED_2863,
  SV2V_UNCONNECTED_2864,SV2V_UNCONNECTED_2865,SV2V_UNCONNECTED_2866,
  SV2V_UNCONNECTED_2867,SV2V_UNCONNECTED_2868,SV2V_UNCONNECTED_2869,
  SV2V_UNCONNECTED_2870,SV2V_UNCONNECTED_2871,SV2V_UNCONNECTED_2872,
  SV2V_UNCONNECTED_2873,SV2V_UNCONNECTED_2874,SV2V_UNCONNECTED_2875,
  SV2V_UNCONNECTED_2876,SV2V_UNCONNECTED_2877,SV2V_UNCONNECTED_2878,
  SV2V_UNCONNECTED_2879,SV2V_UNCONNECTED_2880,SV2V_UNCONNECTED_2881,
  SV2V_UNCONNECTED_2882,SV2V_UNCONNECTED_2883,SV2V_UNCONNECTED_2884,
  SV2V_UNCONNECTED_2885,SV2V_UNCONNECTED_2886,SV2V_UNCONNECTED_2887,
  SV2V_UNCONNECTED_2888,SV2V_UNCONNECTED_2889,SV2V_UNCONNECTED_2890,
  SV2V_UNCONNECTED_2891,SV2V_UNCONNECTED_2892,SV2V_UNCONNECTED_2893,
  SV2V_UNCONNECTED_2894,SV2V_UNCONNECTED_2895,SV2V_UNCONNECTED_2896,SV2V_UNCONNECTED_2897,
  SV2V_UNCONNECTED_2898,SV2V_UNCONNECTED_2899,SV2V_UNCONNECTED_2900,
  SV2V_UNCONNECTED_2901,SV2V_UNCONNECTED_2902,SV2V_UNCONNECTED_2903,
  SV2V_UNCONNECTED_2904,SV2V_UNCONNECTED_2905,SV2V_UNCONNECTED_2906,
  SV2V_UNCONNECTED_2907,SV2V_UNCONNECTED_2908,SV2V_UNCONNECTED_2909,
  SV2V_UNCONNECTED_2910,SV2V_UNCONNECTED_2911,SV2V_UNCONNECTED_2912,
  SV2V_UNCONNECTED_2913,SV2V_UNCONNECTED_2914,SV2V_UNCONNECTED_2915,
  SV2V_UNCONNECTED_2916,SV2V_UNCONNECTED_2917,SV2V_UNCONNECTED_2918,
  SV2V_UNCONNECTED_2919,SV2V_UNCONNECTED_2920,SV2V_UNCONNECTED_2921,
  SV2V_UNCONNECTED_2922,SV2V_UNCONNECTED_2923,SV2V_UNCONNECTED_2924,
  SV2V_UNCONNECTED_2925,SV2V_UNCONNECTED_2926,SV2V_UNCONNECTED_2927,
  SV2V_UNCONNECTED_2928,SV2V_UNCONNECTED_2929,SV2V_UNCONNECTED_2930,
  SV2V_UNCONNECTED_2931,SV2V_UNCONNECTED_2932,SV2V_UNCONNECTED_2933,
  SV2V_UNCONNECTED_2934,SV2V_UNCONNECTED_2935,SV2V_UNCONNECTED_2936,SV2V_UNCONNECTED_2937,
  SV2V_UNCONNECTED_2938,SV2V_UNCONNECTED_2939,SV2V_UNCONNECTED_2940,
  SV2V_UNCONNECTED_2941,SV2V_UNCONNECTED_2942,SV2V_UNCONNECTED_2943,
  SV2V_UNCONNECTED_2944,SV2V_UNCONNECTED_2945,SV2V_UNCONNECTED_2946,
  SV2V_UNCONNECTED_2947,SV2V_UNCONNECTED_2948,SV2V_UNCONNECTED_2949,
  SV2V_UNCONNECTED_2950,SV2V_UNCONNECTED_2951,SV2V_UNCONNECTED_2952,
  SV2V_UNCONNECTED_2953,SV2V_UNCONNECTED_2954,SV2V_UNCONNECTED_2955,
  SV2V_UNCONNECTED_2956,SV2V_UNCONNECTED_2957,SV2V_UNCONNECTED_2958,
  SV2V_UNCONNECTED_2959,SV2V_UNCONNECTED_2960,SV2V_UNCONNECTED_2961,
  SV2V_UNCONNECTED_2962,SV2V_UNCONNECTED_2963,SV2V_UNCONNECTED_2964,
  SV2V_UNCONNECTED_2965,SV2V_UNCONNECTED_2966,SV2V_UNCONNECTED_2967,
  SV2V_UNCONNECTED_2968,SV2V_UNCONNECTED_2969,SV2V_UNCONNECTED_2970,
  SV2V_UNCONNECTED_2971,SV2V_UNCONNECTED_2972,SV2V_UNCONNECTED_2973,
  SV2V_UNCONNECTED_2974,SV2V_UNCONNECTED_2975,SV2V_UNCONNECTED_2976,SV2V_UNCONNECTED_2977,
  SV2V_UNCONNECTED_2978,SV2V_UNCONNECTED_2979,SV2V_UNCONNECTED_2980,
  SV2V_UNCONNECTED_2981,SV2V_UNCONNECTED_2982,SV2V_UNCONNECTED_2983,
  SV2V_UNCONNECTED_2984,SV2V_UNCONNECTED_2985,SV2V_UNCONNECTED_2986,
  SV2V_UNCONNECTED_2987,SV2V_UNCONNECTED_2988,SV2V_UNCONNECTED_2989,
  SV2V_UNCONNECTED_2990,SV2V_UNCONNECTED_2991,SV2V_UNCONNECTED_2992,
  SV2V_UNCONNECTED_2993,SV2V_UNCONNECTED_2994,SV2V_UNCONNECTED_2995,
  SV2V_UNCONNECTED_2996,SV2V_UNCONNECTED_2997,SV2V_UNCONNECTED_2998,
  SV2V_UNCONNECTED_2999,SV2V_UNCONNECTED_3000,SV2V_UNCONNECTED_3001,
  SV2V_UNCONNECTED_3002,SV2V_UNCONNECTED_3003,SV2V_UNCONNECTED_3004,
  SV2V_UNCONNECTED_3005,SV2V_UNCONNECTED_3006,SV2V_UNCONNECTED_3007,
  SV2V_UNCONNECTED_3008,SV2V_UNCONNECTED_3009,SV2V_UNCONNECTED_3010,
  SV2V_UNCONNECTED_3011,SV2V_UNCONNECTED_3012,SV2V_UNCONNECTED_3013,
  SV2V_UNCONNECTED_3014,SV2V_UNCONNECTED_3015,SV2V_UNCONNECTED_3016,SV2V_UNCONNECTED_3017,
  SV2V_UNCONNECTED_3018,SV2V_UNCONNECTED_3019,SV2V_UNCONNECTED_3020,
  SV2V_UNCONNECTED_3021,SV2V_UNCONNECTED_3022,SV2V_UNCONNECTED_3023,
  SV2V_UNCONNECTED_3024,SV2V_UNCONNECTED_3025,SV2V_UNCONNECTED_3026,
  SV2V_UNCONNECTED_3027,SV2V_UNCONNECTED_3028,SV2V_UNCONNECTED_3029,
  SV2V_UNCONNECTED_3030,SV2V_UNCONNECTED_3031,SV2V_UNCONNECTED_3032,
  SV2V_UNCONNECTED_3033,SV2V_UNCONNECTED_3034,SV2V_UNCONNECTED_3035,
  SV2V_UNCONNECTED_3036,SV2V_UNCONNECTED_3037,SV2V_UNCONNECTED_3038,
  SV2V_UNCONNECTED_3039,SV2V_UNCONNECTED_3040,SV2V_UNCONNECTED_3041,
  SV2V_UNCONNECTED_3042,SV2V_UNCONNECTED_3043,SV2V_UNCONNECTED_3044,
  SV2V_UNCONNECTED_3045,SV2V_UNCONNECTED_3046,SV2V_UNCONNECTED_3047,
  SV2V_UNCONNECTED_3048,SV2V_UNCONNECTED_3049,SV2V_UNCONNECTED_3050,
  SV2V_UNCONNECTED_3051,SV2V_UNCONNECTED_3052,SV2V_UNCONNECTED_3053,
  SV2V_UNCONNECTED_3054,SV2V_UNCONNECTED_3055,SV2V_UNCONNECTED_3056,SV2V_UNCONNECTED_3057,
  SV2V_UNCONNECTED_3058,SV2V_UNCONNECTED_3059,SV2V_UNCONNECTED_3060,
  SV2V_UNCONNECTED_3061,SV2V_UNCONNECTED_3062,SV2V_UNCONNECTED_3063,
  SV2V_UNCONNECTED_3064,SV2V_UNCONNECTED_3065,SV2V_UNCONNECTED_3066,
  SV2V_UNCONNECTED_3067,SV2V_UNCONNECTED_3068,SV2V_UNCONNECTED_3069,
  SV2V_UNCONNECTED_3070,SV2V_UNCONNECTED_3071,SV2V_UNCONNECTED_3072,
  SV2V_UNCONNECTED_3073,SV2V_UNCONNECTED_3074,SV2V_UNCONNECTED_3075,
  SV2V_UNCONNECTED_3076,SV2V_UNCONNECTED_3077,SV2V_UNCONNECTED_3078,
  SV2V_UNCONNECTED_3079,SV2V_UNCONNECTED_3080,SV2V_UNCONNECTED_3081,
  SV2V_UNCONNECTED_3082,SV2V_UNCONNECTED_3083,SV2V_UNCONNECTED_3084,
  SV2V_UNCONNECTED_3085,SV2V_UNCONNECTED_3086,SV2V_UNCONNECTED_3087,
  SV2V_UNCONNECTED_3088,SV2V_UNCONNECTED_3089,SV2V_UNCONNECTED_3090,
  SV2V_UNCONNECTED_3091,SV2V_UNCONNECTED_3092,SV2V_UNCONNECTED_3093,
  SV2V_UNCONNECTED_3094,SV2V_UNCONNECTED_3095,SV2V_UNCONNECTED_3096,SV2V_UNCONNECTED_3097,
  SV2V_UNCONNECTED_3098,SV2V_UNCONNECTED_3099,SV2V_UNCONNECTED_3100,
  SV2V_UNCONNECTED_3101,SV2V_UNCONNECTED_3102,SV2V_UNCONNECTED_3103,
  SV2V_UNCONNECTED_3104,SV2V_UNCONNECTED_3105,SV2V_UNCONNECTED_3106,
  SV2V_UNCONNECTED_3107,SV2V_UNCONNECTED_3108,SV2V_UNCONNECTED_3109,
  SV2V_UNCONNECTED_3110,SV2V_UNCONNECTED_3111,SV2V_UNCONNECTED_3112,
  SV2V_UNCONNECTED_3113,SV2V_UNCONNECTED_3114,SV2V_UNCONNECTED_3115,
  SV2V_UNCONNECTED_3116,SV2V_UNCONNECTED_3117,SV2V_UNCONNECTED_3118,
  SV2V_UNCONNECTED_3119,SV2V_UNCONNECTED_3120,SV2V_UNCONNECTED_3121,
  SV2V_UNCONNECTED_3122,SV2V_UNCONNECTED_3123,SV2V_UNCONNECTED_3124,
  SV2V_UNCONNECTED_3125,SV2V_UNCONNECTED_3126,SV2V_UNCONNECTED_3127,
  SV2V_UNCONNECTED_3128,SV2V_UNCONNECTED_3129,SV2V_UNCONNECTED_3130,
  SV2V_UNCONNECTED_3131,SV2V_UNCONNECTED_3132,SV2V_UNCONNECTED_3133,
  SV2V_UNCONNECTED_3134,SV2V_UNCONNECTED_3135,SV2V_UNCONNECTED_3136,SV2V_UNCONNECTED_3137,
  SV2V_UNCONNECTED_3138,SV2V_UNCONNECTED_3139,SV2V_UNCONNECTED_3140,
  SV2V_UNCONNECTED_3141,SV2V_UNCONNECTED_3142,SV2V_UNCONNECTED_3143,
  SV2V_UNCONNECTED_3144,SV2V_UNCONNECTED_3145,SV2V_UNCONNECTED_3146,
  SV2V_UNCONNECTED_3147,SV2V_UNCONNECTED_3148,SV2V_UNCONNECTED_3149,
  SV2V_UNCONNECTED_3150,SV2V_UNCONNECTED_3151,SV2V_UNCONNECTED_3152,
  SV2V_UNCONNECTED_3153,SV2V_UNCONNECTED_3154,SV2V_UNCONNECTED_3155,
  SV2V_UNCONNECTED_3156,SV2V_UNCONNECTED_3157,SV2V_UNCONNECTED_3158,
  SV2V_UNCONNECTED_3159,SV2V_UNCONNECTED_3160,SV2V_UNCONNECTED_3161,
  SV2V_UNCONNECTED_3162,SV2V_UNCONNECTED_3163,SV2V_UNCONNECTED_3164,
  SV2V_UNCONNECTED_3165,SV2V_UNCONNECTED_3166,SV2V_UNCONNECTED_3167,
  SV2V_UNCONNECTED_3168,SV2V_UNCONNECTED_3169,SV2V_UNCONNECTED_3170,
  SV2V_UNCONNECTED_3171,SV2V_UNCONNECTED_3172,SV2V_UNCONNECTED_3173,
  SV2V_UNCONNECTED_3174,SV2V_UNCONNECTED_3175,SV2V_UNCONNECTED_3176,SV2V_UNCONNECTED_3177,
  SV2V_UNCONNECTED_3178,SV2V_UNCONNECTED_3179,SV2V_UNCONNECTED_3180,
  SV2V_UNCONNECTED_3181,SV2V_UNCONNECTED_3182,SV2V_UNCONNECTED_3183,
  SV2V_UNCONNECTED_3184,SV2V_UNCONNECTED_3185,SV2V_UNCONNECTED_3186,
  SV2V_UNCONNECTED_3187,SV2V_UNCONNECTED_3188,SV2V_UNCONNECTED_3189,
  SV2V_UNCONNECTED_3190,SV2V_UNCONNECTED_3191,SV2V_UNCONNECTED_3192,
  SV2V_UNCONNECTED_3193,SV2V_UNCONNECTED_3194,SV2V_UNCONNECTED_3195,
  SV2V_UNCONNECTED_3196,SV2V_UNCONNECTED_3197,SV2V_UNCONNECTED_3198,
  SV2V_UNCONNECTED_3199,SV2V_UNCONNECTED_3200,SV2V_UNCONNECTED_3201,
  SV2V_UNCONNECTED_3202,SV2V_UNCONNECTED_3203,SV2V_UNCONNECTED_3204,
  SV2V_UNCONNECTED_3205,SV2V_UNCONNECTED_3206,SV2V_UNCONNECTED_3207,
  SV2V_UNCONNECTED_3208,SV2V_UNCONNECTED_3209,SV2V_UNCONNECTED_3210,
  SV2V_UNCONNECTED_3211,SV2V_UNCONNECTED_3212,SV2V_UNCONNECTED_3213,
  SV2V_UNCONNECTED_3214,SV2V_UNCONNECTED_3215,SV2V_UNCONNECTED_3216,SV2V_UNCONNECTED_3217,
  SV2V_UNCONNECTED_3218,SV2V_UNCONNECTED_3219,SV2V_UNCONNECTED_3220,
  SV2V_UNCONNECTED_3221,SV2V_UNCONNECTED_3222,SV2V_UNCONNECTED_3223,
  SV2V_UNCONNECTED_3224,SV2V_UNCONNECTED_3225,SV2V_UNCONNECTED_3226,
  SV2V_UNCONNECTED_3227,SV2V_UNCONNECTED_3228,SV2V_UNCONNECTED_3229,
  SV2V_UNCONNECTED_3230,SV2V_UNCONNECTED_3231,SV2V_UNCONNECTED_3232,
  SV2V_UNCONNECTED_3233,SV2V_UNCONNECTED_3234,SV2V_UNCONNECTED_3235,
  SV2V_UNCONNECTED_3236,SV2V_UNCONNECTED_3237,SV2V_UNCONNECTED_3238,
  SV2V_UNCONNECTED_3239,SV2V_UNCONNECTED_3240,SV2V_UNCONNECTED_3241,
  SV2V_UNCONNECTED_3242,SV2V_UNCONNECTED_3243,SV2V_UNCONNECTED_3244,
  SV2V_UNCONNECTED_3245,SV2V_UNCONNECTED_3246,SV2V_UNCONNECTED_3247,
  SV2V_UNCONNECTED_3248,SV2V_UNCONNECTED_3249,SV2V_UNCONNECTED_3250,
  SV2V_UNCONNECTED_3251,SV2V_UNCONNECTED_3252,SV2V_UNCONNECTED_3253,
  SV2V_UNCONNECTED_3254,SV2V_UNCONNECTED_3255,SV2V_UNCONNECTED_3256,SV2V_UNCONNECTED_3257,
  SV2V_UNCONNECTED_3258,SV2V_UNCONNECTED_3259,SV2V_UNCONNECTED_3260,
  SV2V_UNCONNECTED_3261,SV2V_UNCONNECTED_3262,SV2V_UNCONNECTED_3263,
  SV2V_UNCONNECTED_3264,SV2V_UNCONNECTED_3265,SV2V_UNCONNECTED_3266,
  SV2V_UNCONNECTED_3267,SV2V_UNCONNECTED_3268,SV2V_UNCONNECTED_3269,
  SV2V_UNCONNECTED_3270,SV2V_UNCONNECTED_3271,SV2V_UNCONNECTED_3272,
  SV2V_UNCONNECTED_3273,SV2V_UNCONNECTED_3274,SV2V_UNCONNECTED_3275,
  SV2V_UNCONNECTED_3276,SV2V_UNCONNECTED_3277,SV2V_UNCONNECTED_3278,
  SV2V_UNCONNECTED_3279,SV2V_UNCONNECTED_3280,SV2V_UNCONNECTED_3281,
  SV2V_UNCONNECTED_3282,SV2V_UNCONNECTED_3283,SV2V_UNCONNECTED_3284,
  SV2V_UNCONNECTED_3285,SV2V_UNCONNECTED_3286,SV2V_UNCONNECTED_3287,
  SV2V_UNCONNECTED_3288,SV2V_UNCONNECTED_3289,SV2V_UNCONNECTED_3290,
  SV2V_UNCONNECTED_3291,SV2V_UNCONNECTED_3292,SV2V_UNCONNECTED_3293,
  SV2V_UNCONNECTED_3294,SV2V_UNCONNECTED_3295,SV2V_UNCONNECTED_3296,SV2V_UNCONNECTED_3297,
  SV2V_UNCONNECTED_3298,SV2V_UNCONNECTED_3299,SV2V_UNCONNECTED_3300,
  SV2V_UNCONNECTED_3301,SV2V_UNCONNECTED_3302,SV2V_UNCONNECTED_3303,
  SV2V_UNCONNECTED_3304,SV2V_UNCONNECTED_3305,SV2V_UNCONNECTED_3306,
  SV2V_UNCONNECTED_3307,SV2V_UNCONNECTED_3308,SV2V_UNCONNECTED_3309,
  SV2V_UNCONNECTED_3310,SV2V_UNCONNECTED_3311,SV2V_UNCONNECTED_3312,
  SV2V_UNCONNECTED_3313,SV2V_UNCONNECTED_3314,SV2V_UNCONNECTED_3315,
  SV2V_UNCONNECTED_3316,SV2V_UNCONNECTED_3317,SV2V_UNCONNECTED_3318,
  SV2V_UNCONNECTED_3319,SV2V_UNCONNECTED_3320,SV2V_UNCONNECTED_3321,
  SV2V_UNCONNECTED_3322,SV2V_UNCONNECTED_3323,SV2V_UNCONNECTED_3324,
  SV2V_UNCONNECTED_3325,SV2V_UNCONNECTED_3326,SV2V_UNCONNECTED_3327,
  SV2V_UNCONNECTED_3328,SV2V_UNCONNECTED_3329,SV2V_UNCONNECTED_3330,
  SV2V_UNCONNECTED_3331,SV2V_UNCONNECTED_3332,SV2V_UNCONNECTED_3333,
  SV2V_UNCONNECTED_3334,SV2V_UNCONNECTED_3335,SV2V_UNCONNECTED_3336,SV2V_UNCONNECTED_3337,
  SV2V_UNCONNECTED_3338,SV2V_UNCONNECTED_3339,SV2V_UNCONNECTED_3340,
  SV2V_UNCONNECTED_3341,SV2V_UNCONNECTED_3342,SV2V_UNCONNECTED_3343,
  SV2V_UNCONNECTED_3344,SV2V_UNCONNECTED_3345,SV2V_UNCONNECTED_3346,
  SV2V_UNCONNECTED_3347,SV2V_UNCONNECTED_3348,SV2V_UNCONNECTED_3349,
  SV2V_UNCONNECTED_3350,SV2V_UNCONNECTED_3351,SV2V_UNCONNECTED_3352,
  SV2V_UNCONNECTED_3353,SV2V_UNCONNECTED_3354,SV2V_UNCONNECTED_3355,
  SV2V_UNCONNECTED_3356,SV2V_UNCONNECTED_3357,SV2V_UNCONNECTED_3358,
  SV2V_UNCONNECTED_3359,SV2V_UNCONNECTED_3360,SV2V_UNCONNECTED_3361,
  SV2V_UNCONNECTED_3362,SV2V_UNCONNECTED_3363,SV2V_UNCONNECTED_3364,
  SV2V_UNCONNECTED_3365,SV2V_UNCONNECTED_3366,SV2V_UNCONNECTED_3367,
  SV2V_UNCONNECTED_3368,SV2V_UNCONNECTED_3369,SV2V_UNCONNECTED_3370,
  SV2V_UNCONNECTED_3371,SV2V_UNCONNECTED_3372,SV2V_UNCONNECTED_3373,
  SV2V_UNCONNECTED_3374,SV2V_UNCONNECTED_3375,SV2V_UNCONNECTED_3376,SV2V_UNCONNECTED_3377,
  SV2V_UNCONNECTED_3378,SV2V_UNCONNECTED_3379,SV2V_UNCONNECTED_3380,
  SV2V_UNCONNECTED_3381,SV2V_UNCONNECTED_3382,SV2V_UNCONNECTED_3383,
  SV2V_UNCONNECTED_3384,SV2V_UNCONNECTED_3385,SV2V_UNCONNECTED_3386,
  SV2V_UNCONNECTED_3387,SV2V_UNCONNECTED_3388,SV2V_UNCONNECTED_3389,
  SV2V_UNCONNECTED_3390,SV2V_UNCONNECTED_3391,SV2V_UNCONNECTED_3392,
  SV2V_UNCONNECTED_3393,SV2V_UNCONNECTED_3394,SV2V_UNCONNECTED_3395,
  SV2V_UNCONNECTED_3396,SV2V_UNCONNECTED_3397,SV2V_UNCONNECTED_3398,
  SV2V_UNCONNECTED_3399,SV2V_UNCONNECTED_3400,SV2V_UNCONNECTED_3401,
  SV2V_UNCONNECTED_3402,SV2V_UNCONNECTED_3403,SV2V_UNCONNECTED_3404,
  SV2V_UNCONNECTED_3405,SV2V_UNCONNECTED_3406,SV2V_UNCONNECTED_3407,
  SV2V_UNCONNECTED_3408,SV2V_UNCONNECTED_3409,SV2V_UNCONNECTED_3410,
  SV2V_UNCONNECTED_3411,SV2V_UNCONNECTED_3412,SV2V_UNCONNECTED_3413,
  SV2V_UNCONNECTED_3414,SV2V_UNCONNECTED_3415,SV2V_UNCONNECTED_3416,SV2V_UNCONNECTED_3417,
  SV2V_UNCONNECTED_3418,SV2V_UNCONNECTED_3419,SV2V_UNCONNECTED_3420,
  SV2V_UNCONNECTED_3421,SV2V_UNCONNECTED_3422,SV2V_UNCONNECTED_3423,
  SV2V_UNCONNECTED_3424,SV2V_UNCONNECTED_3425,SV2V_UNCONNECTED_3426,
  SV2V_UNCONNECTED_3427,SV2V_UNCONNECTED_3428,SV2V_UNCONNECTED_3429,
  SV2V_UNCONNECTED_3430,SV2V_UNCONNECTED_3431,SV2V_UNCONNECTED_3432,
  SV2V_UNCONNECTED_3433,SV2V_UNCONNECTED_3434,SV2V_UNCONNECTED_3435,
  SV2V_UNCONNECTED_3436,SV2V_UNCONNECTED_3437,SV2V_UNCONNECTED_3438,
  SV2V_UNCONNECTED_3439,SV2V_UNCONNECTED_3440,SV2V_UNCONNECTED_3441,
  SV2V_UNCONNECTED_3442,SV2V_UNCONNECTED_3443,SV2V_UNCONNECTED_3444,
  SV2V_UNCONNECTED_3445,SV2V_UNCONNECTED_3446,SV2V_UNCONNECTED_3447,
  SV2V_UNCONNECTED_3448,SV2V_UNCONNECTED_3449,SV2V_UNCONNECTED_3450,
  SV2V_UNCONNECTED_3451,SV2V_UNCONNECTED_3452,SV2V_UNCONNECTED_3453,
  SV2V_UNCONNECTED_3454,SV2V_UNCONNECTED_3455,SV2V_UNCONNECTED_3456,SV2V_UNCONNECTED_3457,
  SV2V_UNCONNECTED_3458,SV2V_UNCONNECTED_3459,SV2V_UNCONNECTED_3460,
  SV2V_UNCONNECTED_3461,SV2V_UNCONNECTED_3462,SV2V_UNCONNECTED_3463,
  SV2V_UNCONNECTED_3464,SV2V_UNCONNECTED_3465,SV2V_UNCONNECTED_3466,
  SV2V_UNCONNECTED_3467,SV2V_UNCONNECTED_3468,SV2V_UNCONNECTED_3469,
  SV2V_UNCONNECTED_3470,SV2V_UNCONNECTED_3471,SV2V_UNCONNECTED_3472,
  SV2V_UNCONNECTED_3473,SV2V_UNCONNECTED_3474,SV2V_UNCONNECTED_3475,
  SV2V_UNCONNECTED_3476,SV2V_UNCONNECTED_3477,SV2V_UNCONNECTED_3478,
  SV2V_UNCONNECTED_3479,SV2V_UNCONNECTED_3480,SV2V_UNCONNECTED_3481,
  SV2V_UNCONNECTED_3482,SV2V_UNCONNECTED_3483,SV2V_UNCONNECTED_3484,
  SV2V_UNCONNECTED_3485,SV2V_UNCONNECTED_3486,SV2V_UNCONNECTED_3487,
  SV2V_UNCONNECTED_3488,SV2V_UNCONNECTED_3489,SV2V_UNCONNECTED_3490,
  SV2V_UNCONNECTED_3491,SV2V_UNCONNECTED_3492,SV2V_UNCONNECTED_3493,
  SV2V_UNCONNECTED_3494,SV2V_UNCONNECTED_3495,SV2V_UNCONNECTED_3496,SV2V_UNCONNECTED_3497,
  SV2V_UNCONNECTED_3498,SV2V_UNCONNECTED_3499,SV2V_UNCONNECTED_3500,
  SV2V_UNCONNECTED_3501,SV2V_UNCONNECTED_3502,SV2V_UNCONNECTED_3503,
  SV2V_UNCONNECTED_3504,SV2V_UNCONNECTED_3505,SV2V_UNCONNECTED_3506,
  SV2V_UNCONNECTED_3507,SV2V_UNCONNECTED_3508,SV2V_UNCONNECTED_3509,
  SV2V_UNCONNECTED_3510,SV2V_UNCONNECTED_3511,SV2V_UNCONNECTED_3512,
  SV2V_UNCONNECTED_3513,SV2V_UNCONNECTED_3514,SV2V_UNCONNECTED_3515,
  SV2V_UNCONNECTED_3516,SV2V_UNCONNECTED_3517,SV2V_UNCONNECTED_3518,
  SV2V_UNCONNECTED_3519,SV2V_UNCONNECTED_3520,SV2V_UNCONNECTED_3521,
  SV2V_UNCONNECTED_3522,SV2V_UNCONNECTED_3523,SV2V_UNCONNECTED_3524,
  SV2V_UNCONNECTED_3525,SV2V_UNCONNECTED_3526,SV2V_UNCONNECTED_3527,
  SV2V_UNCONNECTED_3528,SV2V_UNCONNECTED_3529,SV2V_UNCONNECTED_3530,
  SV2V_UNCONNECTED_3531,SV2V_UNCONNECTED_3532,SV2V_UNCONNECTED_3533,
  SV2V_UNCONNECTED_3534,SV2V_UNCONNECTED_3535,SV2V_UNCONNECTED_3536,SV2V_UNCONNECTED_3537,
  SV2V_UNCONNECTED_3538,SV2V_UNCONNECTED_3539,SV2V_UNCONNECTED_3540,
  SV2V_UNCONNECTED_3541,SV2V_UNCONNECTED_3542,SV2V_UNCONNECTED_3543,
  SV2V_UNCONNECTED_3544,SV2V_UNCONNECTED_3545,SV2V_UNCONNECTED_3546,
  SV2V_UNCONNECTED_3547,SV2V_UNCONNECTED_3548,SV2V_UNCONNECTED_3549,
  SV2V_UNCONNECTED_3550,SV2V_UNCONNECTED_3551,SV2V_UNCONNECTED_3552,
  SV2V_UNCONNECTED_3553,SV2V_UNCONNECTED_3554,SV2V_UNCONNECTED_3555,
  SV2V_UNCONNECTED_3556,SV2V_UNCONNECTED_3557,SV2V_UNCONNECTED_3558,
  SV2V_UNCONNECTED_3559,SV2V_UNCONNECTED_3560,SV2V_UNCONNECTED_3561,
  SV2V_UNCONNECTED_3562,SV2V_UNCONNECTED_3563,SV2V_UNCONNECTED_3564,
  SV2V_UNCONNECTED_3565,SV2V_UNCONNECTED_3566,SV2V_UNCONNECTED_3567,
  SV2V_UNCONNECTED_3568,SV2V_UNCONNECTED_3569,SV2V_UNCONNECTED_3570,
  SV2V_UNCONNECTED_3571,SV2V_UNCONNECTED_3572,SV2V_UNCONNECTED_3573,
  SV2V_UNCONNECTED_3574,SV2V_UNCONNECTED_3575,SV2V_UNCONNECTED_3576,SV2V_UNCONNECTED_3577,
  SV2V_UNCONNECTED_3578,SV2V_UNCONNECTED_3579,SV2V_UNCONNECTED_3580,
  SV2V_UNCONNECTED_3581,SV2V_UNCONNECTED_3582,SV2V_UNCONNECTED_3583,
  SV2V_UNCONNECTED_3584,SV2V_UNCONNECTED_3585,SV2V_UNCONNECTED_3586,
  SV2V_UNCONNECTED_3587,SV2V_UNCONNECTED_3588,SV2V_UNCONNECTED_3589,
  SV2V_UNCONNECTED_3590,SV2V_UNCONNECTED_3591,SV2V_UNCONNECTED_3592,
  SV2V_UNCONNECTED_3593,SV2V_UNCONNECTED_3594,SV2V_UNCONNECTED_3595,
  SV2V_UNCONNECTED_3596,SV2V_UNCONNECTED_3597,SV2V_UNCONNECTED_3598,
  SV2V_UNCONNECTED_3599,SV2V_UNCONNECTED_3600,SV2V_UNCONNECTED_3601,
  SV2V_UNCONNECTED_3602,SV2V_UNCONNECTED_3603,SV2V_UNCONNECTED_3604,
  SV2V_UNCONNECTED_3605,SV2V_UNCONNECTED_3606,SV2V_UNCONNECTED_3607,
  SV2V_UNCONNECTED_3608,SV2V_UNCONNECTED_3609,SV2V_UNCONNECTED_3610,
  SV2V_UNCONNECTED_3611,SV2V_UNCONNECTED_3612,SV2V_UNCONNECTED_3613,
  SV2V_UNCONNECTED_3614,SV2V_UNCONNECTED_3615,SV2V_UNCONNECTED_3616,SV2V_UNCONNECTED_3617,
  SV2V_UNCONNECTED_3618,SV2V_UNCONNECTED_3619,SV2V_UNCONNECTED_3620,
  SV2V_UNCONNECTED_3621,SV2V_UNCONNECTED_3622,SV2V_UNCONNECTED_3623,
  SV2V_UNCONNECTED_3624,SV2V_UNCONNECTED_3625,SV2V_UNCONNECTED_3626,
  SV2V_UNCONNECTED_3627,SV2V_UNCONNECTED_3628,SV2V_UNCONNECTED_3629,
  SV2V_UNCONNECTED_3630,SV2V_UNCONNECTED_3631,SV2V_UNCONNECTED_3632,
  SV2V_UNCONNECTED_3633,SV2V_UNCONNECTED_3634,SV2V_UNCONNECTED_3635,
  SV2V_UNCONNECTED_3636,SV2V_UNCONNECTED_3637,SV2V_UNCONNECTED_3638,
  SV2V_UNCONNECTED_3639,SV2V_UNCONNECTED_3640,SV2V_UNCONNECTED_3641,
  SV2V_UNCONNECTED_3642,SV2V_UNCONNECTED_3643,SV2V_UNCONNECTED_3644,
  SV2V_UNCONNECTED_3645,SV2V_UNCONNECTED_3646,SV2V_UNCONNECTED_3647,
  SV2V_UNCONNECTED_3648,SV2V_UNCONNECTED_3649,SV2V_UNCONNECTED_3650,
  SV2V_UNCONNECTED_3651,SV2V_UNCONNECTED_3652,SV2V_UNCONNECTED_3653,
  SV2V_UNCONNECTED_3654,SV2V_UNCONNECTED_3655,SV2V_UNCONNECTED_3656,SV2V_UNCONNECTED_3657,
  SV2V_UNCONNECTED_3658,SV2V_UNCONNECTED_3659,SV2V_UNCONNECTED_3660,
  SV2V_UNCONNECTED_3661,SV2V_UNCONNECTED_3662,SV2V_UNCONNECTED_3663,
  SV2V_UNCONNECTED_3664,SV2V_UNCONNECTED_3665,SV2V_UNCONNECTED_3666,
  SV2V_UNCONNECTED_3667,SV2V_UNCONNECTED_3668,SV2V_UNCONNECTED_3669,
  SV2V_UNCONNECTED_3670,SV2V_UNCONNECTED_3671,SV2V_UNCONNECTED_3672,
  SV2V_UNCONNECTED_3673,SV2V_UNCONNECTED_3674,SV2V_UNCONNECTED_3675,
  SV2V_UNCONNECTED_3676,SV2V_UNCONNECTED_3677,SV2V_UNCONNECTED_3678,
  SV2V_UNCONNECTED_3679,SV2V_UNCONNECTED_3680,SV2V_UNCONNECTED_3681,
  SV2V_UNCONNECTED_3682,SV2V_UNCONNECTED_3683,SV2V_UNCONNECTED_3684,
  SV2V_UNCONNECTED_3685,SV2V_UNCONNECTED_3686,SV2V_UNCONNECTED_3687,
  SV2V_UNCONNECTED_3688,SV2V_UNCONNECTED_3689,SV2V_UNCONNECTED_3690,
  SV2V_UNCONNECTED_3691,SV2V_UNCONNECTED_3692,SV2V_UNCONNECTED_3693,
  SV2V_UNCONNECTED_3694,SV2V_UNCONNECTED_3695,SV2V_UNCONNECTED_3696,SV2V_UNCONNECTED_3697,
  SV2V_UNCONNECTED_3698,SV2V_UNCONNECTED_3699,SV2V_UNCONNECTED_3700,
  SV2V_UNCONNECTED_3701,SV2V_UNCONNECTED_3702,SV2V_UNCONNECTED_3703,
  SV2V_UNCONNECTED_3704,SV2V_UNCONNECTED_3705,SV2V_UNCONNECTED_3706,
  SV2V_UNCONNECTED_3707,SV2V_UNCONNECTED_3708,SV2V_UNCONNECTED_3709,
  SV2V_UNCONNECTED_3710,SV2V_UNCONNECTED_3711,SV2V_UNCONNECTED_3712,
  SV2V_UNCONNECTED_3713,SV2V_UNCONNECTED_3714,SV2V_UNCONNECTED_3715,
  SV2V_UNCONNECTED_3716,SV2V_UNCONNECTED_3717,SV2V_UNCONNECTED_3718,
  SV2V_UNCONNECTED_3719,SV2V_UNCONNECTED_3720,SV2V_UNCONNECTED_3721,
  SV2V_UNCONNECTED_3722,SV2V_UNCONNECTED_3723,SV2V_UNCONNECTED_3724,
  SV2V_UNCONNECTED_3725,SV2V_UNCONNECTED_3726,SV2V_UNCONNECTED_3727,
  SV2V_UNCONNECTED_3728,SV2V_UNCONNECTED_3729,SV2V_UNCONNECTED_3730,
  SV2V_UNCONNECTED_3731,SV2V_UNCONNECTED_3732,SV2V_UNCONNECTED_3733,
  SV2V_UNCONNECTED_3734,SV2V_UNCONNECTED_3735,SV2V_UNCONNECTED_3736,SV2V_UNCONNECTED_3737,
  SV2V_UNCONNECTED_3738,SV2V_UNCONNECTED_3739,SV2V_UNCONNECTED_3740,
  SV2V_UNCONNECTED_3741,SV2V_UNCONNECTED_3742,SV2V_UNCONNECTED_3743,
  SV2V_UNCONNECTED_3744,SV2V_UNCONNECTED_3745,SV2V_UNCONNECTED_3746,
  SV2V_UNCONNECTED_3747,SV2V_UNCONNECTED_3748,SV2V_UNCONNECTED_3749,
  SV2V_UNCONNECTED_3750,SV2V_UNCONNECTED_3751,SV2V_UNCONNECTED_3752,
  SV2V_UNCONNECTED_3753,SV2V_UNCONNECTED_3754,SV2V_UNCONNECTED_3755,
  SV2V_UNCONNECTED_3756,SV2V_UNCONNECTED_3757,SV2V_UNCONNECTED_3758,
  SV2V_UNCONNECTED_3759,SV2V_UNCONNECTED_3760,SV2V_UNCONNECTED_3761,
  SV2V_UNCONNECTED_3762,SV2V_UNCONNECTED_3763,SV2V_UNCONNECTED_3764,
  SV2V_UNCONNECTED_3765,SV2V_UNCONNECTED_3766,SV2V_UNCONNECTED_3767,
  SV2V_UNCONNECTED_3768,SV2V_UNCONNECTED_3769,SV2V_UNCONNECTED_3770,
  SV2V_UNCONNECTED_3771,SV2V_UNCONNECTED_3772,SV2V_UNCONNECTED_3773,
  SV2V_UNCONNECTED_3774,SV2V_UNCONNECTED_3775,SV2V_UNCONNECTED_3776,SV2V_UNCONNECTED_3777,
  SV2V_UNCONNECTED_3778,SV2V_UNCONNECTED_3779,SV2V_UNCONNECTED_3780,
  SV2V_UNCONNECTED_3781,SV2V_UNCONNECTED_3782,SV2V_UNCONNECTED_3783,
  SV2V_UNCONNECTED_3784,SV2V_UNCONNECTED_3785,SV2V_UNCONNECTED_3786,
  SV2V_UNCONNECTED_3787,SV2V_UNCONNECTED_3788,SV2V_UNCONNECTED_3789,
  SV2V_UNCONNECTED_3790,SV2V_UNCONNECTED_3791,SV2V_UNCONNECTED_3792,
  SV2V_UNCONNECTED_3793,SV2V_UNCONNECTED_3794,SV2V_UNCONNECTED_3795,
  SV2V_UNCONNECTED_3796,SV2V_UNCONNECTED_3797,SV2V_UNCONNECTED_3798,
  SV2V_UNCONNECTED_3799,SV2V_UNCONNECTED_3800,SV2V_UNCONNECTED_3801,
  SV2V_UNCONNECTED_3802,SV2V_UNCONNECTED_3803,SV2V_UNCONNECTED_3804,
  SV2V_UNCONNECTED_3805,SV2V_UNCONNECTED_3806,SV2V_UNCONNECTED_3807,
  SV2V_UNCONNECTED_3808,SV2V_UNCONNECTED_3809,SV2V_UNCONNECTED_3810,
  SV2V_UNCONNECTED_3811,SV2V_UNCONNECTED_3812,SV2V_UNCONNECTED_3813,
  SV2V_UNCONNECTED_3814,SV2V_UNCONNECTED_3815,SV2V_UNCONNECTED_3816,SV2V_UNCONNECTED_3817,
  SV2V_UNCONNECTED_3818,SV2V_UNCONNECTED_3819,SV2V_UNCONNECTED_3820,
  SV2V_UNCONNECTED_3821,SV2V_UNCONNECTED_3822,SV2V_UNCONNECTED_3823,
  SV2V_UNCONNECTED_3824,SV2V_UNCONNECTED_3825,SV2V_UNCONNECTED_3826,
  SV2V_UNCONNECTED_3827,SV2V_UNCONNECTED_3828,SV2V_UNCONNECTED_3829,
  SV2V_UNCONNECTED_3830,SV2V_UNCONNECTED_3831,SV2V_UNCONNECTED_3832,
  SV2V_UNCONNECTED_3833,SV2V_UNCONNECTED_3834,SV2V_UNCONNECTED_3835,
  SV2V_UNCONNECTED_3836,SV2V_UNCONNECTED_3837,SV2V_UNCONNECTED_3838,
  SV2V_UNCONNECTED_3839,SV2V_UNCONNECTED_3840,SV2V_UNCONNECTED_3841,
  SV2V_UNCONNECTED_3842,SV2V_UNCONNECTED_3843,SV2V_UNCONNECTED_3844,
  SV2V_UNCONNECTED_3845,SV2V_UNCONNECTED_3846,SV2V_UNCONNECTED_3847,
  SV2V_UNCONNECTED_3848,SV2V_UNCONNECTED_3849,SV2V_UNCONNECTED_3850,
  SV2V_UNCONNECTED_3851,SV2V_UNCONNECTED_3852,SV2V_UNCONNECTED_3853,
  SV2V_UNCONNECTED_3854,SV2V_UNCONNECTED_3855,SV2V_UNCONNECTED_3856,SV2V_UNCONNECTED_3857,
  SV2V_UNCONNECTED_3858,SV2V_UNCONNECTED_3859,SV2V_UNCONNECTED_3860,
  SV2V_UNCONNECTED_3861,SV2V_UNCONNECTED_3862,SV2V_UNCONNECTED_3863,
  SV2V_UNCONNECTED_3864,SV2V_UNCONNECTED_3865,SV2V_UNCONNECTED_3866,
  SV2V_UNCONNECTED_3867,SV2V_UNCONNECTED_3868,SV2V_UNCONNECTED_3869,
  SV2V_UNCONNECTED_3870,SV2V_UNCONNECTED_3871,SV2V_UNCONNECTED_3872,
  SV2V_UNCONNECTED_3873,SV2V_UNCONNECTED_3874,SV2V_UNCONNECTED_3875,
  SV2V_UNCONNECTED_3876,SV2V_UNCONNECTED_3877,SV2V_UNCONNECTED_3878,
  SV2V_UNCONNECTED_3879,SV2V_UNCONNECTED_3880,SV2V_UNCONNECTED_3881,
  SV2V_UNCONNECTED_3882,SV2V_UNCONNECTED_3883,SV2V_UNCONNECTED_3884,
  SV2V_UNCONNECTED_3885,SV2V_UNCONNECTED_3886,SV2V_UNCONNECTED_3887,
  SV2V_UNCONNECTED_3888,SV2V_UNCONNECTED_3889,SV2V_UNCONNECTED_3890,
  SV2V_UNCONNECTED_3891,SV2V_UNCONNECTED_3892,SV2V_UNCONNECTED_3893,
  SV2V_UNCONNECTED_3894,SV2V_UNCONNECTED_3895,SV2V_UNCONNECTED_3896,SV2V_UNCONNECTED_3897,
  SV2V_UNCONNECTED_3898,SV2V_UNCONNECTED_3899,SV2V_UNCONNECTED_3900,
  SV2V_UNCONNECTED_3901,SV2V_UNCONNECTED_3902,SV2V_UNCONNECTED_3903,
  SV2V_UNCONNECTED_3904,SV2V_UNCONNECTED_3905,SV2V_UNCONNECTED_3906,
  SV2V_UNCONNECTED_3907,SV2V_UNCONNECTED_3908,SV2V_UNCONNECTED_3909,
  SV2V_UNCONNECTED_3910,SV2V_UNCONNECTED_3911,SV2V_UNCONNECTED_3912,
  SV2V_UNCONNECTED_3913,SV2V_UNCONNECTED_3914,SV2V_UNCONNECTED_3915,
  SV2V_UNCONNECTED_3916,SV2V_UNCONNECTED_3917,SV2V_UNCONNECTED_3918,
  SV2V_UNCONNECTED_3919,SV2V_UNCONNECTED_3920,SV2V_UNCONNECTED_3921,
  SV2V_UNCONNECTED_3922,SV2V_UNCONNECTED_3923,SV2V_UNCONNECTED_3924,
  SV2V_UNCONNECTED_3925,SV2V_UNCONNECTED_3926,SV2V_UNCONNECTED_3927,
  SV2V_UNCONNECTED_3928,SV2V_UNCONNECTED_3929,SV2V_UNCONNECTED_3930,
  SV2V_UNCONNECTED_3931,SV2V_UNCONNECTED_3932,SV2V_UNCONNECTED_3933,
  SV2V_UNCONNECTED_3934,SV2V_UNCONNECTED_3935,SV2V_UNCONNECTED_3936,SV2V_UNCONNECTED_3937,
  SV2V_UNCONNECTED_3938,SV2V_UNCONNECTED_3939,SV2V_UNCONNECTED_3940,
  SV2V_UNCONNECTED_3941,SV2V_UNCONNECTED_3942,SV2V_UNCONNECTED_3943,
  SV2V_UNCONNECTED_3944,SV2V_UNCONNECTED_3945,SV2V_UNCONNECTED_3946,
  SV2V_UNCONNECTED_3947,SV2V_UNCONNECTED_3948,SV2V_UNCONNECTED_3949,
  SV2V_UNCONNECTED_3950,SV2V_UNCONNECTED_3951,SV2V_UNCONNECTED_3952,
  SV2V_UNCONNECTED_3953,SV2V_UNCONNECTED_3954,SV2V_UNCONNECTED_3955,
  SV2V_UNCONNECTED_3956,SV2V_UNCONNECTED_3957,SV2V_UNCONNECTED_3958,
  SV2V_UNCONNECTED_3959,SV2V_UNCONNECTED_3960,SV2V_UNCONNECTED_3961,
  SV2V_UNCONNECTED_3962,SV2V_UNCONNECTED_3963,SV2V_UNCONNECTED_3964,
  SV2V_UNCONNECTED_3965,SV2V_UNCONNECTED_3966,SV2V_UNCONNECTED_3967,
  SV2V_UNCONNECTED_3968,SV2V_UNCONNECTED_3969,SV2V_UNCONNECTED_3970,
  SV2V_UNCONNECTED_3971,SV2V_UNCONNECTED_3972,SV2V_UNCONNECTED_3973,
  SV2V_UNCONNECTED_3974,SV2V_UNCONNECTED_3975,SV2V_UNCONNECTED_3976,SV2V_UNCONNECTED_3977,
  SV2V_UNCONNECTED_3978,SV2V_UNCONNECTED_3979,SV2V_UNCONNECTED_3980,
  SV2V_UNCONNECTED_3981,SV2V_UNCONNECTED_3982,SV2V_UNCONNECTED_3983,
  SV2V_UNCONNECTED_3984,SV2V_UNCONNECTED_3985,SV2V_UNCONNECTED_3986,
  SV2V_UNCONNECTED_3987,SV2V_UNCONNECTED_3988,SV2V_UNCONNECTED_3989,
  SV2V_UNCONNECTED_3990,SV2V_UNCONNECTED_3991,SV2V_UNCONNECTED_3992,
  SV2V_UNCONNECTED_3993,SV2V_UNCONNECTED_3994,SV2V_UNCONNECTED_3995,
  SV2V_UNCONNECTED_3996,SV2V_UNCONNECTED_3997,SV2V_UNCONNECTED_3998,
  SV2V_UNCONNECTED_3999,SV2V_UNCONNECTED_4000,SV2V_UNCONNECTED_4001,
  SV2V_UNCONNECTED_4002,SV2V_UNCONNECTED_4003,SV2V_UNCONNECTED_4004,
  SV2V_UNCONNECTED_4005,SV2V_UNCONNECTED_4006,SV2V_UNCONNECTED_4007,
  SV2V_UNCONNECTED_4008,SV2V_UNCONNECTED_4009,SV2V_UNCONNECTED_4010,
  SV2V_UNCONNECTED_4011,SV2V_UNCONNECTED_4012,SV2V_UNCONNECTED_4013,
  SV2V_UNCONNECTED_4014,SV2V_UNCONNECTED_4015,SV2V_UNCONNECTED_4016,SV2V_UNCONNECTED_4017,
  SV2V_UNCONNECTED_4018,SV2V_UNCONNECTED_4019,SV2V_UNCONNECTED_4020,
  SV2V_UNCONNECTED_4021,SV2V_UNCONNECTED_4022,SV2V_UNCONNECTED_4023,
  SV2V_UNCONNECTED_4024,SV2V_UNCONNECTED_4025,SV2V_UNCONNECTED_4026,
  SV2V_UNCONNECTED_4027,SV2V_UNCONNECTED_4028,SV2V_UNCONNECTED_4029,
  SV2V_UNCONNECTED_4030,SV2V_UNCONNECTED_4031,SV2V_UNCONNECTED_4032,
  SV2V_UNCONNECTED_4033,SV2V_UNCONNECTED_4034,SV2V_UNCONNECTED_4035,
  SV2V_UNCONNECTED_4036,SV2V_UNCONNECTED_4037,SV2V_UNCONNECTED_4038,
  SV2V_UNCONNECTED_4039,SV2V_UNCONNECTED_4040,SV2V_UNCONNECTED_4041,
  SV2V_UNCONNECTED_4042,SV2V_UNCONNECTED_4043,SV2V_UNCONNECTED_4044,
  SV2V_UNCONNECTED_4045,SV2V_UNCONNECTED_4046,SV2V_UNCONNECTED_4047,
  SV2V_UNCONNECTED_4048,SV2V_UNCONNECTED_4049,SV2V_UNCONNECTED_4050,
  SV2V_UNCONNECTED_4051,SV2V_UNCONNECTED_4052,SV2V_UNCONNECTED_4053,
  SV2V_UNCONNECTED_4054,SV2V_UNCONNECTED_4055,SV2V_UNCONNECTED_4056,SV2V_UNCONNECTED_4057,
  SV2V_UNCONNECTED_4058,SV2V_UNCONNECTED_4059,SV2V_UNCONNECTED_4060,
  SV2V_UNCONNECTED_4061,SV2V_UNCONNECTED_4062,SV2V_UNCONNECTED_4063,
  SV2V_UNCONNECTED_4064,SV2V_UNCONNECTED_4065,SV2V_UNCONNECTED_4066,
  SV2V_UNCONNECTED_4067,SV2V_UNCONNECTED_4068,SV2V_UNCONNECTED_4069,
  SV2V_UNCONNECTED_4070,SV2V_UNCONNECTED_4071,SV2V_UNCONNECTED_4072,
  SV2V_UNCONNECTED_4073,SV2V_UNCONNECTED_4074,SV2V_UNCONNECTED_4075,
  SV2V_UNCONNECTED_4076,SV2V_UNCONNECTED_4077,SV2V_UNCONNECTED_4078,
  SV2V_UNCONNECTED_4079,SV2V_UNCONNECTED_4080,SV2V_UNCONNECTED_4081,
  SV2V_UNCONNECTED_4082,SV2V_UNCONNECTED_4083,SV2V_UNCONNECTED_4084,
  SV2V_UNCONNECTED_4085,SV2V_UNCONNECTED_4086,SV2V_UNCONNECTED_4087,
  SV2V_UNCONNECTED_4088,SV2V_UNCONNECTED_4089,SV2V_UNCONNECTED_4090,
  SV2V_UNCONNECTED_4091,SV2V_UNCONNECTED_4092,SV2V_UNCONNECTED_4093,
  SV2V_UNCONNECTED_4094,SV2V_UNCONNECTED_4095,SV2V_UNCONNECTED_4096,SV2V_UNCONNECTED_4097,
  SV2V_UNCONNECTED_4098,SV2V_UNCONNECTED_4099,SV2V_UNCONNECTED_4100,
  SV2V_UNCONNECTED_4101,SV2V_UNCONNECTED_4102,SV2V_UNCONNECTED_4103,
  SV2V_UNCONNECTED_4104,SV2V_UNCONNECTED_4105,SV2V_UNCONNECTED_4106,
  SV2V_UNCONNECTED_4107,SV2V_UNCONNECTED_4108,SV2V_UNCONNECTED_4109,
  SV2V_UNCONNECTED_4110,SV2V_UNCONNECTED_4111,SV2V_UNCONNECTED_4112,
  SV2V_UNCONNECTED_4113,SV2V_UNCONNECTED_4114,SV2V_UNCONNECTED_4115,
  SV2V_UNCONNECTED_4116,SV2V_UNCONNECTED_4117,SV2V_UNCONNECTED_4118,
  SV2V_UNCONNECTED_4119,SV2V_UNCONNECTED_4120,SV2V_UNCONNECTED_4121,
  SV2V_UNCONNECTED_4122,SV2V_UNCONNECTED_4123,SV2V_UNCONNECTED_4124,
  SV2V_UNCONNECTED_4125,SV2V_UNCONNECTED_4126,SV2V_UNCONNECTED_4127,
  SV2V_UNCONNECTED_4128,SV2V_UNCONNECTED_4129,SV2V_UNCONNECTED_4130,
  SV2V_UNCONNECTED_4131,SV2V_UNCONNECTED_4132,SV2V_UNCONNECTED_4133,
  SV2V_UNCONNECTED_4134,SV2V_UNCONNECTED_4135,SV2V_UNCONNECTED_4136,SV2V_UNCONNECTED_4137,
  SV2V_UNCONNECTED_4138,SV2V_UNCONNECTED_4139,SV2V_UNCONNECTED_4140,
  SV2V_UNCONNECTED_4141,SV2V_UNCONNECTED_4142,SV2V_UNCONNECTED_4143,
  SV2V_UNCONNECTED_4144,SV2V_UNCONNECTED_4145,SV2V_UNCONNECTED_4146,
  SV2V_UNCONNECTED_4147,SV2V_UNCONNECTED_4148,SV2V_UNCONNECTED_4149,
  SV2V_UNCONNECTED_4150,SV2V_UNCONNECTED_4151,SV2V_UNCONNECTED_4152,
  SV2V_UNCONNECTED_4153,SV2V_UNCONNECTED_4154,SV2V_UNCONNECTED_4155,
  SV2V_UNCONNECTED_4156,SV2V_UNCONNECTED_4157,SV2V_UNCONNECTED_4158,
  SV2V_UNCONNECTED_4159,SV2V_UNCONNECTED_4160,SV2V_UNCONNECTED_4161,
  SV2V_UNCONNECTED_4162,SV2V_UNCONNECTED_4163,SV2V_UNCONNECTED_4164,
  SV2V_UNCONNECTED_4165,SV2V_UNCONNECTED_4166,SV2V_UNCONNECTED_4167,
  SV2V_UNCONNECTED_4168,SV2V_UNCONNECTED_4169,SV2V_UNCONNECTED_4170,
  SV2V_UNCONNECTED_4171,SV2V_UNCONNECTED_4172,SV2V_UNCONNECTED_4173,
  SV2V_UNCONNECTED_4174,SV2V_UNCONNECTED_4175,SV2V_UNCONNECTED_4176,SV2V_UNCONNECTED_4177,
  SV2V_UNCONNECTED_4178,SV2V_UNCONNECTED_4179,SV2V_UNCONNECTED_4180,
  SV2V_UNCONNECTED_4181,SV2V_UNCONNECTED_4182,SV2V_UNCONNECTED_4183,
  SV2V_UNCONNECTED_4184,SV2V_UNCONNECTED_4185,SV2V_UNCONNECTED_4186,
  SV2V_UNCONNECTED_4187,SV2V_UNCONNECTED_4188,SV2V_UNCONNECTED_4189,
  SV2V_UNCONNECTED_4190,SV2V_UNCONNECTED_4191,SV2V_UNCONNECTED_4192,
  SV2V_UNCONNECTED_4193,SV2V_UNCONNECTED_4194,SV2V_UNCONNECTED_4195,
  SV2V_UNCONNECTED_4196,SV2V_UNCONNECTED_4197,SV2V_UNCONNECTED_4198,
  SV2V_UNCONNECTED_4199,SV2V_UNCONNECTED_4200,SV2V_UNCONNECTED_4201,
  SV2V_UNCONNECTED_4202,SV2V_UNCONNECTED_4203,SV2V_UNCONNECTED_4204,
  SV2V_UNCONNECTED_4205,SV2V_UNCONNECTED_4206,SV2V_UNCONNECTED_4207,
  SV2V_UNCONNECTED_4208,SV2V_UNCONNECTED_4209,SV2V_UNCONNECTED_4210,
  SV2V_UNCONNECTED_4211,SV2V_UNCONNECTED_4212,SV2V_UNCONNECTED_4213,
  SV2V_UNCONNECTED_4214,SV2V_UNCONNECTED_4215,SV2V_UNCONNECTED_4216,SV2V_UNCONNECTED_4217,
  SV2V_UNCONNECTED_4218,SV2V_UNCONNECTED_4219,SV2V_UNCONNECTED_4220,
  SV2V_UNCONNECTED_4221,SV2V_UNCONNECTED_4222,SV2V_UNCONNECTED_4223,
  SV2V_UNCONNECTED_4224,SV2V_UNCONNECTED_4225,SV2V_UNCONNECTED_4226,
  SV2V_UNCONNECTED_4227,SV2V_UNCONNECTED_4228,SV2V_UNCONNECTED_4229,
  SV2V_UNCONNECTED_4230,SV2V_UNCONNECTED_4231,SV2V_UNCONNECTED_4232,
  SV2V_UNCONNECTED_4233,SV2V_UNCONNECTED_4234,SV2V_UNCONNECTED_4235,
  SV2V_UNCONNECTED_4236,SV2V_UNCONNECTED_4237,SV2V_UNCONNECTED_4238,
  SV2V_UNCONNECTED_4239,SV2V_UNCONNECTED_4240,SV2V_UNCONNECTED_4241,
  SV2V_UNCONNECTED_4242,SV2V_UNCONNECTED_4243,SV2V_UNCONNECTED_4244,
  SV2V_UNCONNECTED_4245,SV2V_UNCONNECTED_4246,SV2V_UNCONNECTED_4247,
  SV2V_UNCONNECTED_4248,SV2V_UNCONNECTED_4249,SV2V_UNCONNECTED_4250,
  SV2V_UNCONNECTED_4251,SV2V_UNCONNECTED_4252,SV2V_UNCONNECTED_4253,
  SV2V_UNCONNECTED_4254,SV2V_UNCONNECTED_4255,SV2V_UNCONNECTED_4256,SV2V_UNCONNECTED_4257,
  SV2V_UNCONNECTED_4258,SV2V_UNCONNECTED_4259,SV2V_UNCONNECTED_4260,
  SV2V_UNCONNECTED_4261,SV2V_UNCONNECTED_4262,SV2V_UNCONNECTED_4263,
  SV2V_UNCONNECTED_4264,SV2V_UNCONNECTED_4265,SV2V_UNCONNECTED_4266,
  SV2V_UNCONNECTED_4267,SV2V_UNCONNECTED_4268,SV2V_UNCONNECTED_4269,
  SV2V_UNCONNECTED_4270,SV2V_UNCONNECTED_4271,SV2V_UNCONNECTED_4272,
  SV2V_UNCONNECTED_4273,SV2V_UNCONNECTED_4274,SV2V_UNCONNECTED_4275,
  SV2V_UNCONNECTED_4276,SV2V_UNCONNECTED_4277,SV2V_UNCONNECTED_4278,
  SV2V_UNCONNECTED_4279,SV2V_UNCONNECTED_4280,SV2V_UNCONNECTED_4281,
  SV2V_UNCONNECTED_4282,SV2V_UNCONNECTED_4283,SV2V_UNCONNECTED_4284,
  SV2V_UNCONNECTED_4285,SV2V_UNCONNECTED_4286,SV2V_UNCONNECTED_4287,
  SV2V_UNCONNECTED_4288,SV2V_UNCONNECTED_4289,SV2V_UNCONNECTED_4290,
  SV2V_UNCONNECTED_4291,SV2V_UNCONNECTED_4292,SV2V_UNCONNECTED_4293,
  SV2V_UNCONNECTED_4294,SV2V_UNCONNECTED_4295,SV2V_UNCONNECTED_4296,SV2V_UNCONNECTED_4297,
  SV2V_UNCONNECTED_4298,SV2V_UNCONNECTED_4299,SV2V_UNCONNECTED_4300,
  SV2V_UNCONNECTED_4301,SV2V_UNCONNECTED_4302,SV2V_UNCONNECTED_4303,
  SV2V_UNCONNECTED_4304,SV2V_UNCONNECTED_4305,SV2V_UNCONNECTED_4306,
  SV2V_UNCONNECTED_4307,SV2V_UNCONNECTED_4308,SV2V_UNCONNECTED_4309,
  SV2V_UNCONNECTED_4310,SV2V_UNCONNECTED_4311,SV2V_UNCONNECTED_4312,
  SV2V_UNCONNECTED_4313,SV2V_UNCONNECTED_4314,SV2V_UNCONNECTED_4315,
  SV2V_UNCONNECTED_4316,SV2V_UNCONNECTED_4317,SV2V_UNCONNECTED_4318,
  SV2V_UNCONNECTED_4319,SV2V_UNCONNECTED_4320,SV2V_UNCONNECTED_4321,
  SV2V_UNCONNECTED_4322,SV2V_UNCONNECTED_4323,SV2V_UNCONNECTED_4324,
  SV2V_UNCONNECTED_4325,SV2V_UNCONNECTED_4326,SV2V_UNCONNECTED_4327,
  SV2V_UNCONNECTED_4328,SV2V_UNCONNECTED_4329,SV2V_UNCONNECTED_4330,
  SV2V_UNCONNECTED_4331,SV2V_UNCONNECTED_4332,SV2V_UNCONNECTED_4333,
  SV2V_UNCONNECTED_4334,SV2V_UNCONNECTED_4335,SV2V_UNCONNECTED_4336,SV2V_UNCONNECTED_4337,
  SV2V_UNCONNECTED_4338,SV2V_UNCONNECTED_4339,SV2V_UNCONNECTED_4340,
  SV2V_UNCONNECTED_4341,SV2V_UNCONNECTED_4342,SV2V_UNCONNECTED_4343,
  SV2V_UNCONNECTED_4344,SV2V_UNCONNECTED_4345,SV2V_UNCONNECTED_4346,
  SV2V_UNCONNECTED_4347,SV2V_UNCONNECTED_4348,SV2V_UNCONNECTED_4349,
  SV2V_UNCONNECTED_4350,SV2V_UNCONNECTED_4351,SV2V_UNCONNECTED_4352,
  SV2V_UNCONNECTED_4353,SV2V_UNCONNECTED_4354,SV2V_UNCONNECTED_4355,
  SV2V_UNCONNECTED_4356,SV2V_UNCONNECTED_4357,SV2V_UNCONNECTED_4358,
  SV2V_UNCONNECTED_4359,SV2V_UNCONNECTED_4360,SV2V_UNCONNECTED_4361,
  SV2V_UNCONNECTED_4362,SV2V_UNCONNECTED_4363,SV2V_UNCONNECTED_4364,
  SV2V_UNCONNECTED_4365,SV2V_UNCONNECTED_4366,SV2V_UNCONNECTED_4367,
  SV2V_UNCONNECTED_4368,SV2V_UNCONNECTED_4369,SV2V_UNCONNECTED_4370,
  SV2V_UNCONNECTED_4371,SV2V_UNCONNECTED_4372,SV2V_UNCONNECTED_4373,
  SV2V_UNCONNECTED_4374,SV2V_UNCONNECTED_4375,SV2V_UNCONNECTED_4376,SV2V_UNCONNECTED_4377,
  SV2V_UNCONNECTED_4378,SV2V_UNCONNECTED_4379,SV2V_UNCONNECTED_4380,
  SV2V_UNCONNECTED_4381,SV2V_UNCONNECTED_4382,SV2V_UNCONNECTED_4383,
  SV2V_UNCONNECTED_4384,SV2V_UNCONNECTED_4385,SV2V_UNCONNECTED_4386,
  SV2V_UNCONNECTED_4387,SV2V_UNCONNECTED_4388,SV2V_UNCONNECTED_4389,
  SV2V_UNCONNECTED_4390,SV2V_UNCONNECTED_4391,SV2V_UNCONNECTED_4392,
  SV2V_UNCONNECTED_4393,SV2V_UNCONNECTED_4394,SV2V_UNCONNECTED_4395,
  SV2V_UNCONNECTED_4396,SV2V_UNCONNECTED_4397,SV2V_UNCONNECTED_4398,
  SV2V_UNCONNECTED_4399,SV2V_UNCONNECTED_4400,SV2V_UNCONNECTED_4401,
  SV2V_UNCONNECTED_4402,SV2V_UNCONNECTED_4403,SV2V_UNCONNECTED_4404,
  SV2V_UNCONNECTED_4405,SV2V_UNCONNECTED_4406,SV2V_UNCONNECTED_4407,
  SV2V_UNCONNECTED_4408,SV2V_UNCONNECTED_4409,SV2V_UNCONNECTED_4410,
  SV2V_UNCONNECTED_4411,SV2V_UNCONNECTED_4412,SV2V_UNCONNECTED_4413,
  SV2V_UNCONNECTED_4414,SV2V_UNCONNECTED_4415,SV2V_UNCONNECTED_4416,SV2V_UNCONNECTED_4417,
  SV2V_UNCONNECTED_4418,SV2V_UNCONNECTED_4419,SV2V_UNCONNECTED_4420,
  SV2V_UNCONNECTED_4421,SV2V_UNCONNECTED_4422,SV2V_UNCONNECTED_4423,
  SV2V_UNCONNECTED_4424,SV2V_UNCONNECTED_4425,SV2V_UNCONNECTED_4426,
  SV2V_UNCONNECTED_4427,SV2V_UNCONNECTED_4428,SV2V_UNCONNECTED_4429,
  SV2V_UNCONNECTED_4430,SV2V_UNCONNECTED_4431,SV2V_UNCONNECTED_4432,
  SV2V_UNCONNECTED_4433,SV2V_UNCONNECTED_4434,SV2V_UNCONNECTED_4435,
  SV2V_UNCONNECTED_4436,SV2V_UNCONNECTED_4437,SV2V_UNCONNECTED_4438,
  SV2V_UNCONNECTED_4439,SV2V_UNCONNECTED_4440,SV2V_UNCONNECTED_4441,
  SV2V_UNCONNECTED_4442,SV2V_UNCONNECTED_4443,SV2V_UNCONNECTED_4444,
  SV2V_UNCONNECTED_4445,SV2V_UNCONNECTED_4446,SV2V_UNCONNECTED_4447,
  SV2V_UNCONNECTED_4448,SV2V_UNCONNECTED_4449,SV2V_UNCONNECTED_4450,
  SV2V_UNCONNECTED_4451,SV2V_UNCONNECTED_4452,SV2V_UNCONNECTED_4453,
  SV2V_UNCONNECTED_4454,SV2V_UNCONNECTED_4455,SV2V_UNCONNECTED_4456,SV2V_UNCONNECTED_4457,
  SV2V_UNCONNECTED_4458,SV2V_UNCONNECTED_4459,SV2V_UNCONNECTED_4460,
  SV2V_UNCONNECTED_4461,SV2V_UNCONNECTED_4462,SV2V_UNCONNECTED_4463,
  SV2V_UNCONNECTED_4464,SV2V_UNCONNECTED_4465,SV2V_UNCONNECTED_4466,
  SV2V_UNCONNECTED_4467,SV2V_UNCONNECTED_4468,SV2V_UNCONNECTED_4469,
  SV2V_UNCONNECTED_4470,SV2V_UNCONNECTED_4471,SV2V_UNCONNECTED_4472,
  SV2V_UNCONNECTED_4473,SV2V_UNCONNECTED_4474,SV2V_UNCONNECTED_4475,
  SV2V_UNCONNECTED_4476,SV2V_UNCONNECTED_4477,SV2V_UNCONNECTED_4478,
  SV2V_UNCONNECTED_4479,SV2V_UNCONNECTED_4480,SV2V_UNCONNECTED_4481,
  SV2V_UNCONNECTED_4482,SV2V_UNCONNECTED_4483,SV2V_UNCONNECTED_4484,
  SV2V_UNCONNECTED_4485,SV2V_UNCONNECTED_4486,SV2V_UNCONNECTED_4487,
  SV2V_UNCONNECTED_4488,SV2V_UNCONNECTED_4489,SV2V_UNCONNECTED_4490,
  SV2V_UNCONNECTED_4491,SV2V_UNCONNECTED_4492,SV2V_UNCONNECTED_4493,
  SV2V_UNCONNECTED_4494,SV2V_UNCONNECTED_4495,SV2V_UNCONNECTED_4496,SV2V_UNCONNECTED_4497,
  SV2V_UNCONNECTED_4498,SV2V_UNCONNECTED_4499,SV2V_UNCONNECTED_4500,
  SV2V_UNCONNECTED_4501,SV2V_UNCONNECTED_4502,SV2V_UNCONNECTED_4503,
  SV2V_UNCONNECTED_4504,SV2V_UNCONNECTED_4505,SV2V_UNCONNECTED_4506,
  SV2V_UNCONNECTED_4507,SV2V_UNCONNECTED_4508,SV2V_UNCONNECTED_4509,
  SV2V_UNCONNECTED_4510,SV2V_UNCONNECTED_4511,SV2V_UNCONNECTED_4512,
  SV2V_UNCONNECTED_4513,SV2V_UNCONNECTED_4514,SV2V_UNCONNECTED_4515,
  SV2V_UNCONNECTED_4516,SV2V_UNCONNECTED_4517,SV2V_UNCONNECTED_4518,
  SV2V_UNCONNECTED_4519,SV2V_UNCONNECTED_4520,SV2V_UNCONNECTED_4521,
  SV2V_UNCONNECTED_4522,SV2V_UNCONNECTED_4523,SV2V_UNCONNECTED_4524,
  SV2V_UNCONNECTED_4525,SV2V_UNCONNECTED_4526,SV2V_UNCONNECTED_4527,
  SV2V_UNCONNECTED_4528,SV2V_UNCONNECTED_4529,SV2V_UNCONNECTED_4530,
  SV2V_UNCONNECTED_4531,SV2V_UNCONNECTED_4532,SV2V_UNCONNECTED_4533,
  SV2V_UNCONNECTED_4534,SV2V_UNCONNECTED_4535,SV2V_UNCONNECTED_4536,SV2V_UNCONNECTED_4537,
  SV2V_UNCONNECTED_4538,SV2V_UNCONNECTED_4539,SV2V_UNCONNECTED_4540,
  SV2V_UNCONNECTED_4541,SV2V_UNCONNECTED_4542,SV2V_UNCONNECTED_4543,
  SV2V_UNCONNECTED_4544,SV2V_UNCONNECTED_4545,SV2V_UNCONNECTED_4546,
  SV2V_UNCONNECTED_4547,SV2V_UNCONNECTED_4548,SV2V_UNCONNECTED_4549,
  SV2V_UNCONNECTED_4550,SV2V_UNCONNECTED_4551,SV2V_UNCONNECTED_4552,
  SV2V_UNCONNECTED_4553,SV2V_UNCONNECTED_4554,SV2V_UNCONNECTED_4555,
  SV2V_UNCONNECTED_4556,SV2V_UNCONNECTED_4557,SV2V_UNCONNECTED_4558,
  SV2V_UNCONNECTED_4559,SV2V_UNCONNECTED_4560,SV2V_UNCONNECTED_4561,
  SV2V_UNCONNECTED_4562,SV2V_UNCONNECTED_4563,SV2V_UNCONNECTED_4564,
  SV2V_UNCONNECTED_4565,SV2V_UNCONNECTED_4566,SV2V_UNCONNECTED_4567,
  SV2V_UNCONNECTED_4568,SV2V_UNCONNECTED_4569,SV2V_UNCONNECTED_4570,
  SV2V_UNCONNECTED_4571,SV2V_UNCONNECTED_4572,SV2V_UNCONNECTED_4573,
  SV2V_UNCONNECTED_4574,SV2V_UNCONNECTED_4575,SV2V_UNCONNECTED_4576,SV2V_UNCONNECTED_4577,
  SV2V_UNCONNECTED_4578,SV2V_UNCONNECTED_4579,SV2V_UNCONNECTED_4580,
  SV2V_UNCONNECTED_4581,SV2V_UNCONNECTED_4582,SV2V_UNCONNECTED_4583,
  SV2V_UNCONNECTED_4584,SV2V_UNCONNECTED_4585,SV2V_UNCONNECTED_4586,
  SV2V_UNCONNECTED_4587,SV2V_UNCONNECTED_4588,SV2V_UNCONNECTED_4589,
  SV2V_UNCONNECTED_4590,SV2V_UNCONNECTED_4591,SV2V_UNCONNECTED_4592,
  SV2V_UNCONNECTED_4593,SV2V_UNCONNECTED_4594,SV2V_UNCONNECTED_4595,
  SV2V_UNCONNECTED_4596,SV2V_UNCONNECTED_4597,SV2V_UNCONNECTED_4598,
  SV2V_UNCONNECTED_4599,SV2V_UNCONNECTED_4600,SV2V_UNCONNECTED_4601,
  SV2V_UNCONNECTED_4602,SV2V_UNCONNECTED_4603,SV2V_UNCONNECTED_4604,
  SV2V_UNCONNECTED_4605,SV2V_UNCONNECTED_4606,SV2V_UNCONNECTED_4607,
  SV2V_UNCONNECTED_4608,SV2V_UNCONNECTED_4609,SV2V_UNCONNECTED_4610,
  SV2V_UNCONNECTED_4611,SV2V_UNCONNECTED_4612,SV2V_UNCONNECTED_4613,
  SV2V_UNCONNECTED_4614,SV2V_UNCONNECTED_4615,SV2V_UNCONNECTED_4616,SV2V_UNCONNECTED_4617,
  SV2V_UNCONNECTED_4618,SV2V_UNCONNECTED_4619,SV2V_UNCONNECTED_4620,
  SV2V_UNCONNECTED_4621,SV2V_UNCONNECTED_4622,SV2V_UNCONNECTED_4623,
  SV2V_UNCONNECTED_4624,SV2V_UNCONNECTED_4625,SV2V_UNCONNECTED_4626,
  SV2V_UNCONNECTED_4627,SV2V_UNCONNECTED_4628,SV2V_UNCONNECTED_4629,
  SV2V_UNCONNECTED_4630,SV2V_UNCONNECTED_4631,SV2V_UNCONNECTED_4632,
  SV2V_UNCONNECTED_4633,SV2V_UNCONNECTED_4634,SV2V_UNCONNECTED_4635,
  SV2V_UNCONNECTED_4636,SV2V_UNCONNECTED_4637,SV2V_UNCONNECTED_4638,
  SV2V_UNCONNECTED_4639,SV2V_UNCONNECTED_4640,SV2V_UNCONNECTED_4641,
  SV2V_UNCONNECTED_4642,SV2V_UNCONNECTED_4643,SV2V_UNCONNECTED_4644,
  SV2V_UNCONNECTED_4645,SV2V_UNCONNECTED_4646,SV2V_UNCONNECTED_4647,
  SV2V_UNCONNECTED_4648,SV2V_UNCONNECTED_4649,SV2V_UNCONNECTED_4650,
  SV2V_UNCONNECTED_4651,SV2V_UNCONNECTED_4652,SV2V_UNCONNECTED_4653,
  SV2V_UNCONNECTED_4654,SV2V_UNCONNECTED_4655,SV2V_UNCONNECTED_4656,SV2V_UNCONNECTED_4657,
  SV2V_UNCONNECTED_4658,SV2V_UNCONNECTED_4659,SV2V_UNCONNECTED_4660,
  SV2V_UNCONNECTED_4661,SV2V_UNCONNECTED_4662,SV2V_UNCONNECTED_4663,
  SV2V_UNCONNECTED_4664,SV2V_UNCONNECTED_4665,SV2V_UNCONNECTED_4666,
  SV2V_UNCONNECTED_4667,SV2V_UNCONNECTED_4668,SV2V_UNCONNECTED_4669,
  SV2V_UNCONNECTED_4670,SV2V_UNCONNECTED_4671,SV2V_UNCONNECTED_4672,
  SV2V_UNCONNECTED_4673,SV2V_UNCONNECTED_4674,SV2V_UNCONNECTED_4675,
  SV2V_UNCONNECTED_4676,SV2V_UNCONNECTED_4677,SV2V_UNCONNECTED_4678,
  SV2V_UNCONNECTED_4679,SV2V_UNCONNECTED_4680,SV2V_UNCONNECTED_4681,
  SV2V_UNCONNECTED_4682,SV2V_UNCONNECTED_4683,SV2V_UNCONNECTED_4684,
  SV2V_UNCONNECTED_4685,SV2V_UNCONNECTED_4686,SV2V_UNCONNECTED_4687,
  SV2V_UNCONNECTED_4688,SV2V_UNCONNECTED_4689,SV2V_UNCONNECTED_4690,
  SV2V_UNCONNECTED_4691,SV2V_UNCONNECTED_4692,SV2V_UNCONNECTED_4693,
  SV2V_UNCONNECTED_4694,SV2V_UNCONNECTED_4695,SV2V_UNCONNECTED_4696,SV2V_UNCONNECTED_4697,
  SV2V_UNCONNECTED_4698,SV2V_UNCONNECTED_4699,SV2V_UNCONNECTED_4700,
  SV2V_UNCONNECTED_4701,SV2V_UNCONNECTED_4702,SV2V_UNCONNECTED_4703,
  SV2V_UNCONNECTED_4704,SV2V_UNCONNECTED_4705,SV2V_UNCONNECTED_4706,
  SV2V_UNCONNECTED_4707,SV2V_UNCONNECTED_4708,SV2V_UNCONNECTED_4709,
  SV2V_UNCONNECTED_4710,SV2V_UNCONNECTED_4711,SV2V_UNCONNECTED_4712,
  SV2V_UNCONNECTED_4713,SV2V_UNCONNECTED_4714,SV2V_UNCONNECTED_4715,
  SV2V_UNCONNECTED_4716,SV2V_UNCONNECTED_4717,SV2V_UNCONNECTED_4718,
  SV2V_UNCONNECTED_4719,SV2V_UNCONNECTED_4720,SV2V_UNCONNECTED_4721,
  SV2V_UNCONNECTED_4722,SV2V_UNCONNECTED_4723,SV2V_UNCONNECTED_4724,
  SV2V_UNCONNECTED_4725,SV2V_UNCONNECTED_4726,SV2V_UNCONNECTED_4727,
  SV2V_UNCONNECTED_4728,SV2V_UNCONNECTED_4729,SV2V_UNCONNECTED_4730,
  SV2V_UNCONNECTED_4731,SV2V_UNCONNECTED_4732,SV2V_UNCONNECTED_4733,
  SV2V_UNCONNECTED_4734,SV2V_UNCONNECTED_4735,SV2V_UNCONNECTED_4736,SV2V_UNCONNECTED_4737,
  SV2V_UNCONNECTED_4738,SV2V_UNCONNECTED_4739,SV2V_UNCONNECTED_4740,
  SV2V_UNCONNECTED_4741,SV2V_UNCONNECTED_4742,SV2V_UNCONNECTED_4743,
  SV2V_UNCONNECTED_4744,SV2V_UNCONNECTED_4745,SV2V_UNCONNECTED_4746,
  SV2V_UNCONNECTED_4747,SV2V_UNCONNECTED_4748,SV2V_UNCONNECTED_4749,
  SV2V_UNCONNECTED_4750,SV2V_UNCONNECTED_4751,SV2V_UNCONNECTED_4752,
  SV2V_UNCONNECTED_4753,SV2V_UNCONNECTED_4754,SV2V_UNCONNECTED_4755,
  SV2V_UNCONNECTED_4756,SV2V_UNCONNECTED_4757,SV2V_UNCONNECTED_4758,
  SV2V_UNCONNECTED_4759,SV2V_UNCONNECTED_4760,SV2V_UNCONNECTED_4761,
  SV2V_UNCONNECTED_4762,SV2V_UNCONNECTED_4763,SV2V_UNCONNECTED_4764,
  SV2V_UNCONNECTED_4765,SV2V_UNCONNECTED_4766,SV2V_UNCONNECTED_4767,
  SV2V_UNCONNECTED_4768,SV2V_UNCONNECTED_4769,SV2V_UNCONNECTED_4770,
  SV2V_UNCONNECTED_4771,SV2V_UNCONNECTED_4772,SV2V_UNCONNECTED_4773,
  SV2V_UNCONNECTED_4774,SV2V_UNCONNECTED_4775,SV2V_UNCONNECTED_4776,SV2V_UNCONNECTED_4777,
  SV2V_UNCONNECTED_4778,SV2V_UNCONNECTED_4779,SV2V_UNCONNECTED_4780,
  SV2V_UNCONNECTED_4781,SV2V_UNCONNECTED_4782,SV2V_UNCONNECTED_4783,
  SV2V_UNCONNECTED_4784,SV2V_UNCONNECTED_4785,SV2V_UNCONNECTED_4786,
  SV2V_UNCONNECTED_4787,SV2V_UNCONNECTED_4788,SV2V_UNCONNECTED_4789,
  SV2V_UNCONNECTED_4790,SV2V_UNCONNECTED_4791,SV2V_UNCONNECTED_4792,
  SV2V_UNCONNECTED_4793,SV2V_UNCONNECTED_4794,SV2V_UNCONNECTED_4795,
  SV2V_UNCONNECTED_4796,SV2V_UNCONNECTED_4797,SV2V_UNCONNECTED_4798,
  SV2V_UNCONNECTED_4799,SV2V_UNCONNECTED_4800,SV2V_UNCONNECTED_4801,
  SV2V_UNCONNECTED_4802,SV2V_UNCONNECTED_4803,SV2V_UNCONNECTED_4804,
  SV2V_UNCONNECTED_4805,SV2V_UNCONNECTED_4806,SV2V_UNCONNECTED_4807,
  SV2V_UNCONNECTED_4808,SV2V_UNCONNECTED_4809,SV2V_UNCONNECTED_4810,
  SV2V_UNCONNECTED_4811,SV2V_UNCONNECTED_4812,SV2V_UNCONNECTED_4813,
  SV2V_UNCONNECTED_4814,SV2V_UNCONNECTED_4815,SV2V_UNCONNECTED_4816,SV2V_UNCONNECTED_4817,
  SV2V_UNCONNECTED_4818,SV2V_UNCONNECTED_4819,SV2V_UNCONNECTED_4820,
  SV2V_UNCONNECTED_4821,SV2V_UNCONNECTED_4822,SV2V_UNCONNECTED_4823,
  SV2V_UNCONNECTED_4824,SV2V_UNCONNECTED_4825,SV2V_UNCONNECTED_4826,
  SV2V_UNCONNECTED_4827,SV2V_UNCONNECTED_4828,SV2V_UNCONNECTED_4829,
  SV2V_UNCONNECTED_4830,SV2V_UNCONNECTED_4831,SV2V_UNCONNECTED_4832,
  SV2V_UNCONNECTED_4833,SV2V_UNCONNECTED_4834,SV2V_UNCONNECTED_4835,
  SV2V_UNCONNECTED_4836,SV2V_UNCONNECTED_4837,SV2V_UNCONNECTED_4838,
  SV2V_UNCONNECTED_4839,SV2V_UNCONNECTED_4840,SV2V_UNCONNECTED_4841,
  SV2V_UNCONNECTED_4842,SV2V_UNCONNECTED_4843,SV2V_UNCONNECTED_4844,
  SV2V_UNCONNECTED_4845,SV2V_UNCONNECTED_4846,SV2V_UNCONNECTED_4847,
  SV2V_UNCONNECTED_4848,SV2V_UNCONNECTED_4849,SV2V_UNCONNECTED_4850,
  SV2V_UNCONNECTED_4851,SV2V_UNCONNECTED_4852,SV2V_UNCONNECTED_4853,
  SV2V_UNCONNECTED_4854,SV2V_UNCONNECTED_4855,SV2V_UNCONNECTED_4856,SV2V_UNCONNECTED_4857,
  SV2V_UNCONNECTED_4858,SV2V_UNCONNECTED_4859,SV2V_UNCONNECTED_4860,
  SV2V_UNCONNECTED_4861,SV2V_UNCONNECTED_4862,SV2V_UNCONNECTED_4863,
  SV2V_UNCONNECTED_4864,SV2V_UNCONNECTED_4865,SV2V_UNCONNECTED_4866,
  SV2V_UNCONNECTED_4867,SV2V_UNCONNECTED_4868,SV2V_UNCONNECTED_4869,
  SV2V_UNCONNECTED_4870,SV2V_UNCONNECTED_4871,SV2V_UNCONNECTED_4872,
  SV2V_UNCONNECTED_4873,SV2V_UNCONNECTED_4874,SV2V_UNCONNECTED_4875,
  SV2V_UNCONNECTED_4876,SV2V_UNCONNECTED_4877,SV2V_UNCONNECTED_4878,
  SV2V_UNCONNECTED_4879,SV2V_UNCONNECTED_4880,SV2V_UNCONNECTED_4881,
  SV2V_UNCONNECTED_4882,SV2V_UNCONNECTED_4883,SV2V_UNCONNECTED_4884,
  SV2V_UNCONNECTED_4885,SV2V_UNCONNECTED_4886,SV2V_UNCONNECTED_4887,
  SV2V_UNCONNECTED_4888,SV2V_UNCONNECTED_4889,SV2V_UNCONNECTED_4890,
  SV2V_UNCONNECTED_4891,SV2V_UNCONNECTED_4892,SV2V_UNCONNECTED_4893,
  SV2V_UNCONNECTED_4894,SV2V_UNCONNECTED_4895,SV2V_UNCONNECTED_4896,SV2V_UNCONNECTED_4897,
  SV2V_UNCONNECTED_4898,SV2V_UNCONNECTED_4899,SV2V_UNCONNECTED_4900,
  SV2V_UNCONNECTED_4901,SV2V_UNCONNECTED_4902,SV2V_UNCONNECTED_4903,
  SV2V_UNCONNECTED_4904,SV2V_UNCONNECTED_4905,SV2V_UNCONNECTED_4906,
  SV2V_UNCONNECTED_4907,SV2V_UNCONNECTED_4908,SV2V_UNCONNECTED_4909,
  SV2V_UNCONNECTED_4910,SV2V_UNCONNECTED_4911,SV2V_UNCONNECTED_4912,
  SV2V_UNCONNECTED_4913,SV2V_UNCONNECTED_4914,SV2V_UNCONNECTED_4915,
  SV2V_UNCONNECTED_4916,SV2V_UNCONNECTED_4917,SV2V_UNCONNECTED_4918,
  SV2V_UNCONNECTED_4919,SV2V_UNCONNECTED_4920,SV2V_UNCONNECTED_4921,
  SV2V_UNCONNECTED_4922,SV2V_UNCONNECTED_4923,SV2V_UNCONNECTED_4924,
  SV2V_UNCONNECTED_4925,SV2V_UNCONNECTED_4926,SV2V_UNCONNECTED_4927,
  SV2V_UNCONNECTED_4928,SV2V_UNCONNECTED_4929,SV2V_UNCONNECTED_4930,
  SV2V_UNCONNECTED_4931,SV2V_UNCONNECTED_4932,SV2V_UNCONNECTED_4933,
  SV2V_UNCONNECTED_4934,SV2V_UNCONNECTED_4935,SV2V_UNCONNECTED_4936,SV2V_UNCONNECTED_4937,
  SV2V_UNCONNECTED_4938,SV2V_UNCONNECTED_4939,SV2V_UNCONNECTED_4940,
  SV2V_UNCONNECTED_4941,SV2V_UNCONNECTED_4942,SV2V_UNCONNECTED_4943,
  SV2V_UNCONNECTED_4944,SV2V_UNCONNECTED_4945,SV2V_UNCONNECTED_4946,
  SV2V_UNCONNECTED_4947,SV2V_UNCONNECTED_4948,SV2V_UNCONNECTED_4949,
  SV2V_UNCONNECTED_4950,SV2V_UNCONNECTED_4951,SV2V_UNCONNECTED_4952,
  SV2V_UNCONNECTED_4953,SV2V_UNCONNECTED_4954,SV2V_UNCONNECTED_4955,
  SV2V_UNCONNECTED_4956,SV2V_UNCONNECTED_4957,SV2V_UNCONNECTED_4958,
  SV2V_UNCONNECTED_4959,SV2V_UNCONNECTED_4960,SV2V_UNCONNECTED_4961,
  SV2V_UNCONNECTED_4962,SV2V_UNCONNECTED_4963,SV2V_UNCONNECTED_4964,
  SV2V_UNCONNECTED_4965,SV2V_UNCONNECTED_4966,SV2V_UNCONNECTED_4967,
  SV2V_UNCONNECTED_4968,SV2V_UNCONNECTED_4969,SV2V_UNCONNECTED_4970,
  SV2V_UNCONNECTED_4971,SV2V_UNCONNECTED_4972,SV2V_UNCONNECTED_4973,
  SV2V_UNCONNECTED_4974,SV2V_UNCONNECTED_4975,SV2V_UNCONNECTED_4976,SV2V_UNCONNECTED_4977,
  SV2V_UNCONNECTED_4978,SV2V_UNCONNECTED_4979,SV2V_UNCONNECTED_4980,
  SV2V_UNCONNECTED_4981,SV2V_UNCONNECTED_4982,SV2V_UNCONNECTED_4983,
  SV2V_UNCONNECTED_4984,SV2V_UNCONNECTED_4985,SV2V_UNCONNECTED_4986,
  SV2V_UNCONNECTED_4987,SV2V_UNCONNECTED_4988,SV2V_UNCONNECTED_4989,
  SV2V_UNCONNECTED_4990,SV2V_UNCONNECTED_4991,SV2V_UNCONNECTED_4992,
  SV2V_UNCONNECTED_4993,SV2V_UNCONNECTED_4994,SV2V_UNCONNECTED_4995,
  SV2V_UNCONNECTED_4996,SV2V_UNCONNECTED_4997,SV2V_UNCONNECTED_4998,
  SV2V_UNCONNECTED_4999,SV2V_UNCONNECTED_5000,SV2V_UNCONNECTED_5001,
  SV2V_UNCONNECTED_5002,SV2V_UNCONNECTED_5003,SV2V_UNCONNECTED_5004,
  SV2V_UNCONNECTED_5005,SV2V_UNCONNECTED_5006,SV2V_UNCONNECTED_5007,
  SV2V_UNCONNECTED_5008,SV2V_UNCONNECTED_5009,SV2V_UNCONNECTED_5010,
  SV2V_UNCONNECTED_5011,SV2V_UNCONNECTED_5012,SV2V_UNCONNECTED_5013,
  SV2V_UNCONNECTED_5014,SV2V_UNCONNECTED_5015,SV2V_UNCONNECTED_5016,SV2V_UNCONNECTED_5017,
  SV2V_UNCONNECTED_5018,SV2V_UNCONNECTED_5019,SV2V_UNCONNECTED_5020,
  SV2V_UNCONNECTED_5021,SV2V_UNCONNECTED_5022,SV2V_UNCONNECTED_5023,
  SV2V_UNCONNECTED_5024,SV2V_UNCONNECTED_5025,SV2V_UNCONNECTED_5026,
  SV2V_UNCONNECTED_5027,SV2V_UNCONNECTED_5028,SV2V_UNCONNECTED_5029,
  SV2V_UNCONNECTED_5030,SV2V_UNCONNECTED_5031,SV2V_UNCONNECTED_5032,
  SV2V_UNCONNECTED_5033,SV2V_UNCONNECTED_5034,SV2V_UNCONNECTED_5035,
  SV2V_UNCONNECTED_5036,SV2V_UNCONNECTED_5037,SV2V_UNCONNECTED_5038,
  SV2V_UNCONNECTED_5039,SV2V_UNCONNECTED_5040,SV2V_UNCONNECTED_5041,
  SV2V_UNCONNECTED_5042,SV2V_UNCONNECTED_5043,SV2V_UNCONNECTED_5044,
  SV2V_UNCONNECTED_5045,SV2V_UNCONNECTED_5046,SV2V_UNCONNECTED_5047,
  SV2V_UNCONNECTED_5048,SV2V_UNCONNECTED_5049,SV2V_UNCONNECTED_5050,
  SV2V_UNCONNECTED_5051,SV2V_UNCONNECTED_5052,SV2V_UNCONNECTED_5053,
  SV2V_UNCONNECTED_5054,SV2V_UNCONNECTED_5055,SV2V_UNCONNECTED_5056,SV2V_UNCONNECTED_5057,
  SV2V_UNCONNECTED_5058,SV2V_UNCONNECTED_5059,SV2V_UNCONNECTED_5060,
  SV2V_UNCONNECTED_5061,SV2V_UNCONNECTED_5062,SV2V_UNCONNECTED_5063,
  SV2V_UNCONNECTED_5064,SV2V_UNCONNECTED_5065,SV2V_UNCONNECTED_5066,
  SV2V_UNCONNECTED_5067,SV2V_UNCONNECTED_5068,SV2V_UNCONNECTED_5069,
  SV2V_UNCONNECTED_5070,SV2V_UNCONNECTED_5071,SV2V_UNCONNECTED_5072,
  SV2V_UNCONNECTED_5073,SV2V_UNCONNECTED_5074,SV2V_UNCONNECTED_5075,
  SV2V_UNCONNECTED_5076,SV2V_UNCONNECTED_5077,SV2V_UNCONNECTED_5078,
  SV2V_UNCONNECTED_5079,SV2V_UNCONNECTED_5080,SV2V_UNCONNECTED_5081,
  SV2V_UNCONNECTED_5082,SV2V_UNCONNECTED_5083,SV2V_UNCONNECTED_5084,
  SV2V_UNCONNECTED_5085,SV2V_UNCONNECTED_5086,SV2V_UNCONNECTED_5087,
  SV2V_UNCONNECTED_5088,SV2V_UNCONNECTED_5089,SV2V_UNCONNECTED_5090,
  SV2V_UNCONNECTED_5091,SV2V_UNCONNECTED_5092,SV2V_UNCONNECTED_5093,
  SV2V_UNCONNECTED_5094,SV2V_UNCONNECTED_5095,SV2V_UNCONNECTED_5096,SV2V_UNCONNECTED_5097,
  SV2V_UNCONNECTED_5098,SV2V_UNCONNECTED_5099,SV2V_UNCONNECTED_5100,
  SV2V_UNCONNECTED_5101,SV2V_UNCONNECTED_5102,SV2V_UNCONNECTED_5103,
  SV2V_UNCONNECTED_5104,SV2V_UNCONNECTED_5105,SV2V_UNCONNECTED_5106,
  SV2V_UNCONNECTED_5107,SV2V_UNCONNECTED_5108,SV2V_UNCONNECTED_5109,
  SV2V_UNCONNECTED_5110,SV2V_UNCONNECTED_5111,SV2V_UNCONNECTED_5112,
  SV2V_UNCONNECTED_5113,SV2V_UNCONNECTED_5114,SV2V_UNCONNECTED_5115,
  SV2V_UNCONNECTED_5116,SV2V_UNCONNECTED_5117,SV2V_UNCONNECTED_5118,
  SV2V_UNCONNECTED_5119,SV2V_UNCONNECTED_5120,SV2V_UNCONNECTED_5121,
  SV2V_UNCONNECTED_5122,SV2V_UNCONNECTED_5123,SV2V_UNCONNECTED_5124,
  SV2V_UNCONNECTED_5125,SV2V_UNCONNECTED_5126,SV2V_UNCONNECTED_5127,
  SV2V_UNCONNECTED_5128,SV2V_UNCONNECTED_5129,SV2V_UNCONNECTED_5130,
  SV2V_UNCONNECTED_5131,SV2V_UNCONNECTED_5132,SV2V_UNCONNECTED_5133,
  SV2V_UNCONNECTED_5134,SV2V_UNCONNECTED_5135,SV2V_UNCONNECTED_5136,SV2V_UNCONNECTED_5137,
  SV2V_UNCONNECTED_5138,SV2V_UNCONNECTED_5139,SV2V_UNCONNECTED_5140,
  SV2V_UNCONNECTED_5141,SV2V_UNCONNECTED_5142,SV2V_UNCONNECTED_5143,
  SV2V_UNCONNECTED_5144,SV2V_UNCONNECTED_5145,SV2V_UNCONNECTED_5146,
  SV2V_UNCONNECTED_5147,SV2V_UNCONNECTED_5148,SV2V_UNCONNECTED_5149,
  SV2V_UNCONNECTED_5150,SV2V_UNCONNECTED_5151,SV2V_UNCONNECTED_5152,
  SV2V_UNCONNECTED_5153,SV2V_UNCONNECTED_5154,SV2V_UNCONNECTED_5155,
  SV2V_UNCONNECTED_5156,SV2V_UNCONNECTED_5157,SV2V_UNCONNECTED_5158,
  SV2V_UNCONNECTED_5159,SV2V_UNCONNECTED_5160,SV2V_UNCONNECTED_5161,
  SV2V_UNCONNECTED_5162,SV2V_UNCONNECTED_5163,SV2V_UNCONNECTED_5164,
  SV2V_UNCONNECTED_5165,SV2V_UNCONNECTED_5166,SV2V_UNCONNECTED_5167,
  SV2V_UNCONNECTED_5168,SV2V_UNCONNECTED_5169,SV2V_UNCONNECTED_5170,
  SV2V_UNCONNECTED_5171,SV2V_UNCONNECTED_5172,SV2V_UNCONNECTED_5173,
  SV2V_UNCONNECTED_5174,SV2V_UNCONNECTED_5175,SV2V_UNCONNECTED_5176,SV2V_UNCONNECTED_5177,
  SV2V_UNCONNECTED_5178,SV2V_UNCONNECTED_5179,SV2V_UNCONNECTED_5180,
  SV2V_UNCONNECTED_5181,SV2V_UNCONNECTED_5182,SV2V_UNCONNECTED_5183,
  SV2V_UNCONNECTED_5184,SV2V_UNCONNECTED_5185,SV2V_UNCONNECTED_5186,
  SV2V_UNCONNECTED_5187,SV2V_UNCONNECTED_5188,SV2V_UNCONNECTED_5189,
  SV2V_UNCONNECTED_5190,SV2V_UNCONNECTED_5191,SV2V_UNCONNECTED_5192,
  SV2V_UNCONNECTED_5193,SV2V_UNCONNECTED_5194,SV2V_UNCONNECTED_5195,
  SV2V_UNCONNECTED_5196,SV2V_UNCONNECTED_5197,SV2V_UNCONNECTED_5198,
  SV2V_UNCONNECTED_5199,SV2V_UNCONNECTED_5200,SV2V_UNCONNECTED_5201,
  SV2V_UNCONNECTED_5202,SV2V_UNCONNECTED_5203,SV2V_UNCONNECTED_5204,
  SV2V_UNCONNECTED_5205,SV2V_UNCONNECTED_5206,SV2V_UNCONNECTED_5207,
  SV2V_UNCONNECTED_5208,SV2V_UNCONNECTED_5209,SV2V_UNCONNECTED_5210,
  SV2V_UNCONNECTED_5211,SV2V_UNCONNECTED_5212,SV2V_UNCONNECTED_5213,
  SV2V_UNCONNECTED_5214,SV2V_UNCONNECTED_5215,SV2V_UNCONNECTED_5216,SV2V_UNCONNECTED_5217,
  SV2V_UNCONNECTED_5218,SV2V_UNCONNECTED_5219,SV2V_UNCONNECTED_5220,
  SV2V_UNCONNECTED_5221,SV2V_UNCONNECTED_5222,SV2V_UNCONNECTED_5223,
  SV2V_UNCONNECTED_5224,SV2V_UNCONNECTED_5225,SV2V_UNCONNECTED_5226,
  SV2V_UNCONNECTED_5227,SV2V_UNCONNECTED_5228,SV2V_UNCONNECTED_5229,
  SV2V_UNCONNECTED_5230,SV2V_UNCONNECTED_5231,SV2V_UNCONNECTED_5232,
  SV2V_UNCONNECTED_5233,SV2V_UNCONNECTED_5234,SV2V_UNCONNECTED_5235,
  SV2V_UNCONNECTED_5236,SV2V_UNCONNECTED_5237,SV2V_UNCONNECTED_5238,
  SV2V_UNCONNECTED_5239,SV2V_UNCONNECTED_5240,SV2V_UNCONNECTED_5241,
  SV2V_UNCONNECTED_5242,SV2V_UNCONNECTED_5243,SV2V_UNCONNECTED_5244,
  SV2V_UNCONNECTED_5245,SV2V_UNCONNECTED_5246,SV2V_UNCONNECTED_5247,
  SV2V_UNCONNECTED_5248,SV2V_UNCONNECTED_5249,SV2V_UNCONNECTED_5250,
  SV2V_UNCONNECTED_5251,SV2V_UNCONNECTED_5252,SV2V_UNCONNECTED_5253,
  SV2V_UNCONNECTED_5254,SV2V_UNCONNECTED_5255,SV2V_UNCONNECTED_5256,SV2V_UNCONNECTED_5257,
  SV2V_UNCONNECTED_5258,SV2V_UNCONNECTED_5259,SV2V_UNCONNECTED_5260,
  SV2V_UNCONNECTED_5261,SV2V_UNCONNECTED_5262,SV2V_UNCONNECTED_5263,
  SV2V_UNCONNECTED_5264,SV2V_UNCONNECTED_5265,SV2V_UNCONNECTED_5266,
  SV2V_UNCONNECTED_5267,SV2V_UNCONNECTED_5268,SV2V_UNCONNECTED_5269,
  SV2V_UNCONNECTED_5270,SV2V_UNCONNECTED_5271,SV2V_UNCONNECTED_5272,
  SV2V_UNCONNECTED_5273,SV2V_UNCONNECTED_5274,SV2V_UNCONNECTED_5275,
  SV2V_UNCONNECTED_5276,SV2V_UNCONNECTED_5277,SV2V_UNCONNECTED_5278,
  SV2V_UNCONNECTED_5279,SV2V_UNCONNECTED_5280,SV2V_UNCONNECTED_5281,
  SV2V_UNCONNECTED_5282,SV2V_UNCONNECTED_5283,SV2V_UNCONNECTED_5284,
  SV2V_UNCONNECTED_5285,SV2V_UNCONNECTED_5286,SV2V_UNCONNECTED_5287,
  SV2V_UNCONNECTED_5288,SV2V_UNCONNECTED_5289,SV2V_UNCONNECTED_5290,
  SV2V_UNCONNECTED_5291,SV2V_UNCONNECTED_5292,SV2V_UNCONNECTED_5293,
  SV2V_UNCONNECTED_5294,SV2V_UNCONNECTED_5295,SV2V_UNCONNECTED_5296,SV2V_UNCONNECTED_5297,
  SV2V_UNCONNECTED_5298,SV2V_UNCONNECTED_5299,SV2V_UNCONNECTED_5300,
  SV2V_UNCONNECTED_5301,SV2V_UNCONNECTED_5302,SV2V_UNCONNECTED_5303,
  SV2V_UNCONNECTED_5304,SV2V_UNCONNECTED_5305,SV2V_UNCONNECTED_5306,
  SV2V_UNCONNECTED_5307,SV2V_UNCONNECTED_5308,SV2V_UNCONNECTED_5309,
  SV2V_UNCONNECTED_5310,SV2V_UNCONNECTED_5311,SV2V_UNCONNECTED_5312,
  SV2V_UNCONNECTED_5313,SV2V_UNCONNECTED_5314,SV2V_UNCONNECTED_5315,
  SV2V_UNCONNECTED_5316,SV2V_UNCONNECTED_5317,SV2V_UNCONNECTED_5318,
  SV2V_UNCONNECTED_5319,SV2V_UNCONNECTED_5320,SV2V_UNCONNECTED_5321,
  SV2V_UNCONNECTED_5322,SV2V_UNCONNECTED_5323,SV2V_UNCONNECTED_5324,
  SV2V_UNCONNECTED_5325,SV2V_UNCONNECTED_5326,SV2V_UNCONNECTED_5327,
  SV2V_UNCONNECTED_5328,SV2V_UNCONNECTED_5329,SV2V_UNCONNECTED_5330,
  SV2V_UNCONNECTED_5331,SV2V_UNCONNECTED_5332,SV2V_UNCONNECTED_5333,
  SV2V_UNCONNECTED_5334,SV2V_UNCONNECTED_5335,SV2V_UNCONNECTED_5336,SV2V_UNCONNECTED_5337,
  SV2V_UNCONNECTED_5338,SV2V_UNCONNECTED_5339,SV2V_UNCONNECTED_5340,
  SV2V_UNCONNECTED_5341,SV2V_UNCONNECTED_5342,SV2V_UNCONNECTED_5343,
  SV2V_UNCONNECTED_5344,SV2V_UNCONNECTED_5345,SV2V_UNCONNECTED_5346,
  SV2V_UNCONNECTED_5347,SV2V_UNCONNECTED_5348,SV2V_UNCONNECTED_5349,
  SV2V_UNCONNECTED_5350,SV2V_UNCONNECTED_5351,SV2V_UNCONNECTED_5352,
  SV2V_UNCONNECTED_5353,SV2V_UNCONNECTED_5354,SV2V_UNCONNECTED_5355,
  SV2V_UNCONNECTED_5356,SV2V_UNCONNECTED_5357,SV2V_UNCONNECTED_5358,
  SV2V_UNCONNECTED_5359,SV2V_UNCONNECTED_5360,SV2V_UNCONNECTED_5361,
  SV2V_UNCONNECTED_5362,SV2V_UNCONNECTED_5363,SV2V_UNCONNECTED_5364,
  SV2V_UNCONNECTED_5365,SV2V_UNCONNECTED_5366,SV2V_UNCONNECTED_5367,
  SV2V_UNCONNECTED_5368,SV2V_UNCONNECTED_5369,SV2V_UNCONNECTED_5370,
  SV2V_UNCONNECTED_5371,SV2V_UNCONNECTED_5372,SV2V_UNCONNECTED_5373,
  SV2V_UNCONNECTED_5374,SV2V_UNCONNECTED_5375,SV2V_UNCONNECTED_5376,SV2V_UNCONNECTED_5377,
  SV2V_UNCONNECTED_5378,SV2V_UNCONNECTED_5379,SV2V_UNCONNECTED_5380,
  SV2V_UNCONNECTED_5381,SV2V_UNCONNECTED_5382,SV2V_UNCONNECTED_5383,
  SV2V_UNCONNECTED_5384,SV2V_UNCONNECTED_5385,SV2V_UNCONNECTED_5386,
  SV2V_UNCONNECTED_5387,SV2V_UNCONNECTED_5388,SV2V_UNCONNECTED_5389,
  SV2V_UNCONNECTED_5390,SV2V_UNCONNECTED_5391,SV2V_UNCONNECTED_5392,
  SV2V_UNCONNECTED_5393,SV2V_UNCONNECTED_5394,SV2V_UNCONNECTED_5395,
  SV2V_UNCONNECTED_5396,SV2V_UNCONNECTED_5397,SV2V_UNCONNECTED_5398,
  SV2V_UNCONNECTED_5399,SV2V_UNCONNECTED_5400,SV2V_UNCONNECTED_5401,
  SV2V_UNCONNECTED_5402,SV2V_UNCONNECTED_5403,SV2V_UNCONNECTED_5404,
  SV2V_UNCONNECTED_5405,SV2V_UNCONNECTED_5406,SV2V_UNCONNECTED_5407,
  SV2V_UNCONNECTED_5408,SV2V_UNCONNECTED_5409,SV2V_UNCONNECTED_5410,
  SV2V_UNCONNECTED_5411,SV2V_UNCONNECTED_5412,SV2V_UNCONNECTED_5413,
  SV2V_UNCONNECTED_5414,SV2V_UNCONNECTED_5415,SV2V_UNCONNECTED_5416,SV2V_UNCONNECTED_5417,
  SV2V_UNCONNECTED_5418,SV2V_UNCONNECTED_5419,SV2V_UNCONNECTED_5420,
  SV2V_UNCONNECTED_5421,SV2V_UNCONNECTED_5422,SV2V_UNCONNECTED_5423,
  SV2V_UNCONNECTED_5424,SV2V_UNCONNECTED_5425,SV2V_UNCONNECTED_5426,
  SV2V_UNCONNECTED_5427,SV2V_UNCONNECTED_5428,SV2V_UNCONNECTED_5429,
  SV2V_UNCONNECTED_5430,SV2V_UNCONNECTED_5431,SV2V_UNCONNECTED_5432,
  SV2V_UNCONNECTED_5433,SV2V_UNCONNECTED_5434,SV2V_UNCONNECTED_5435,
  SV2V_UNCONNECTED_5436,SV2V_UNCONNECTED_5437,SV2V_UNCONNECTED_5438,
  SV2V_UNCONNECTED_5439,SV2V_UNCONNECTED_5440,SV2V_UNCONNECTED_5441,
  SV2V_UNCONNECTED_5442,SV2V_UNCONNECTED_5443,SV2V_UNCONNECTED_5444,
  SV2V_UNCONNECTED_5445,SV2V_UNCONNECTED_5446,SV2V_UNCONNECTED_5447,
  SV2V_UNCONNECTED_5448,SV2V_UNCONNECTED_5449,SV2V_UNCONNECTED_5450,
  SV2V_UNCONNECTED_5451,SV2V_UNCONNECTED_5452,SV2V_UNCONNECTED_5453,
  SV2V_UNCONNECTED_5454,SV2V_UNCONNECTED_5455,SV2V_UNCONNECTED_5456,SV2V_UNCONNECTED_5457,
  SV2V_UNCONNECTED_5458,SV2V_UNCONNECTED_5459,SV2V_UNCONNECTED_5460,
  SV2V_UNCONNECTED_5461,SV2V_UNCONNECTED_5462,SV2V_UNCONNECTED_5463,
  SV2V_UNCONNECTED_5464,SV2V_UNCONNECTED_5465,SV2V_UNCONNECTED_5466,
  SV2V_UNCONNECTED_5467,SV2V_UNCONNECTED_5468,SV2V_UNCONNECTED_5469,
  SV2V_UNCONNECTED_5470,SV2V_UNCONNECTED_5471,SV2V_UNCONNECTED_5472,
  SV2V_UNCONNECTED_5473,SV2V_UNCONNECTED_5474,SV2V_UNCONNECTED_5475,
  SV2V_UNCONNECTED_5476,SV2V_UNCONNECTED_5477,SV2V_UNCONNECTED_5478,
  SV2V_UNCONNECTED_5479,SV2V_UNCONNECTED_5480,SV2V_UNCONNECTED_5481,
  SV2V_UNCONNECTED_5482,SV2V_UNCONNECTED_5483,SV2V_UNCONNECTED_5484,
  SV2V_UNCONNECTED_5485,SV2V_UNCONNECTED_5486,SV2V_UNCONNECTED_5487,
  SV2V_UNCONNECTED_5488,SV2V_UNCONNECTED_5489,SV2V_UNCONNECTED_5490,
  SV2V_UNCONNECTED_5491,SV2V_UNCONNECTED_5492,SV2V_UNCONNECTED_5493,
  SV2V_UNCONNECTED_5494,SV2V_UNCONNECTED_5495,SV2V_UNCONNECTED_5496,SV2V_UNCONNECTED_5497,
  SV2V_UNCONNECTED_5498,SV2V_UNCONNECTED_5499,SV2V_UNCONNECTED_5500,
  SV2V_UNCONNECTED_5501,SV2V_UNCONNECTED_5502,SV2V_UNCONNECTED_5503,
  SV2V_UNCONNECTED_5504,SV2V_UNCONNECTED_5505,SV2V_UNCONNECTED_5506,
  SV2V_UNCONNECTED_5507,SV2V_UNCONNECTED_5508,SV2V_UNCONNECTED_5509,
  SV2V_UNCONNECTED_5510,SV2V_UNCONNECTED_5511,SV2V_UNCONNECTED_5512,
  SV2V_UNCONNECTED_5513,SV2V_UNCONNECTED_5514,SV2V_UNCONNECTED_5515,
  SV2V_UNCONNECTED_5516,SV2V_UNCONNECTED_5517,SV2V_UNCONNECTED_5518,
  SV2V_UNCONNECTED_5519,SV2V_UNCONNECTED_5520,SV2V_UNCONNECTED_5521,
  SV2V_UNCONNECTED_5522,SV2V_UNCONNECTED_5523,SV2V_UNCONNECTED_5524,
  SV2V_UNCONNECTED_5525,SV2V_UNCONNECTED_5526,SV2V_UNCONNECTED_5527,
  SV2V_UNCONNECTED_5528,SV2V_UNCONNECTED_5529,SV2V_UNCONNECTED_5530,
  SV2V_UNCONNECTED_5531,SV2V_UNCONNECTED_5532,SV2V_UNCONNECTED_5533,
  SV2V_UNCONNECTED_5534,SV2V_UNCONNECTED_5535,SV2V_UNCONNECTED_5536,SV2V_UNCONNECTED_5537,
  SV2V_UNCONNECTED_5538,SV2V_UNCONNECTED_5539,SV2V_UNCONNECTED_5540,
  SV2V_UNCONNECTED_5541,SV2V_UNCONNECTED_5542,SV2V_UNCONNECTED_5543,
  SV2V_UNCONNECTED_5544,SV2V_UNCONNECTED_5545,SV2V_UNCONNECTED_5546,
  SV2V_UNCONNECTED_5547,SV2V_UNCONNECTED_5548,SV2V_UNCONNECTED_5549,
  SV2V_UNCONNECTED_5550,SV2V_UNCONNECTED_5551,SV2V_UNCONNECTED_5552,
  SV2V_UNCONNECTED_5553,SV2V_UNCONNECTED_5554,SV2V_UNCONNECTED_5555,
  SV2V_UNCONNECTED_5556,SV2V_UNCONNECTED_5557,SV2V_UNCONNECTED_5558,
  SV2V_UNCONNECTED_5559,SV2V_UNCONNECTED_5560,SV2V_UNCONNECTED_5561,
  SV2V_UNCONNECTED_5562,SV2V_UNCONNECTED_5563,SV2V_UNCONNECTED_5564,
  SV2V_UNCONNECTED_5565,SV2V_UNCONNECTED_5566,SV2V_UNCONNECTED_5567,
  SV2V_UNCONNECTED_5568,SV2V_UNCONNECTED_5569,SV2V_UNCONNECTED_5570,
  SV2V_UNCONNECTED_5571,SV2V_UNCONNECTED_5572,SV2V_UNCONNECTED_5573,
  SV2V_UNCONNECTED_5574,SV2V_UNCONNECTED_5575,SV2V_UNCONNECTED_5576,SV2V_UNCONNECTED_5577,
  SV2V_UNCONNECTED_5578,SV2V_UNCONNECTED_5579,SV2V_UNCONNECTED_5580,
  SV2V_UNCONNECTED_5581,SV2V_UNCONNECTED_5582,SV2V_UNCONNECTED_5583,
  SV2V_UNCONNECTED_5584,SV2V_UNCONNECTED_5585,SV2V_UNCONNECTED_5586,
  SV2V_UNCONNECTED_5587,SV2V_UNCONNECTED_5588,SV2V_UNCONNECTED_5589,
  SV2V_UNCONNECTED_5590,SV2V_UNCONNECTED_5591,SV2V_UNCONNECTED_5592,
  SV2V_UNCONNECTED_5593,SV2V_UNCONNECTED_5594,SV2V_UNCONNECTED_5595,
  SV2V_UNCONNECTED_5596,SV2V_UNCONNECTED_5597,SV2V_UNCONNECTED_5598,
  SV2V_UNCONNECTED_5599,SV2V_UNCONNECTED_5600,SV2V_UNCONNECTED_5601,
  SV2V_UNCONNECTED_5602,SV2V_UNCONNECTED_5603,SV2V_UNCONNECTED_5604,
  SV2V_UNCONNECTED_5605,SV2V_UNCONNECTED_5606,SV2V_UNCONNECTED_5607,
  SV2V_UNCONNECTED_5608,SV2V_UNCONNECTED_5609,SV2V_UNCONNECTED_5610,
  SV2V_UNCONNECTED_5611,SV2V_UNCONNECTED_5612,SV2V_UNCONNECTED_5613,
  SV2V_UNCONNECTED_5614,SV2V_UNCONNECTED_5615,SV2V_UNCONNECTED_5616,SV2V_UNCONNECTED_5617,
  SV2V_UNCONNECTED_5618,SV2V_UNCONNECTED_5619,SV2V_UNCONNECTED_5620,
  SV2V_UNCONNECTED_5621,SV2V_UNCONNECTED_5622,SV2V_UNCONNECTED_5623,
  SV2V_UNCONNECTED_5624,SV2V_UNCONNECTED_5625,SV2V_UNCONNECTED_5626,
  SV2V_UNCONNECTED_5627,SV2V_UNCONNECTED_5628,SV2V_UNCONNECTED_5629,
  SV2V_UNCONNECTED_5630,SV2V_UNCONNECTED_5631,SV2V_UNCONNECTED_5632,
  SV2V_UNCONNECTED_5633,SV2V_UNCONNECTED_5634,SV2V_UNCONNECTED_5635,
  SV2V_UNCONNECTED_5636,SV2V_UNCONNECTED_5637,SV2V_UNCONNECTED_5638,
  SV2V_UNCONNECTED_5639,SV2V_UNCONNECTED_5640,SV2V_UNCONNECTED_5641,
  SV2V_UNCONNECTED_5642,SV2V_UNCONNECTED_5643,SV2V_UNCONNECTED_5644,
  SV2V_UNCONNECTED_5645,SV2V_UNCONNECTED_5646,SV2V_UNCONNECTED_5647,
  SV2V_UNCONNECTED_5648,SV2V_UNCONNECTED_5649,SV2V_UNCONNECTED_5650,
  SV2V_UNCONNECTED_5651,SV2V_UNCONNECTED_5652,SV2V_UNCONNECTED_5653,
  SV2V_UNCONNECTED_5654,SV2V_UNCONNECTED_5655,SV2V_UNCONNECTED_5656,SV2V_UNCONNECTED_5657,
  SV2V_UNCONNECTED_5658,SV2V_UNCONNECTED_5659,SV2V_UNCONNECTED_5660,
  SV2V_UNCONNECTED_5661,SV2V_UNCONNECTED_5662,SV2V_UNCONNECTED_5663,
  SV2V_UNCONNECTED_5664,SV2V_UNCONNECTED_5665,SV2V_UNCONNECTED_5666,
  SV2V_UNCONNECTED_5667,SV2V_UNCONNECTED_5668,SV2V_UNCONNECTED_5669,
  SV2V_UNCONNECTED_5670,SV2V_UNCONNECTED_5671,SV2V_UNCONNECTED_5672,
  SV2V_UNCONNECTED_5673,SV2V_UNCONNECTED_5674,SV2V_UNCONNECTED_5675,
  SV2V_UNCONNECTED_5676,SV2V_UNCONNECTED_5677,SV2V_UNCONNECTED_5678,
  SV2V_UNCONNECTED_5679,SV2V_UNCONNECTED_5680,SV2V_UNCONNECTED_5681,
  SV2V_UNCONNECTED_5682,SV2V_UNCONNECTED_5683,SV2V_UNCONNECTED_5684,
  SV2V_UNCONNECTED_5685,SV2V_UNCONNECTED_5686,SV2V_UNCONNECTED_5687,
  SV2V_UNCONNECTED_5688,SV2V_UNCONNECTED_5689,SV2V_UNCONNECTED_5690,
  SV2V_UNCONNECTED_5691,SV2V_UNCONNECTED_5692,SV2V_UNCONNECTED_5693,
  SV2V_UNCONNECTED_5694,SV2V_UNCONNECTED_5695,SV2V_UNCONNECTED_5696,SV2V_UNCONNECTED_5697,
  SV2V_UNCONNECTED_5698,SV2V_UNCONNECTED_5699,SV2V_UNCONNECTED_5700,
  SV2V_UNCONNECTED_5701,SV2V_UNCONNECTED_5702,SV2V_UNCONNECTED_5703,
  SV2V_UNCONNECTED_5704,SV2V_UNCONNECTED_5705,SV2V_UNCONNECTED_5706,
  SV2V_UNCONNECTED_5707,SV2V_UNCONNECTED_5708,SV2V_UNCONNECTED_5709,
  SV2V_UNCONNECTED_5710,SV2V_UNCONNECTED_5711,SV2V_UNCONNECTED_5712,
  SV2V_UNCONNECTED_5713,SV2V_UNCONNECTED_5714,SV2V_UNCONNECTED_5715,
  SV2V_UNCONNECTED_5716,SV2V_UNCONNECTED_5717,SV2V_UNCONNECTED_5718,
  SV2V_UNCONNECTED_5719,SV2V_UNCONNECTED_5720,SV2V_UNCONNECTED_5721,
  SV2V_UNCONNECTED_5722,SV2V_UNCONNECTED_5723,SV2V_UNCONNECTED_5724,
  SV2V_UNCONNECTED_5725,SV2V_UNCONNECTED_5726,SV2V_UNCONNECTED_5727,
  SV2V_UNCONNECTED_5728,SV2V_UNCONNECTED_5729,SV2V_UNCONNECTED_5730,
  SV2V_UNCONNECTED_5731,SV2V_UNCONNECTED_5732,SV2V_UNCONNECTED_5733,
  SV2V_UNCONNECTED_5734,SV2V_UNCONNECTED_5735,SV2V_UNCONNECTED_5736,SV2V_UNCONNECTED_5737,
  SV2V_UNCONNECTED_5738,SV2V_UNCONNECTED_5739,SV2V_UNCONNECTED_5740,
  SV2V_UNCONNECTED_5741,SV2V_UNCONNECTED_5742,SV2V_UNCONNECTED_5743,
  SV2V_UNCONNECTED_5744,SV2V_UNCONNECTED_5745,SV2V_UNCONNECTED_5746,
  SV2V_UNCONNECTED_5747,SV2V_UNCONNECTED_5748,SV2V_UNCONNECTED_5749,
  SV2V_UNCONNECTED_5750,SV2V_UNCONNECTED_5751,SV2V_UNCONNECTED_5752,
  SV2V_UNCONNECTED_5753,SV2V_UNCONNECTED_5754,SV2V_UNCONNECTED_5755,
  SV2V_UNCONNECTED_5756,SV2V_UNCONNECTED_5757,SV2V_UNCONNECTED_5758,
  SV2V_UNCONNECTED_5759,SV2V_UNCONNECTED_5760,SV2V_UNCONNECTED_5761,
  SV2V_UNCONNECTED_5762,SV2V_UNCONNECTED_5763,SV2V_UNCONNECTED_5764,
  SV2V_UNCONNECTED_5765,SV2V_UNCONNECTED_5766,SV2V_UNCONNECTED_5767,
  SV2V_UNCONNECTED_5768,SV2V_UNCONNECTED_5769,SV2V_UNCONNECTED_5770,
  SV2V_UNCONNECTED_5771,SV2V_UNCONNECTED_5772,SV2V_UNCONNECTED_5773,
  SV2V_UNCONNECTED_5774,SV2V_UNCONNECTED_5775,SV2V_UNCONNECTED_5776,SV2V_UNCONNECTED_5777,
  SV2V_UNCONNECTED_5778,SV2V_UNCONNECTED_5779,SV2V_UNCONNECTED_5780,
  SV2V_UNCONNECTED_5781,SV2V_UNCONNECTED_5782,SV2V_UNCONNECTED_5783,
  SV2V_UNCONNECTED_5784,SV2V_UNCONNECTED_5785,SV2V_UNCONNECTED_5786,
  SV2V_UNCONNECTED_5787,SV2V_UNCONNECTED_5788,SV2V_UNCONNECTED_5789,
  SV2V_UNCONNECTED_5790,SV2V_UNCONNECTED_5791,SV2V_UNCONNECTED_5792,
  SV2V_UNCONNECTED_5793,SV2V_UNCONNECTED_5794,SV2V_UNCONNECTED_5795,
  SV2V_UNCONNECTED_5796,SV2V_UNCONNECTED_5797,SV2V_UNCONNECTED_5798,
  SV2V_UNCONNECTED_5799,SV2V_UNCONNECTED_5800,SV2V_UNCONNECTED_5801,
  SV2V_UNCONNECTED_5802,SV2V_UNCONNECTED_5803,SV2V_UNCONNECTED_5804,
  SV2V_UNCONNECTED_5805,SV2V_UNCONNECTED_5806,SV2V_UNCONNECTED_5807,
  SV2V_UNCONNECTED_5808,SV2V_UNCONNECTED_5809,SV2V_UNCONNECTED_5810,
  SV2V_UNCONNECTED_5811,SV2V_UNCONNECTED_5812,SV2V_UNCONNECTED_5813,
  SV2V_UNCONNECTED_5814,SV2V_UNCONNECTED_5815,SV2V_UNCONNECTED_5816,SV2V_UNCONNECTED_5817,
  SV2V_UNCONNECTED_5818,SV2V_UNCONNECTED_5819,SV2V_UNCONNECTED_5820,
  SV2V_UNCONNECTED_5821,SV2V_UNCONNECTED_5822,SV2V_UNCONNECTED_5823,
  SV2V_UNCONNECTED_5824,SV2V_UNCONNECTED_5825,SV2V_UNCONNECTED_5826,
  SV2V_UNCONNECTED_5827,SV2V_UNCONNECTED_5828,SV2V_UNCONNECTED_5829,
  SV2V_UNCONNECTED_5830,SV2V_UNCONNECTED_5831,SV2V_UNCONNECTED_5832,
  SV2V_UNCONNECTED_5833,SV2V_UNCONNECTED_5834,SV2V_UNCONNECTED_5835,
  SV2V_UNCONNECTED_5836,SV2V_UNCONNECTED_5837,SV2V_UNCONNECTED_5838,
  SV2V_UNCONNECTED_5839,SV2V_UNCONNECTED_5840,SV2V_UNCONNECTED_5841,
  SV2V_UNCONNECTED_5842,SV2V_UNCONNECTED_5843,SV2V_UNCONNECTED_5844,
  SV2V_UNCONNECTED_5845,SV2V_UNCONNECTED_5846,SV2V_UNCONNECTED_5847,
  SV2V_UNCONNECTED_5848,SV2V_UNCONNECTED_5849,SV2V_UNCONNECTED_5850,
  SV2V_UNCONNECTED_5851,SV2V_UNCONNECTED_5852,SV2V_UNCONNECTED_5853,
  SV2V_UNCONNECTED_5854,SV2V_UNCONNECTED_5855,SV2V_UNCONNECTED_5856,SV2V_UNCONNECTED_5857,
  SV2V_UNCONNECTED_5858,SV2V_UNCONNECTED_5859,SV2V_UNCONNECTED_5860,
  SV2V_UNCONNECTED_5861,SV2V_UNCONNECTED_5862,SV2V_UNCONNECTED_5863,
  SV2V_UNCONNECTED_5864,SV2V_UNCONNECTED_5865,SV2V_UNCONNECTED_5866,
  SV2V_UNCONNECTED_5867,SV2V_UNCONNECTED_5868,SV2V_UNCONNECTED_5869,
  SV2V_UNCONNECTED_5870,SV2V_UNCONNECTED_5871,SV2V_UNCONNECTED_5872,
  SV2V_UNCONNECTED_5873,SV2V_UNCONNECTED_5874,SV2V_UNCONNECTED_5875,
  SV2V_UNCONNECTED_5876,SV2V_UNCONNECTED_5877,SV2V_UNCONNECTED_5878,
  SV2V_UNCONNECTED_5879,SV2V_UNCONNECTED_5880,SV2V_UNCONNECTED_5881,
  SV2V_UNCONNECTED_5882,SV2V_UNCONNECTED_5883,SV2V_UNCONNECTED_5884,
  SV2V_UNCONNECTED_5885,SV2V_UNCONNECTED_5886,SV2V_UNCONNECTED_5887,
  SV2V_UNCONNECTED_5888,SV2V_UNCONNECTED_5889,SV2V_UNCONNECTED_5890,
  SV2V_UNCONNECTED_5891,SV2V_UNCONNECTED_5892,SV2V_UNCONNECTED_5893,
  SV2V_UNCONNECTED_5894,SV2V_UNCONNECTED_5895,SV2V_UNCONNECTED_5896,SV2V_UNCONNECTED_5897,
  SV2V_UNCONNECTED_5898,SV2V_UNCONNECTED_5899,SV2V_UNCONNECTED_5900,
  SV2V_UNCONNECTED_5901,SV2V_UNCONNECTED_5902,SV2V_UNCONNECTED_5903,
  SV2V_UNCONNECTED_5904,SV2V_UNCONNECTED_5905,SV2V_UNCONNECTED_5906,
  SV2V_UNCONNECTED_5907,SV2V_UNCONNECTED_5908,SV2V_UNCONNECTED_5909,
  SV2V_UNCONNECTED_5910,SV2V_UNCONNECTED_5911,SV2V_UNCONNECTED_5912,
  SV2V_UNCONNECTED_5913,SV2V_UNCONNECTED_5914,SV2V_UNCONNECTED_5915,
  SV2V_UNCONNECTED_5916,SV2V_UNCONNECTED_5917,SV2V_UNCONNECTED_5918,
  SV2V_UNCONNECTED_5919,SV2V_UNCONNECTED_5920,SV2V_UNCONNECTED_5921,
  SV2V_UNCONNECTED_5922,SV2V_UNCONNECTED_5923,SV2V_UNCONNECTED_5924,
  SV2V_UNCONNECTED_5925,SV2V_UNCONNECTED_5926,SV2V_UNCONNECTED_5927,
  SV2V_UNCONNECTED_5928,SV2V_UNCONNECTED_5929,SV2V_UNCONNECTED_5930,
  SV2V_UNCONNECTED_5931,SV2V_UNCONNECTED_5932,SV2V_UNCONNECTED_5933,
  SV2V_UNCONNECTED_5934,SV2V_UNCONNECTED_5935,SV2V_UNCONNECTED_5936,SV2V_UNCONNECTED_5937,
  SV2V_UNCONNECTED_5938,SV2V_UNCONNECTED_5939,SV2V_UNCONNECTED_5940,
  SV2V_UNCONNECTED_5941,SV2V_UNCONNECTED_5942,SV2V_UNCONNECTED_5943,
  SV2V_UNCONNECTED_5944,SV2V_UNCONNECTED_5945,SV2V_UNCONNECTED_5946,
  SV2V_UNCONNECTED_5947,SV2V_UNCONNECTED_5948,SV2V_UNCONNECTED_5949,
  SV2V_UNCONNECTED_5950,SV2V_UNCONNECTED_5951,SV2V_UNCONNECTED_5952,
  SV2V_UNCONNECTED_5953,SV2V_UNCONNECTED_5954,SV2V_UNCONNECTED_5955,
  SV2V_UNCONNECTED_5956,SV2V_UNCONNECTED_5957,SV2V_UNCONNECTED_5958,
  SV2V_UNCONNECTED_5959,SV2V_UNCONNECTED_5960,SV2V_UNCONNECTED_5961,
  SV2V_UNCONNECTED_5962,SV2V_UNCONNECTED_5963,SV2V_UNCONNECTED_5964,
  SV2V_UNCONNECTED_5965,SV2V_UNCONNECTED_5966,SV2V_UNCONNECTED_5967,
  SV2V_UNCONNECTED_5968,SV2V_UNCONNECTED_5969,SV2V_UNCONNECTED_5970,
  SV2V_UNCONNECTED_5971,SV2V_UNCONNECTED_5972,SV2V_UNCONNECTED_5973,
  SV2V_UNCONNECTED_5974,SV2V_UNCONNECTED_5975,SV2V_UNCONNECTED_5976,SV2V_UNCONNECTED_5977,
  SV2V_UNCONNECTED_5978,SV2V_UNCONNECTED_5979,SV2V_UNCONNECTED_5980,
  SV2V_UNCONNECTED_5981,SV2V_UNCONNECTED_5982,SV2V_UNCONNECTED_5983,
  SV2V_UNCONNECTED_5984,SV2V_UNCONNECTED_5985,SV2V_UNCONNECTED_5986,
  SV2V_UNCONNECTED_5987,SV2V_UNCONNECTED_5988,SV2V_UNCONNECTED_5989,
  SV2V_UNCONNECTED_5990,SV2V_UNCONNECTED_5991,SV2V_UNCONNECTED_5992,
  SV2V_UNCONNECTED_5993,SV2V_UNCONNECTED_5994,SV2V_UNCONNECTED_5995,
  SV2V_UNCONNECTED_5996,SV2V_UNCONNECTED_5997,SV2V_UNCONNECTED_5998,
  SV2V_UNCONNECTED_5999,SV2V_UNCONNECTED_6000,SV2V_UNCONNECTED_6001,
  SV2V_UNCONNECTED_6002,SV2V_UNCONNECTED_6003,SV2V_UNCONNECTED_6004,
  SV2V_UNCONNECTED_6005,SV2V_UNCONNECTED_6006,SV2V_UNCONNECTED_6007,
  SV2V_UNCONNECTED_6008,SV2V_UNCONNECTED_6009,SV2V_UNCONNECTED_6010,
  SV2V_UNCONNECTED_6011,SV2V_UNCONNECTED_6012,SV2V_UNCONNECTED_6013,
  SV2V_UNCONNECTED_6014,SV2V_UNCONNECTED_6015,SV2V_UNCONNECTED_6016,SV2V_UNCONNECTED_6017,
  SV2V_UNCONNECTED_6018,SV2V_UNCONNECTED_6019,SV2V_UNCONNECTED_6020,
  SV2V_UNCONNECTED_6021,SV2V_UNCONNECTED_6022,SV2V_UNCONNECTED_6023,
  SV2V_UNCONNECTED_6024,SV2V_UNCONNECTED_6025,SV2V_UNCONNECTED_6026,
  SV2V_UNCONNECTED_6027,SV2V_UNCONNECTED_6028,SV2V_UNCONNECTED_6029,
  SV2V_UNCONNECTED_6030,SV2V_UNCONNECTED_6031,SV2V_UNCONNECTED_6032,
  SV2V_UNCONNECTED_6033,SV2V_UNCONNECTED_6034,SV2V_UNCONNECTED_6035,
  SV2V_UNCONNECTED_6036,SV2V_UNCONNECTED_6037,SV2V_UNCONNECTED_6038,
  SV2V_UNCONNECTED_6039,SV2V_UNCONNECTED_6040,SV2V_UNCONNECTED_6041,
  SV2V_UNCONNECTED_6042,SV2V_UNCONNECTED_6043,SV2V_UNCONNECTED_6044,
  SV2V_UNCONNECTED_6045,SV2V_UNCONNECTED_6046,SV2V_UNCONNECTED_6047,
  SV2V_UNCONNECTED_6048,SV2V_UNCONNECTED_6049,SV2V_UNCONNECTED_6050,
  SV2V_UNCONNECTED_6051,SV2V_UNCONNECTED_6052,SV2V_UNCONNECTED_6053,
  SV2V_UNCONNECTED_6054,SV2V_UNCONNECTED_6055,SV2V_UNCONNECTED_6056,SV2V_UNCONNECTED_6057,
  SV2V_UNCONNECTED_6058,SV2V_UNCONNECTED_6059,SV2V_UNCONNECTED_6060,
  SV2V_UNCONNECTED_6061,SV2V_UNCONNECTED_6062,SV2V_UNCONNECTED_6063,
  SV2V_UNCONNECTED_6064,SV2V_UNCONNECTED_6065,SV2V_UNCONNECTED_6066,
  SV2V_UNCONNECTED_6067,SV2V_UNCONNECTED_6068,SV2V_UNCONNECTED_6069,
  SV2V_UNCONNECTED_6070,SV2V_UNCONNECTED_6071,SV2V_UNCONNECTED_6072,
  SV2V_UNCONNECTED_6073,SV2V_UNCONNECTED_6074,SV2V_UNCONNECTED_6075,
  SV2V_UNCONNECTED_6076,SV2V_UNCONNECTED_6077,SV2V_UNCONNECTED_6078,
  SV2V_UNCONNECTED_6079,SV2V_UNCONNECTED_6080,SV2V_UNCONNECTED_6081,
  SV2V_UNCONNECTED_6082,SV2V_UNCONNECTED_6083,SV2V_UNCONNECTED_6084,
  SV2V_UNCONNECTED_6085,SV2V_UNCONNECTED_6086,SV2V_UNCONNECTED_6087,
  SV2V_UNCONNECTED_6088,SV2V_UNCONNECTED_6089,SV2V_UNCONNECTED_6090,
  SV2V_UNCONNECTED_6091,SV2V_UNCONNECTED_6092,SV2V_UNCONNECTED_6093,
  SV2V_UNCONNECTED_6094,SV2V_UNCONNECTED_6095,SV2V_UNCONNECTED_6096,SV2V_UNCONNECTED_6097,
  SV2V_UNCONNECTED_6098,SV2V_UNCONNECTED_6099,SV2V_UNCONNECTED_6100,
  SV2V_UNCONNECTED_6101,SV2V_UNCONNECTED_6102,SV2V_UNCONNECTED_6103,
  SV2V_UNCONNECTED_6104,SV2V_UNCONNECTED_6105,SV2V_UNCONNECTED_6106,
  SV2V_UNCONNECTED_6107,SV2V_UNCONNECTED_6108,SV2V_UNCONNECTED_6109,
  SV2V_UNCONNECTED_6110,SV2V_UNCONNECTED_6111,SV2V_UNCONNECTED_6112,
  SV2V_UNCONNECTED_6113,SV2V_UNCONNECTED_6114,SV2V_UNCONNECTED_6115,
  SV2V_UNCONNECTED_6116,SV2V_UNCONNECTED_6117,SV2V_UNCONNECTED_6118,
  SV2V_UNCONNECTED_6119,SV2V_UNCONNECTED_6120,SV2V_UNCONNECTED_6121,
  SV2V_UNCONNECTED_6122,SV2V_UNCONNECTED_6123,SV2V_UNCONNECTED_6124,
  SV2V_UNCONNECTED_6125,SV2V_UNCONNECTED_6126,SV2V_UNCONNECTED_6127,
  SV2V_UNCONNECTED_6128,SV2V_UNCONNECTED_6129,SV2V_UNCONNECTED_6130,
  SV2V_UNCONNECTED_6131,SV2V_UNCONNECTED_6132,SV2V_UNCONNECTED_6133,
  SV2V_UNCONNECTED_6134,SV2V_UNCONNECTED_6135,SV2V_UNCONNECTED_6136,SV2V_UNCONNECTED_6137,
  SV2V_UNCONNECTED_6138,SV2V_UNCONNECTED_6139,SV2V_UNCONNECTED_6140,
  SV2V_UNCONNECTED_6141,SV2V_UNCONNECTED_6142,SV2V_UNCONNECTED_6143,
  SV2V_UNCONNECTED_6144,SV2V_UNCONNECTED_6145,SV2V_UNCONNECTED_6146,
  SV2V_UNCONNECTED_6147,SV2V_UNCONNECTED_6148,SV2V_UNCONNECTED_6149,
  SV2V_UNCONNECTED_6150,SV2V_UNCONNECTED_6151,SV2V_UNCONNECTED_6152,
  SV2V_UNCONNECTED_6153,SV2V_UNCONNECTED_6154,SV2V_UNCONNECTED_6155,
  SV2V_UNCONNECTED_6156,SV2V_UNCONNECTED_6157,SV2V_UNCONNECTED_6158,
  SV2V_UNCONNECTED_6159,SV2V_UNCONNECTED_6160,SV2V_UNCONNECTED_6161,
  SV2V_UNCONNECTED_6162,SV2V_UNCONNECTED_6163,SV2V_UNCONNECTED_6164,
  SV2V_UNCONNECTED_6165,SV2V_UNCONNECTED_6166,SV2V_UNCONNECTED_6167,
  SV2V_UNCONNECTED_6168,SV2V_UNCONNECTED_6169,SV2V_UNCONNECTED_6170,
  SV2V_UNCONNECTED_6171,SV2V_UNCONNECTED_6172,SV2V_UNCONNECTED_6173,
  SV2V_UNCONNECTED_6174,SV2V_UNCONNECTED_6175,SV2V_UNCONNECTED_6176,SV2V_UNCONNECTED_6177,
  SV2V_UNCONNECTED_6178,SV2V_UNCONNECTED_6179,SV2V_UNCONNECTED_6180,
  SV2V_UNCONNECTED_6181,SV2V_UNCONNECTED_6182,SV2V_UNCONNECTED_6183,
  SV2V_UNCONNECTED_6184,SV2V_UNCONNECTED_6185,SV2V_UNCONNECTED_6186,
  SV2V_UNCONNECTED_6187,SV2V_UNCONNECTED_6188,SV2V_UNCONNECTED_6189,
  SV2V_UNCONNECTED_6190,SV2V_UNCONNECTED_6191,SV2V_UNCONNECTED_6192,
  SV2V_UNCONNECTED_6193,SV2V_UNCONNECTED_6194,SV2V_UNCONNECTED_6195,
  SV2V_UNCONNECTED_6196,SV2V_UNCONNECTED_6197,SV2V_UNCONNECTED_6198,
  SV2V_UNCONNECTED_6199,SV2V_UNCONNECTED_6200,SV2V_UNCONNECTED_6201,
  SV2V_UNCONNECTED_6202,SV2V_UNCONNECTED_6203,SV2V_UNCONNECTED_6204,
  SV2V_UNCONNECTED_6205,SV2V_UNCONNECTED_6206,SV2V_UNCONNECTED_6207,
  SV2V_UNCONNECTED_6208,SV2V_UNCONNECTED_6209,SV2V_UNCONNECTED_6210,
  SV2V_UNCONNECTED_6211,SV2V_UNCONNECTED_6212,SV2V_UNCONNECTED_6213,
  SV2V_UNCONNECTED_6214,SV2V_UNCONNECTED_6215,SV2V_UNCONNECTED_6216,SV2V_UNCONNECTED_6217,
  SV2V_UNCONNECTED_6218,SV2V_UNCONNECTED_6219,SV2V_UNCONNECTED_6220,
  SV2V_UNCONNECTED_6221,SV2V_UNCONNECTED_6222,SV2V_UNCONNECTED_6223,
  SV2V_UNCONNECTED_6224,SV2V_UNCONNECTED_6225,SV2V_UNCONNECTED_6226,
  SV2V_UNCONNECTED_6227,SV2V_UNCONNECTED_6228,SV2V_UNCONNECTED_6229,
  SV2V_UNCONNECTED_6230,SV2V_UNCONNECTED_6231,SV2V_UNCONNECTED_6232,
  SV2V_UNCONNECTED_6233,SV2V_UNCONNECTED_6234,SV2V_UNCONNECTED_6235,
  SV2V_UNCONNECTED_6236,SV2V_UNCONNECTED_6237,SV2V_UNCONNECTED_6238,
  SV2V_UNCONNECTED_6239,SV2V_UNCONNECTED_6240,SV2V_UNCONNECTED_6241,
  SV2V_UNCONNECTED_6242,SV2V_UNCONNECTED_6243,SV2V_UNCONNECTED_6244,
  SV2V_UNCONNECTED_6245,SV2V_UNCONNECTED_6246,SV2V_UNCONNECTED_6247,
  SV2V_UNCONNECTED_6248,SV2V_UNCONNECTED_6249,SV2V_UNCONNECTED_6250,
  SV2V_UNCONNECTED_6251,SV2V_UNCONNECTED_6252,SV2V_UNCONNECTED_6253,
  SV2V_UNCONNECTED_6254,SV2V_UNCONNECTED_6255,SV2V_UNCONNECTED_6256,SV2V_UNCONNECTED_6257,
  SV2V_UNCONNECTED_6258,SV2V_UNCONNECTED_6259,SV2V_UNCONNECTED_6260,
  SV2V_UNCONNECTED_6261,SV2V_UNCONNECTED_6262,SV2V_UNCONNECTED_6263,
  SV2V_UNCONNECTED_6264,SV2V_UNCONNECTED_6265,SV2V_UNCONNECTED_6266,
  SV2V_UNCONNECTED_6267,SV2V_UNCONNECTED_6268,SV2V_UNCONNECTED_6269,
  SV2V_UNCONNECTED_6270,SV2V_UNCONNECTED_6271,SV2V_UNCONNECTED_6272,
  SV2V_UNCONNECTED_6273,SV2V_UNCONNECTED_6274,SV2V_UNCONNECTED_6275,
  SV2V_UNCONNECTED_6276,SV2V_UNCONNECTED_6277,SV2V_UNCONNECTED_6278,
  SV2V_UNCONNECTED_6279,SV2V_UNCONNECTED_6280,SV2V_UNCONNECTED_6281,
  SV2V_UNCONNECTED_6282,SV2V_UNCONNECTED_6283,SV2V_UNCONNECTED_6284,
  SV2V_UNCONNECTED_6285,SV2V_UNCONNECTED_6286,SV2V_UNCONNECTED_6287,
  SV2V_UNCONNECTED_6288,SV2V_UNCONNECTED_6289,SV2V_UNCONNECTED_6290,
  SV2V_UNCONNECTED_6291,SV2V_UNCONNECTED_6292,SV2V_UNCONNECTED_6293,
  SV2V_UNCONNECTED_6294,SV2V_UNCONNECTED_6295,SV2V_UNCONNECTED_6296,SV2V_UNCONNECTED_6297,
  SV2V_UNCONNECTED_6298,SV2V_UNCONNECTED_6299,SV2V_UNCONNECTED_6300,
  SV2V_UNCONNECTED_6301,SV2V_UNCONNECTED_6302,SV2V_UNCONNECTED_6303,
  SV2V_UNCONNECTED_6304,SV2V_UNCONNECTED_6305,SV2V_UNCONNECTED_6306,
  SV2V_UNCONNECTED_6307,SV2V_UNCONNECTED_6308,SV2V_UNCONNECTED_6309,
  SV2V_UNCONNECTED_6310,SV2V_UNCONNECTED_6311,SV2V_UNCONNECTED_6312,
  SV2V_UNCONNECTED_6313,SV2V_UNCONNECTED_6314,SV2V_UNCONNECTED_6315,
  SV2V_UNCONNECTED_6316,SV2V_UNCONNECTED_6317,SV2V_UNCONNECTED_6318,
  SV2V_UNCONNECTED_6319,SV2V_UNCONNECTED_6320,SV2V_UNCONNECTED_6321,
  SV2V_UNCONNECTED_6322,SV2V_UNCONNECTED_6323,SV2V_UNCONNECTED_6324,
  SV2V_UNCONNECTED_6325,SV2V_UNCONNECTED_6326,SV2V_UNCONNECTED_6327,
  SV2V_UNCONNECTED_6328,SV2V_UNCONNECTED_6329,SV2V_UNCONNECTED_6330,
  SV2V_UNCONNECTED_6331,SV2V_UNCONNECTED_6332,SV2V_UNCONNECTED_6333,
  SV2V_UNCONNECTED_6334,SV2V_UNCONNECTED_6335,SV2V_UNCONNECTED_6336,SV2V_UNCONNECTED_6337,
  SV2V_UNCONNECTED_6338,SV2V_UNCONNECTED_6339,SV2V_UNCONNECTED_6340,
  SV2V_UNCONNECTED_6341,SV2V_UNCONNECTED_6342,SV2V_UNCONNECTED_6343,
  SV2V_UNCONNECTED_6344,SV2V_UNCONNECTED_6345,SV2V_UNCONNECTED_6346,
  SV2V_UNCONNECTED_6347,SV2V_UNCONNECTED_6348,SV2V_UNCONNECTED_6349,
  SV2V_UNCONNECTED_6350,SV2V_UNCONNECTED_6351,SV2V_UNCONNECTED_6352,
  SV2V_UNCONNECTED_6353,SV2V_UNCONNECTED_6354,SV2V_UNCONNECTED_6355,
  SV2V_UNCONNECTED_6356,SV2V_UNCONNECTED_6357,SV2V_UNCONNECTED_6358,
  SV2V_UNCONNECTED_6359,SV2V_UNCONNECTED_6360,SV2V_UNCONNECTED_6361,
  SV2V_UNCONNECTED_6362,SV2V_UNCONNECTED_6363,SV2V_UNCONNECTED_6364,
  SV2V_UNCONNECTED_6365,SV2V_UNCONNECTED_6366,SV2V_UNCONNECTED_6367,
  SV2V_UNCONNECTED_6368,SV2V_UNCONNECTED_6369,SV2V_UNCONNECTED_6370,
  SV2V_UNCONNECTED_6371,SV2V_UNCONNECTED_6372,SV2V_UNCONNECTED_6373,
  SV2V_UNCONNECTED_6374,SV2V_UNCONNECTED_6375,SV2V_UNCONNECTED_6376,SV2V_UNCONNECTED_6377,
  SV2V_UNCONNECTED_6378,SV2V_UNCONNECTED_6379,SV2V_UNCONNECTED_6380,
  SV2V_UNCONNECTED_6381,SV2V_UNCONNECTED_6382,SV2V_UNCONNECTED_6383,
  SV2V_UNCONNECTED_6384,SV2V_UNCONNECTED_6385,SV2V_UNCONNECTED_6386,
  SV2V_UNCONNECTED_6387,SV2V_UNCONNECTED_6388,SV2V_UNCONNECTED_6389,
  SV2V_UNCONNECTED_6390,SV2V_UNCONNECTED_6391,SV2V_UNCONNECTED_6392,
  SV2V_UNCONNECTED_6393,SV2V_UNCONNECTED_6394,SV2V_UNCONNECTED_6395,
  SV2V_UNCONNECTED_6396,SV2V_UNCONNECTED_6397,SV2V_UNCONNECTED_6398,
  SV2V_UNCONNECTED_6399,SV2V_UNCONNECTED_6400,SV2V_UNCONNECTED_6401,
  SV2V_UNCONNECTED_6402,SV2V_UNCONNECTED_6403,SV2V_UNCONNECTED_6404,
  SV2V_UNCONNECTED_6405,SV2V_UNCONNECTED_6406,SV2V_UNCONNECTED_6407,
  SV2V_UNCONNECTED_6408,SV2V_UNCONNECTED_6409,SV2V_UNCONNECTED_6410,
  SV2V_UNCONNECTED_6411,SV2V_UNCONNECTED_6412,SV2V_UNCONNECTED_6413,
  SV2V_UNCONNECTED_6414,SV2V_UNCONNECTED_6415,SV2V_UNCONNECTED_6416,SV2V_UNCONNECTED_6417,
  SV2V_UNCONNECTED_6418,SV2V_UNCONNECTED_6419,SV2V_UNCONNECTED_6420,
  SV2V_UNCONNECTED_6421,SV2V_UNCONNECTED_6422,SV2V_UNCONNECTED_6423,
  SV2V_UNCONNECTED_6424,SV2V_UNCONNECTED_6425,SV2V_UNCONNECTED_6426,
  SV2V_UNCONNECTED_6427,SV2V_UNCONNECTED_6428,SV2V_UNCONNECTED_6429,
  SV2V_UNCONNECTED_6430,SV2V_UNCONNECTED_6431,SV2V_UNCONNECTED_6432,
  SV2V_UNCONNECTED_6433,SV2V_UNCONNECTED_6434,SV2V_UNCONNECTED_6435,
  SV2V_UNCONNECTED_6436,SV2V_UNCONNECTED_6437,SV2V_UNCONNECTED_6438,
  SV2V_UNCONNECTED_6439,SV2V_UNCONNECTED_6440,SV2V_UNCONNECTED_6441,
  SV2V_UNCONNECTED_6442,SV2V_UNCONNECTED_6443,SV2V_UNCONNECTED_6444,
  SV2V_UNCONNECTED_6445,SV2V_UNCONNECTED_6446,SV2V_UNCONNECTED_6447,
  SV2V_UNCONNECTED_6448,SV2V_UNCONNECTED_6449,SV2V_UNCONNECTED_6450,
  SV2V_UNCONNECTED_6451,SV2V_UNCONNECTED_6452,SV2V_UNCONNECTED_6453,
  SV2V_UNCONNECTED_6454,SV2V_UNCONNECTED_6455,SV2V_UNCONNECTED_6456,SV2V_UNCONNECTED_6457,
  SV2V_UNCONNECTED_6458,SV2V_UNCONNECTED_6459,SV2V_UNCONNECTED_6460,
  SV2V_UNCONNECTED_6461,SV2V_UNCONNECTED_6462,SV2V_UNCONNECTED_6463,
  SV2V_UNCONNECTED_6464,SV2V_UNCONNECTED_6465,SV2V_UNCONNECTED_6466,
  SV2V_UNCONNECTED_6467,SV2V_UNCONNECTED_6468,SV2V_UNCONNECTED_6469,
  SV2V_UNCONNECTED_6470,SV2V_UNCONNECTED_6471,SV2V_UNCONNECTED_6472,
  SV2V_UNCONNECTED_6473,SV2V_UNCONNECTED_6474,SV2V_UNCONNECTED_6475,
  SV2V_UNCONNECTED_6476,SV2V_UNCONNECTED_6477,SV2V_UNCONNECTED_6478,
  SV2V_UNCONNECTED_6479,SV2V_UNCONNECTED_6480,SV2V_UNCONNECTED_6481,
  SV2V_UNCONNECTED_6482,SV2V_UNCONNECTED_6483,SV2V_UNCONNECTED_6484,
  SV2V_UNCONNECTED_6485,SV2V_UNCONNECTED_6486,SV2V_UNCONNECTED_6487,
  SV2V_UNCONNECTED_6488,SV2V_UNCONNECTED_6489,SV2V_UNCONNECTED_6490,
  SV2V_UNCONNECTED_6491,SV2V_UNCONNECTED_6492,SV2V_UNCONNECTED_6493,
  SV2V_UNCONNECTED_6494,SV2V_UNCONNECTED_6495,SV2V_UNCONNECTED_6496,SV2V_UNCONNECTED_6497,
  SV2V_UNCONNECTED_6498,SV2V_UNCONNECTED_6499,SV2V_UNCONNECTED_6500,
  SV2V_UNCONNECTED_6501,SV2V_UNCONNECTED_6502,SV2V_UNCONNECTED_6503,
  SV2V_UNCONNECTED_6504,SV2V_UNCONNECTED_6505,SV2V_UNCONNECTED_6506,
  SV2V_UNCONNECTED_6507,SV2V_UNCONNECTED_6508,SV2V_UNCONNECTED_6509,
  SV2V_UNCONNECTED_6510,SV2V_UNCONNECTED_6511,SV2V_UNCONNECTED_6512,
  SV2V_UNCONNECTED_6513,SV2V_UNCONNECTED_6514,SV2V_UNCONNECTED_6515,
  SV2V_UNCONNECTED_6516,SV2V_UNCONNECTED_6517,SV2V_UNCONNECTED_6518,
  SV2V_UNCONNECTED_6519,SV2V_UNCONNECTED_6520,SV2V_UNCONNECTED_6521,
  SV2V_UNCONNECTED_6522,SV2V_UNCONNECTED_6523,SV2V_UNCONNECTED_6524,
  SV2V_UNCONNECTED_6525,SV2V_UNCONNECTED_6526,SV2V_UNCONNECTED_6527,
  SV2V_UNCONNECTED_6528,SV2V_UNCONNECTED_6529,SV2V_UNCONNECTED_6530,
  SV2V_UNCONNECTED_6531,SV2V_UNCONNECTED_6532,SV2V_UNCONNECTED_6533,
  SV2V_UNCONNECTED_6534,SV2V_UNCONNECTED_6535,SV2V_UNCONNECTED_6536,SV2V_UNCONNECTED_6537,
  SV2V_UNCONNECTED_6538,SV2V_UNCONNECTED_6539,SV2V_UNCONNECTED_6540,
  SV2V_UNCONNECTED_6541,SV2V_UNCONNECTED_6542,SV2V_UNCONNECTED_6543,
  SV2V_UNCONNECTED_6544,SV2V_UNCONNECTED_6545,SV2V_UNCONNECTED_6546,
  SV2V_UNCONNECTED_6547,SV2V_UNCONNECTED_6548,SV2V_UNCONNECTED_6549,
  SV2V_UNCONNECTED_6550,SV2V_UNCONNECTED_6551,SV2V_UNCONNECTED_6552,
  SV2V_UNCONNECTED_6553,SV2V_UNCONNECTED_6554,SV2V_UNCONNECTED_6555,
  SV2V_UNCONNECTED_6556,SV2V_UNCONNECTED_6557,SV2V_UNCONNECTED_6558,
  SV2V_UNCONNECTED_6559,SV2V_UNCONNECTED_6560,SV2V_UNCONNECTED_6561,
  SV2V_UNCONNECTED_6562,SV2V_UNCONNECTED_6563,SV2V_UNCONNECTED_6564,
  SV2V_UNCONNECTED_6565,SV2V_UNCONNECTED_6566,SV2V_UNCONNECTED_6567,
  SV2V_UNCONNECTED_6568,SV2V_UNCONNECTED_6569,SV2V_UNCONNECTED_6570,
  SV2V_UNCONNECTED_6571,SV2V_UNCONNECTED_6572,SV2V_UNCONNECTED_6573,
  SV2V_UNCONNECTED_6574,SV2V_UNCONNECTED_6575,SV2V_UNCONNECTED_6576,SV2V_UNCONNECTED_6577,
  SV2V_UNCONNECTED_6578,SV2V_UNCONNECTED_6579,SV2V_UNCONNECTED_6580,
  SV2V_UNCONNECTED_6581,SV2V_UNCONNECTED_6582,SV2V_UNCONNECTED_6583,
  SV2V_UNCONNECTED_6584,SV2V_UNCONNECTED_6585,SV2V_UNCONNECTED_6586,
  SV2V_UNCONNECTED_6587,SV2V_UNCONNECTED_6588,SV2V_UNCONNECTED_6589,
  SV2V_UNCONNECTED_6590,SV2V_UNCONNECTED_6591,SV2V_UNCONNECTED_6592,
  SV2V_UNCONNECTED_6593,SV2V_UNCONNECTED_6594,SV2V_UNCONNECTED_6595,
  SV2V_UNCONNECTED_6596,SV2V_UNCONNECTED_6597,SV2V_UNCONNECTED_6598,
  SV2V_UNCONNECTED_6599,SV2V_UNCONNECTED_6600,SV2V_UNCONNECTED_6601,
  SV2V_UNCONNECTED_6602,SV2V_UNCONNECTED_6603,SV2V_UNCONNECTED_6604,
  SV2V_UNCONNECTED_6605,SV2V_UNCONNECTED_6606,SV2V_UNCONNECTED_6607,
  SV2V_UNCONNECTED_6608,SV2V_UNCONNECTED_6609,SV2V_UNCONNECTED_6610,
  SV2V_UNCONNECTED_6611,SV2V_UNCONNECTED_6612,SV2V_UNCONNECTED_6613,
  SV2V_UNCONNECTED_6614,SV2V_UNCONNECTED_6615,SV2V_UNCONNECTED_6616,SV2V_UNCONNECTED_6617,
  SV2V_UNCONNECTED_6618,SV2V_UNCONNECTED_6619,SV2V_UNCONNECTED_6620,
  SV2V_UNCONNECTED_6621,SV2V_UNCONNECTED_6622,SV2V_UNCONNECTED_6623,
  SV2V_UNCONNECTED_6624,SV2V_UNCONNECTED_6625,SV2V_UNCONNECTED_6626,
  SV2V_UNCONNECTED_6627,SV2V_UNCONNECTED_6628,SV2V_UNCONNECTED_6629,
  SV2V_UNCONNECTED_6630,SV2V_UNCONNECTED_6631,SV2V_UNCONNECTED_6632,
  SV2V_UNCONNECTED_6633,SV2V_UNCONNECTED_6634,SV2V_UNCONNECTED_6635,
  SV2V_UNCONNECTED_6636,SV2V_UNCONNECTED_6637,SV2V_UNCONNECTED_6638,
  SV2V_UNCONNECTED_6639,SV2V_UNCONNECTED_6640,SV2V_UNCONNECTED_6641,
  SV2V_UNCONNECTED_6642,SV2V_UNCONNECTED_6643,SV2V_UNCONNECTED_6644,
  SV2V_UNCONNECTED_6645,SV2V_UNCONNECTED_6646,SV2V_UNCONNECTED_6647,
  SV2V_UNCONNECTED_6648,SV2V_UNCONNECTED_6649,SV2V_UNCONNECTED_6650,
  SV2V_UNCONNECTED_6651,SV2V_UNCONNECTED_6652,SV2V_UNCONNECTED_6653,
  SV2V_UNCONNECTED_6654,SV2V_UNCONNECTED_6655,SV2V_UNCONNECTED_6656,SV2V_UNCONNECTED_6657,
  SV2V_UNCONNECTED_6658,SV2V_UNCONNECTED_6659,SV2V_UNCONNECTED_6660,
  SV2V_UNCONNECTED_6661,SV2V_UNCONNECTED_6662,SV2V_UNCONNECTED_6663,
  SV2V_UNCONNECTED_6664,SV2V_UNCONNECTED_6665,SV2V_UNCONNECTED_6666,
  SV2V_UNCONNECTED_6667,SV2V_UNCONNECTED_6668,SV2V_UNCONNECTED_6669,
  SV2V_UNCONNECTED_6670,SV2V_UNCONNECTED_6671,SV2V_UNCONNECTED_6672,
  SV2V_UNCONNECTED_6673,SV2V_UNCONNECTED_6674,SV2V_UNCONNECTED_6675,
  SV2V_UNCONNECTED_6676,SV2V_UNCONNECTED_6677,SV2V_UNCONNECTED_6678,
  SV2V_UNCONNECTED_6679,SV2V_UNCONNECTED_6680,SV2V_UNCONNECTED_6681,
  SV2V_UNCONNECTED_6682,SV2V_UNCONNECTED_6683,SV2V_UNCONNECTED_6684,
  SV2V_UNCONNECTED_6685,SV2V_UNCONNECTED_6686,SV2V_UNCONNECTED_6687,
  SV2V_UNCONNECTED_6688,SV2V_UNCONNECTED_6689,SV2V_UNCONNECTED_6690,
  SV2V_UNCONNECTED_6691,SV2V_UNCONNECTED_6692,SV2V_UNCONNECTED_6693,
  SV2V_UNCONNECTED_6694,SV2V_UNCONNECTED_6695,SV2V_UNCONNECTED_6696,SV2V_UNCONNECTED_6697,
  SV2V_UNCONNECTED_6698,SV2V_UNCONNECTED_6699,SV2V_UNCONNECTED_6700,
  SV2V_UNCONNECTED_6701,SV2V_UNCONNECTED_6702,SV2V_UNCONNECTED_6703,
  SV2V_UNCONNECTED_6704,SV2V_UNCONNECTED_6705,SV2V_UNCONNECTED_6706,
  SV2V_UNCONNECTED_6707,SV2V_UNCONNECTED_6708,SV2V_UNCONNECTED_6709,
  SV2V_UNCONNECTED_6710,SV2V_UNCONNECTED_6711,SV2V_UNCONNECTED_6712,
  SV2V_UNCONNECTED_6713,SV2V_UNCONNECTED_6714,SV2V_UNCONNECTED_6715,
  SV2V_UNCONNECTED_6716,SV2V_UNCONNECTED_6717,SV2V_UNCONNECTED_6718,
  SV2V_UNCONNECTED_6719,SV2V_UNCONNECTED_6720,SV2V_UNCONNECTED_6721,
  SV2V_UNCONNECTED_6722,SV2V_UNCONNECTED_6723,SV2V_UNCONNECTED_6724,
  SV2V_UNCONNECTED_6725,SV2V_UNCONNECTED_6726,SV2V_UNCONNECTED_6727,
  SV2V_UNCONNECTED_6728,SV2V_UNCONNECTED_6729,SV2V_UNCONNECTED_6730,
  SV2V_UNCONNECTED_6731,SV2V_UNCONNECTED_6732,SV2V_UNCONNECTED_6733,
  SV2V_UNCONNECTED_6734,SV2V_UNCONNECTED_6735,SV2V_UNCONNECTED_6736,SV2V_UNCONNECTED_6737,
  SV2V_UNCONNECTED_6738,SV2V_UNCONNECTED_6739,SV2V_UNCONNECTED_6740,
  SV2V_UNCONNECTED_6741,SV2V_UNCONNECTED_6742,SV2V_UNCONNECTED_6743,
  SV2V_UNCONNECTED_6744,SV2V_UNCONNECTED_6745,SV2V_UNCONNECTED_6746,
  SV2V_UNCONNECTED_6747,SV2V_UNCONNECTED_6748,SV2V_UNCONNECTED_6749,
  SV2V_UNCONNECTED_6750,SV2V_UNCONNECTED_6751,SV2V_UNCONNECTED_6752,
  SV2V_UNCONNECTED_6753,SV2V_UNCONNECTED_6754,SV2V_UNCONNECTED_6755,
  SV2V_UNCONNECTED_6756,SV2V_UNCONNECTED_6757,SV2V_UNCONNECTED_6758,
  SV2V_UNCONNECTED_6759,SV2V_UNCONNECTED_6760,SV2V_UNCONNECTED_6761,
  SV2V_UNCONNECTED_6762,SV2V_UNCONNECTED_6763,SV2V_UNCONNECTED_6764,
  SV2V_UNCONNECTED_6765,SV2V_UNCONNECTED_6766,SV2V_UNCONNECTED_6767,
  SV2V_UNCONNECTED_6768,SV2V_UNCONNECTED_6769,SV2V_UNCONNECTED_6770,
  SV2V_UNCONNECTED_6771,SV2V_UNCONNECTED_6772,SV2V_UNCONNECTED_6773,
  SV2V_UNCONNECTED_6774,SV2V_UNCONNECTED_6775,SV2V_UNCONNECTED_6776,SV2V_UNCONNECTED_6777,
  SV2V_UNCONNECTED_6778,SV2V_UNCONNECTED_6779,SV2V_UNCONNECTED_6780,
  SV2V_UNCONNECTED_6781,SV2V_UNCONNECTED_6782,SV2V_UNCONNECTED_6783,
  SV2V_UNCONNECTED_6784,SV2V_UNCONNECTED_6785,SV2V_UNCONNECTED_6786,
  SV2V_UNCONNECTED_6787,SV2V_UNCONNECTED_6788,SV2V_UNCONNECTED_6789,
  SV2V_UNCONNECTED_6790,SV2V_UNCONNECTED_6791,SV2V_UNCONNECTED_6792,
  SV2V_UNCONNECTED_6793,SV2V_UNCONNECTED_6794,SV2V_UNCONNECTED_6795,
  SV2V_UNCONNECTED_6796,SV2V_UNCONNECTED_6797,SV2V_UNCONNECTED_6798,
  SV2V_UNCONNECTED_6799,SV2V_UNCONNECTED_6800,SV2V_UNCONNECTED_6801,
  SV2V_UNCONNECTED_6802,SV2V_UNCONNECTED_6803,SV2V_UNCONNECTED_6804,
  SV2V_UNCONNECTED_6805,SV2V_UNCONNECTED_6806,SV2V_UNCONNECTED_6807,
  SV2V_UNCONNECTED_6808,SV2V_UNCONNECTED_6809,SV2V_UNCONNECTED_6810,
  SV2V_UNCONNECTED_6811,SV2V_UNCONNECTED_6812,SV2V_UNCONNECTED_6813,
  SV2V_UNCONNECTED_6814,SV2V_UNCONNECTED_6815,SV2V_UNCONNECTED_6816,SV2V_UNCONNECTED_6817,
  SV2V_UNCONNECTED_6818,SV2V_UNCONNECTED_6819,SV2V_UNCONNECTED_6820,
  SV2V_UNCONNECTED_6821,SV2V_UNCONNECTED_6822,SV2V_UNCONNECTED_6823,
  SV2V_UNCONNECTED_6824,SV2V_UNCONNECTED_6825,SV2V_UNCONNECTED_6826,
  SV2V_UNCONNECTED_6827,SV2V_UNCONNECTED_6828,SV2V_UNCONNECTED_6829,
  SV2V_UNCONNECTED_6830,SV2V_UNCONNECTED_6831,SV2V_UNCONNECTED_6832,
  SV2V_UNCONNECTED_6833,SV2V_UNCONNECTED_6834,SV2V_UNCONNECTED_6835,
  SV2V_UNCONNECTED_6836,SV2V_UNCONNECTED_6837,SV2V_UNCONNECTED_6838,
  SV2V_UNCONNECTED_6839,SV2V_UNCONNECTED_6840,SV2V_UNCONNECTED_6841,
  SV2V_UNCONNECTED_6842,SV2V_UNCONNECTED_6843,SV2V_UNCONNECTED_6844,
  SV2V_UNCONNECTED_6845,SV2V_UNCONNECTED_6846,SV2V_UNCONNECTED_6847,
  SV2V_UNCONNECTED_6848,SV2V_UNCONNECTED_6849,SV2V_UNCONNECTED_6850,
  SV2V_UNCONNECTED_6851,SV2V_UNCONNECTED_6852,SV2V_UNCONNECTED_6853,
  SV2V_UNCONNECTED_6854,SV2V_UNCONNECTED_6855,SV2V_UNCONNECTED_6856,SV2V_UNCONNECTED_6857,
  SV2V_UNCONNECTED_6858,SV2V_UNCONNECTED_6859,SV2V_UNCONNECTED_6860,
  SV2V_UNCONNECTED_6861,SV2V_UNCONNECTED_6862,SV2V_UNCONNECTED_6863,
  SV2V_UNCONNECTED_6864,SV2V_UNCONNECTED_6865,SV2V_UNCONNECTED_6866,
  SV2V_UNCONNECTED_6867,SV2V_UNCONNECTED_6868,SV2V_UNCONNECTED_6869,
  SV2V_UNCONNECTED_6870,SV2V_UNCONNECTED_6871,SV2V_UNCONNECTED_6872,
  SV2V_UNCONNECTED_6873,SV2V_UNCONNECTED_6874,SV2V_UNCONNECTED_6875,
  SV2V_UNCONNECTED_6876,SV2V_UNCONNECTED_6877,SV2V_UNCONNECTED_6878,
  SV2V_UNCONNECTED_6879,SV2V_UNCONNECTED_6880,SV2V_UNCONNECTED_6881,
  SV2V_UNCONNECTED_6882,SV2V_UNCONNECTED_6883,SV2V_UNCONNECTED_6884,
  SV2V_UNCONNECTED_6885,SV2V_UNCONNECTED_6886,SV2V_UNCONNECTED_6887,
  SV2V_UNCONNECTED_6888,SV2V_UNCONNECTED_6889,SV2V_UNCONNECTED_6890,
  SV2V_UNCONNECTED_6891,SV2V_UNCONNECTED_6892,SV2V_UNCONNECTED_6893,
  SV2V_UNCONNECTED_6894,SV2V_UNCONNECTED_6895,SV2V_UNCONNECTED_6896,SV2V_UNCONNECTED_6897,
  SV2V_UNCONNECTED_6898,SV2V_UNCONNECTED_6899,SV2V_UNCONNECTED_6900,
  SV2V_UNCONNECTED_6901,SV2V_UNCONNECTED_6902,SV2V_UNCONNECTED_6903,
  SV2V_UNCONNECTED_6904,SV2V_UNCONNECTED_6905,SV2V_UNCONNECTED_6906,
  SV2V_UNCONNECTED_6907,SV2V_UNCONNECTED_6908,SV2V_UNCONNECTED_6909,
  SV2V_UNCONNECTED_6910,SV2V_UNCONNECTED_6911,SV2V_UNCONNECTED_6912,
  SV2V_UNCONNECTED_6913,SV2V_UNCONNECTED_6914,SV2V_UNCONNECTED_6915,
  SV2V_UNCONNECTED_6916,SV2V_UNCONNECTED_6917,SV2V_UNCONNECTED_6918,
  SV2V_UNCONNECTED_6919,SV2V_UNCONNECTED_6920,SV2V_UNCONNECTED_6921,
  SV2V_UNCONNECTED_6922,SV2V_UNCONNECTED_6923,SV2V_UNCONNECTED_6924,
  SV2V_UNCONNECTED_6925,SV2V_UNCONNECTED_6926,SV2V_UNCONNECTED_6927,
  SV2V_UNCONNECTED_6928,SV2V_UNCONNECTED_6929,SV2V_UNCONNECTED_6930,
  SV2V_UNCONNECTED_6931,SV2V_UNCONNECTED_6932,SV2V_UNCONNECTED_6933,
  SV2V_UNCONNECTED_6934,SV2V_UNCONNECTED_6935,SV2V_UNCONNECTED_6936,SV2V_UNCONNECTED_6937,
  SV2V_UNCONNECTED_6938,SV2V_UNCONNECTED_6939,SV2V_UNCONNECTED_6940,
  SV2V_UNCONNECTED_6941,SV2V_UNCONNECTED_6942,SV2V_UNCONNECTED_6943,
  SV2V_UNCONNECTED_6944,SV2V_UNCONNECTED_6945,SV2V_UNCONNECTED_6946,
  SV2V_UNCONNECTED_6947,SV2V_UNCONNECTED_6948,SV2V_UNCONNECTED_6949,
  SV2V_UNCONNECTED_6950,SV2V_UNCONNECTED_6951,SV2V_UNCONNECTED_6952,
  SV2V_UNCONNECTED_6953,SV2V_UNCONNECTED_6954,SV2V_UNCONNECTED_6955,
  SV2V_UNCONNECTED_6956,SV2V_UNCONNECTED_6957,SV2V_UNCONNECTED_6958,
  SV2V_UNCONNECTED_6959,SV2V_UNCONNECTED_6960,SV2V_UNCONNECTED_6961,
  SV2V_UNCONNECTED_6962,SV2V_UNCONNECTED_6963,SV2V_UNCONNECTED_6964,
  SV2V_UNCONNECTED_6965,SV2V_UNCONNECTED_6966,SV2V_UNCONNECTED_6967,
  SV2V_UNCONNECTED_6968,SV2V_UNCONNECTED_6969,SV2V_UNCONNECTED_6970,
  SV2V_UNCONNECTED_6971,SV2V_UNCONNECTED_6972,SV2V_UNCONNECTED_6973,
  SV2V_UNCONNECTED_6974,SV2V_UNCONNECTED_6975,SV2V_UNCONNECTED_6976,SV2V_UNCONNECTED_6977,
  SV2V_UNCONNECTED_6978,SV2V_UNCONNECTED_6979,SV2V_UNCONNECTED_6980,
  SV2V_UNCONNECTED_6981,SV2V_UNCONNECTED_6982,SV2V_UNCONNECTED_6983,
  SV2V_UNCONNECTED_6984,SV2V_UNCONNECTED_6985,SV2V_UNCONNECTED_6986,
  SV2V_UNCONNECTED_6987,SV2V_UNCONNECTED_6988,SV2V_UNCONNECTED_6989,
  SV2V_UNCONNECTED_6990,SV2V_UNCONNECTED_6991,SV2V_UNCONNECTED_6992,
  SV2V_UNCONNECTED_6993,SV2V_UNCONNECTED_6994,SV2V_UNCONNECTED_6995,
  SV2V_UNCONNECTED_6996,SV2V_UNCONNECTED_6997,SV2V_UNCONNECTED_6998,
  SV2V_UNCONNECTED_6999,SV2V_UNCONNECTED_7000,SV2V_UNCONNECTED_7001,
  SV2V_UNCONNECTED_7002,SV2V_UNCONNECTED_7003,SV2V_UNCONNECTED_7004,
  SV2V_UNCONNECTED_7005,SV2V_UNCONNECTED_7006,SV2V_UNCONNECTED_7007,
  SV2V_UNCONNECTED_7008,SV2V_UNCONNECTED_7009,SV2V_UNCONNECTED_7010,
  SV2V_UNCONNECTED_7011,SV2V_UNCONNECTED_7012,SV2V_UNCONNECTED_7013,
  SV2V_UNCONNECTED_7014,SV2V_UNCONNECTED_7015,SV2V_UNCONNECTED_7016,SV2V_UNCONNECTED_7017,
  SV2V_UNCONNECTED_7018,SV2V_UNCONNECTED_7019,SV2V_UNCONNECTED_7020,
  SV2V_UNCONNECTED_7021,SV2V_UNCONNECTED_7022,SV2V_UNCONNECTED_7023,
  SV2V_UNCONNECTED_7024,SV2V_UNCONNECTED_7025,SV2V_UNCONNECTED_7026,
  SV2V_UNCONNECTED_7027,SV2V_UNCONNECTED_7028,SV2V_UNCONNECTED_7029,
  SV2V_UNCONNECTED_7030,SV2V_UNCONNECTED_7031,SV2V_UNCONNECTED_7032,
  SV2V_UNCONNECTED_7033,SV2V_UNCONNECTED_7034,SV2V_UNCONNECTED_7035,
  SV2V_UNCONNECTED_7036,SV2V_UNCONNECTED_7037,SV2V_UNCONNECTED_7038,
  SV2V_UNCONNECTED_7039,SV2V_UNCONNECTED_7040,SV2V_UNCONNECTED_7041,
  SV2V_UNCONNECTED_7042,SV2V_UNCONNECTED_7043,SV2V_UNCONNECTED_7044,
  SV2V_UNCONNECTED_7045,SV2V_UNCONNECTED_7046,SV2V_UNCONNECTED_7047,
  SV2V_UNCONNECTED_7048,SV2V_UNCONNECTED_7049,SV2V_UNCONNECTED_7050,
  SV2V_UNCONNECTED_7051,SV2V_UNCONNECTED_7052,SV2V_UNCONNECTED_7053,
  SV2V_UNCONNECTED_7054,SV2V_UNCONNECTED_7055,SV2V_UNCONNECTED_7056,SV2V_UNCONNECTED_7057,
  SV2V_UNCONNECTED_7058,SV2V_UNCONNECTED_7059,SV2V_UNCONNECTED_7060,
  SV2V_UNCONNECTED_7061,SV2V_UNCONNECTED_7062,SV2V_UNCONNECTED_7063,
  SV2V_UNCONNECTED_7064,SV2V_UNCONNECTED_7065,SV2V_UNCONNECTED_7066,
  SV2V_UNCONNECTED_7067,SV2V_UNCONNECTED_7068,SV2V_UNCONNECTED_7069,
  SV2V_UNCONNECTED_7070,SV2V_UNCONNECTED_7071,SV2V_UNCONNECTED_7072,
  SV2V_UNCONNECTED_7073,SV2V_UNCONNECTED_7074,SV2V_UNCONNECTED_7075,
  SV2V_UNCONNECTED_7076,SV2V_UNCONNECTED_7077,SV2V_UNCONNECTED_7078,
  SV2V_UNCONNECTED_7079,SV2V_UNCONNECTED_7080,SV2V_UNCONNECTED_7081,
  SV2V_UNCONNECTED_7082,SV2V_UNCONNECTED_7083,SV2V_UNCONNECTED_7084,
  SV2V_UNCONNECTED_7085,SV2V_UNCONNECTED_7086,SV2V_UNCONNECTED_7087,
  SV2V_UNCONNECTED_7088,SV2V_UNCONNECTED_7089,SV2V_UNCONNECTED_7090,
  SV2V_UNCONNECTED_7091,SV2V_UNCONNECTED_7092,SV2V_UNCONNECTED_7093,
  SV2V_UNCONNECTED_7094,SV2V_UNCONNECTED_7095,SV2V_UNCONNECTED_7096,SV2V_UNCONNECTED_7097,
  SV2V_UNCONNECTED_7098,SV2V_UNCONNECTED_7099,SV2V_UNCONNECTED_7100,
  SV2V_UNCONNECTED_7101,SV2V_UNCONNECTED_7102,SV2V_UNCONNECTED_7103,
  SV2V_UNCONNECTED_7104,SV2V_UNCONNECTED_7105,SV2V_UNCONNECTED_7106,
  SV2V_UNCONNECTED_7107,SV2V_UNCONNECTED_7108,SV2V_UNCONNECTED_7109,
  SV2V_UNCONNECTED_7110,SV2V_UNCONNECTED_7111,SV2V_UNCONNECTED_7112,
  SV2V_UNCONNECTED_7113,SV2V_UNCONNECTED_7114,SV2V_UNCONNECTED_7115,
  SV2V_UNCONNECTED_7116,SV2V_UNCONNECTED_7117,SV2V_UNCONNECTED_7118,
  SV2V_UNCONNECTED_7119,SV2V_UNCONNECTED_7120,SV2V_UNCONNECTED_7121,
  SV2V_UNCONNECTED_7122,SV2V_UNCONNECTED_7123,SV2V_UNCONNECTED_7124,
  SV2V_UNCONNECTED_7125,SV2V_UNCONNECTED_7126,SV2V_UNCONNECTED_7127,
  SV2V_UNCONNECTED_7128,SV2V_UNCONNECTED_7129,SV2V_UNCONNECTED_7130,
  SV2V_UNCONNECTED_7131,SV2V_UNCONNECTED_7132,SV2V_UNCONNECTED_7133,
  SV2V_UNCONNECTED_7134,SV2V_UNCONNECTED_7135,SV2V_UNCONNECTED_7136,SV2V_UNCONNECTED_7137,
  SV2V_UNCONNECTED_7138,SV2V_UNCONNECTED_7139,SV2V_UNCONNECTED_7140,
  SV2V_UNCONNECTED_7141,SV2V_UNCONNECTED_7142,SV2V_UNCONNECTED_7143,
  SV2V_UNCONNECTED_7144,SV2V_UNCONNECTED_7145,SV2V_UNCONNECTED_7146,
  SV2V_UNCONNECTED_7147,SV2V_UNCONNECTED_7148,SV2V_UNCONNECTED_7149,
  SV2V_UNCONNECTED_7150,SV2V_UNCONNECTED_7151,SV2V_UNCONNECTED_7152,
  SV2V_UNCONNECTED_7153,SV2V_UNCONNECTED_7154,SV2V_UNCONNECTED_7155,
  SV2V_UNCONNECTED_7156,SV2V_UNCONNECTED_7157,SV2V_UNCONNECTED_7158,
  SV2V_UNCONNECTED_7159,SV2V_UNCONNECTED_7160,SV2V_UNCONNECTED_7161,
  SV2V_UNCONNECTED_7162,SV2V_UNCONNECTED_7163,SV2V_UNCONNECTED_7164,
  SV2V_UNCONNECTED_7165,SV2V_UNCONNECTED_7166,SV2V_UNCONNECTED_7167,
  SV2V_UNCONNECTED_7168,SV2V_UNCONNECTED_7169,SV2V_UNCONNECTED_7170,
  SV2V_UNCONNECTED_7171,SV2V_UNCONNECTED_7172,SV2V_UNCONNECTED_7173,
  SV2V_UNCONNECTED_7174,SV2V_UNCONNECTED_7175,SV2V_UNCONNECTED_7176,SV2V_UNCONNECTED_7177,
  SV2V_UNCONNECTED_7178,SV2V_UNCONNECTED_7179,SV2V_UNCONNECTED_7180,
  SV2V_UNCONNECTED_7181,SV2V_UNCONNECTED_7182,SV2V_UNCONNECTED_7183,
  SV2V_UNCONNECTED_7184,SV2V_UNCONNECTED_7185,SV2V_UNCONNECTED_7186,
  SV2V_UNCONNECTED_7187,SV2V_UNCONNECTED_7188,SV2V_UNCONNECTED_7189,
  SV2V_UNCONNECTED_7190,SV2V_UNCONNECTED_7191,SV2V_UNCONNECTED_7192,
  SV2V_UNCONNECTED_7193,SV2V_UNCONNECTED_7194,SV2V_UNCONNECTED_7195,
  SV2V_UNCONNECTED_7196,SV2V_UNCONNECTED_7197;
  wire [56:0] T4,T284,T288,T290;
  wire [54:0] sigX3,T445,T31,T693,T322,T309,T310,roundUp_sigY3,T311,T314,T344,T323,T345;
  wire [0:0] roundMask,T446,T14,T682,T684,T206,T698;
  wire [55:55] T104;
  wire [55:2] T6,T697;
  wire [53:6] T9;
  wire [3:0] T15,T541,T542,T543,T544,T545,T546,T547,T548,T116;
  wire [15:0] T16,T118;
  wire [31:0] T17,T109,T179,T279,T280;
  wire [12:0] T19,sExpX3_13,T352,T305,T306,T355,T353,T356;
  wire [13:13] sExpX3;
  wire [7:0] T447,CDom_estNormDist,T20,T117;
  wire [6:0] T448,T450,T451,T452,T453,T454,T455,T456,T457,T458,T459,T460,T461,T462,T463,T464,
  T465,T466,T467,T468,T469,T470,T471,T472,T473,T474,T475,T476,T477,T478,T479,T480,
  T481,T482,T483,T484,T485,T486,T487,T488,T489,T490,T491,T492;
  wire [5:0] T493,T494,T495,T496,T497,T498,T499,T500,T501,T502,T503,T504,T505,T506,T507,T508,
  T509,T510,T511,T512,T513,T514,T515,T516,T517,T518,T519,T520,T521,T522,T523,T524,
  T663;
  wire [2:0] T549,T550,T551,T552,T304;
  wire [1:0] T553,T554,T115,T695,T308;
  wire [107:1] T22;
  wire [108:107] T25;
  wire [161:109] sigSum;
  wire [15:15] T49,T52,T155,T158;
  wire [14:14] T50,T156;
  wire [15:14] T53,T56,T159,T162;
  wire [13:12] T54,T160;
  wire [15:12] T57,T60,T163,T166;
  wire [11:8] T58,T164;
  wire [31:31] T74,T77;
  wire [30:30] T75;
  wire [31:30] T78,T81;
  wire [29:28] T79;
  wire [31:28] T82,T85;
  wire [27:24] T83;
  wire [31:24] T86,T89;
  wire [23:16] T87;
  wire [31:8] absSigSumExtraMask;
  wire [7:7] T136,T139;
  wire [6:6] T137;
  wire [7:6] T140,T143;
  wire [5:4] T141;
  wire [87:32] cFirstNormAbsSigSum;
  wire [87:0] T257,notCDom_neg_cFirstNormAbsSigSum,T269,T258;
  wire [86:0] T681,CDom_firstNormAbsSigSum,notCDom_pos_firstNormAbsSigSum,T205,T181,T185,T227,
  T219,T237,T228,T247,T238;
  wire [53:53] T182;
  wire [85:85] T186;
  wire [43:0] T199;
  wire [161:44] notSigSum;
  wire [21:21] T213;
  wire [86:86] T686,T687,T688,T689;
  wire [55:0] T692;
  wire [9:0] sExpY;
  wire [52:0] sigY3;
  wire [51:0] T390,T394,fractY;
  wire [51:51] T385,T391;
  wire [11:0] T405,T410,T412,T415,T418,T416,T421,T419,T424,T422,T425;
  wire [11:11] T404,T406,T411,T423,T426;
  wire [9:9] T413,T417;
  wire [10:10] T420;
  assign io_exceptionFlags[3] = 1'b0;
  assign { SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, SV2V_UNCONNECTED_16, SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, sigX3_56, T446[0:0], sigX3[54:1] } = { cFirstNormAbsSigSum, T179[31:1] } >> normTo2ShiftDist;
  assign T300 = sExpX3_13 <= { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T695 };
  assign sigX3Shift1 = { sigX3_56, T446[0:0] } == 1'b0;
  assign isZeroY = { sigX3_56, T446[0:0], sigX3[54:54] } == 1'b0;
  assign T400 = { T304[1:0], sExpY } < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign N374 = io_fromPreMul_highExpB[1] | io_fromPreMul_highExpB[2];
  assign N375 = io_fromPreMul_highExpB[0] | N374;
  assign N376 = ~N375;
  assign N377 = io_fromPreMul_highExpA[1] | io_fromPreMul_highExpA[2];
  assign N378 = io_fromPreMul_highExpA[0] | N377;
  assign N379 = ~N378;
  assign N380 = ~T304[1];
  assign N381 = ~T304[0];
  assign N382 = N380 | T304[2];
  assign N383 = N381 | N382;
  assign N384 = ~N383;
  assign N385 = io_fromPreMul_highExpC[1] & io_fromPreMul_highExpC[2];
  assign N386 = io_fromPreMul_highExpA[1] & io_fromPreMul_highExpA[2];
  assign N387 = io_fromPreMul_highExpB[1] & io_fromPreMul_highExpB[2];
  assign N388 = T308[0] | T308[1];
  assign N389 = ~N388;
  assign N390 = T288[55] | T288[56];
  assign N391 = T288[54] | N390;
  assign N392 = T288[53] | N391;
  assign N393 = T288[52] | N392;
  assign N394 = T288[51] | N393;
  assign N395 = T288[50] | N394;
  assign N396 = T288[49] | N395;
  assign N397 = T288[48] | N396;
  assign N398 = T288[47] | N397;
  assign N399 = T288[46] | N398;
  assign N400 = T288[45] | N399;
  assign N401 = T288[44] | N400;
  assign N402 = T288[43] | N401;
  assign N403 = T288[42] | N402;
  assign N404 = T288[41] | N403;
  assign N405 = T288[40] | N404;
  assign N406 = T288[39] | N405;
  assign N407 = T288[38] | N406;
  assign N408 = T288[37] | N407;
  assign N409 = T288[36] | N408;
  assign N410 = T288[35] | N409;
  assign N411 = T288[34] | N410;
  assign N412 = T288[33] | N411;
  assign N413 = T288[32] | N412;
  assign N414 = T288[31] | N413;
  assign N415 = T288[30] | N414;
  assign N416 = T288[29] | N415;
  assign N417 = T288[28] | N416;
  assign N418 = T288[27] | N417;
  assign N419 = T288[26] | N418;
  assign N420 = T288[25] | N419;
  assign N421 = T288[24] | N420;
  assign N422 = T288[23] | N421;
  assign N423 = T288[22] | N422;
  assign N424 = T288[21] | N423;
  assign N425 = T288[20] | N424;
  assign N426 = T288[19] | N425;
  assign N427 = T288[18] | N426;
  assign N428 = T288[17] | N427;
  assign N429 = T288[16] | N428;
  assign N430 = T288[15] | N429;
  assign N431 = T288[14] | N430;
  assign N432 = T288[13] | N431;
  assign N433 = T288[12] | N432;
  assign N434 = T288[11] | N433;
  assign N435 = T288[10] | N434;
  assign N436 = T288[9] | N435;
  assign N437 = T288[8] | N436;
  assign N438 = T288[7] | N437;
  assign N439 = T288[6] | N438;
  assign N440 = T288[5] | N439;
  assign N441 = T288[4] | N440;
  assign N442 = T288[3] | N441;
  assign N443 = T288[2] | N442;
  assign N444 = T288[1] | N443;
  assign N445 = T288[0] | N444;
  assign N446 = ~N445;
  assign N447 = T284[55] | T284[56];
  assign N448 = T284[54] | N447;
  assign N449 = T284[53] | N448;
  assign N450 = T284[52] | N449;
  assign N451 = T284[51] | N450;
  assign N452 = T284[50] | N451;
  assign N453 = T284[49] | N452;
  assign N454 = T284[48] | N453;
  assign N455 = T284[47] | N454;
  assign N456 = T284[46] | N455;
  assign N457 = T284[45] | N456;
  assign N458 = T284[44] | N457;
  assign N459 = T284[43] | N458;
  assign N460 = T284[42] | N459;
  assign N461 = T284[41] | N460;
  assign N462 = T284[40] | N461;
  assign N463 = T284[39] | N462;
  assign N464 = T284[38] | N463;
  assign N465 = T284[37] | N464;
  assign N466 = T284[36] | N465;
  assign N467 = T284[35] | N466;
  assign N468 = T284[34] | N467;
  assign N469 = T284[33] | N468;
  assign N470 = T284[32] | N469;
  assign N471 = T284[31] | N470;
  assign N472 = T284[30] | N471;
  assign N473 = T284[29] | N472;
  assign N474 = T284[28] | N473;
  assign N475 = T284[27] | N474;
  assign N476 = T284[26] | N475;
  assign N477 = T284[25] | N476;
  assign N478 = T284[24] | N477;
  assign N479 = T284[23] | N478;
  assign N480 = T284[22] | N479;
  assign N481 = T284[21] | N480;
  assign N482 = T284[20] | N481;
  assign N483 = T284[19] | N482;
  assign N484 = T284[18] | N483;
  assign N485 = T284[17] | N484;
  assign N486 = T284[16] | N485;
  assign N487 = T284[15] | N486;
  assign N488 = T284[14] | N487;
  assign N489 = T284[13] | N488;
  assign N490 = T284[12] | N489;
  assign N491 = T284[11] | N490;
  assign N492 = T284[10] | N491;
  assign N493 = T284[9] | N492;
  assign N494 = T284[8] | N493;
  assign N495 = T284[7] | N494;
  assign N496 = T284[6] | N495;
  assign N497 = T284[5] | N496;
  assign N498 = T284[4] | N497;
  assign N499 = T284[3] | N498;
  assign N500 = T284[2] | N499;
  assign N501 = T284[1] | N500;
  assign N502 = T284[0] | N501;
  assign N503 = T4[55] | T4[56];
  assign N504 = T4[54] | N503;
  assign N505 = T4[53] | N504;
  assign N506 = T4[52] | N505;
  assign N507 = T4[51] | N506;
  assign N508 = T4[50] | N507;
  assign N509 = T4[49] | N508;
  assign N510 = T4[48] | N509;
  assign N511 = T4[47] | N510;
  assign N512 = T4[46] | N511;
  assign N513 = T4[45] | N512;
  assign N514 = T4[44] | N513;
  assign N515 = T4[43] | N514;
  assign N516 = T4[42] | N515;
  assign N517 = T4[41] | N516;
  assign N518 = T4[40] | N517;
  assign N519 = T4[39] | N518;
  assign N520 = T4[38] | N519;
  assign N521 = T4[37] | N520;
  assign N522 = T4[36] | N521;
  assign N523 = T4[35] | N522;
  assign N524 = T4[34] | N523;
  assign N525 = T4[33] | N524;
  assign N526 = T4[32] | N525;
  assign N527 = T4[31] | N526;
  assign N528 = T4[30] | N527;
  assign N529 = T4[29] | N528;
  assign N530 = T4[28] | N529;
  assign N531 = T4[27] | N530;
  assign N532 = T4[26] | N531;
  assign N533 = T4[25] | N532;
  assign N534 = T4[24] | N533;
  assign N535 = T4[23] | N534;
  assign N536 = T4[22] | N535;
  assign N537 = T4[21] | N536;
  assign N538 = T4[20] | N537;
  assign N539 = T4[19] | N538;
  assign N540 = T4[18] | N539;
  assign N541 = T4[17] | N540;
  assign N542 = T4[16] | N541;
  assign N543 = T4[15] | N542;
  assign N544 = T4[14] | N543;
  assign N545 = T4[13] | N544;
  assign N546 = T4[12] | N545;
  assign N547 = T4[11] | N546;
  assign N548 = T4[10] | N547;
  assign N549 = T4[9] | N548;
  assign N550 = T4[8] | N549;
  assign N551 = T4[7] | N550;
  assign N552 = T4[6] | N551;
  assign N553 = T4[5] | N552;
  assign N554 = T4[4] | N553;
  assign N555 = T4[3] | N554;
  assign N556 = T4[2] | N555;
  assign N557 = T4[1] | N556;
  assign N558 = T4[0] | N557;
  assign N559 = io_fromPreMul_roundingMode[0] | io_fromPreMul_roundingMode[1];
  assign N560 = ~N559;
  assign N561 = io_fromPreMul_roundingMode[0] & io_fromPreMul_roundingMode[1];
  assign N562 = T279[30] | T279[31];
  assign N563 = T279[29] | N562;
  assign N564 = T279[28] | N563;
  assign N565 = T279[27] | N564;
  assign N566 = T279[26] | N565;
  assign N567 = T279[25] | N566;
  assign N568 = T279[24] | N567;
  assign N569 = T279[23] | N568;
  assign N570 = T279[22] | N569;
  assign N571 = T279[21] | N570;
  assign N572 = T279[20] | N571;
  assign N573 = T279[19] | N572;
  assign N574 = T279[18] | N573;
  assign N575 = T279[17] | N574;
  assign N576 = T279[16] | N575;
  assign N577 = T279[15] | N576;
  assign N578 = T279[14] | N577;
  assign N579 = T279[13] | N578;
  assign N580 = T279[12] | N579;
  assign N581 = T279[11] | N580;
  assign N582 = T279[10] | N581;
  assign N583 = T279[9] | N582;
  assign N584 = T279[8] | N583;
  assign N585 = T279[7] | N584;
  assign N586 = T279[6] | N585;
  assign N587 = T279[5] | N586;
  assign N588 = T279[4] | N587;
  assign N589 = T279[3] | N588;
  assign N590 = T279[2] | N589;
  assign N591 = T279[1] | N590;
  assign N592 = T279[0] | N591;
  assign N593 = ~N592;
  assign N594 = T109[30] | T109[31];
  assign N595 = T109[29] | N594;
  assign N596 = T109[28] | N595;
  assign N597 = T109[27] | N596;
  assign N598 = T109[26] | N597;
  assign N599 = T109[25] | N598;
  assign N600 = T109[24] | N599;
  assign N601 = T109[23] | N600;
  assign N602 = T109[22] | N601;
  assign N603 = T109[21] | N602;
  assign N604 = T109[20] | N603;
  assign N605 = T109[19] | N604;
  assign N606 = T109[18] | N605;
  assign N607 = T109[17] | N606;
  assign N608 = T109[16] | N607;
  assign N609 = T109[15] | N608;
  assign N610 = T109[14] | N609;
  assign N611 = T109[13] | N610;
  assign N612 = T109[12] | N611;
  assign N613 = T109[11] | N612;
  assign N614 = T109[10] | N613;
  assign N615 = T109[9] | N614;
  assign N616 = T109[8] | N615;
  assign N617 = T109[7] | N616;
  assign N618 = T109[6] | N617;
  assign N619 = T109[5] | N618;
  assign N620 = T109[4] | N619;
  assign N621 = T109[3] | N620;
  assign N622 = T109[2] | N621;
  assign N623 = T109[1] | N622;
  assign N624 = T109[0] | N623;
  assign N625 = ~io_fromPreMul_roundingMode[1];
  assign N626 = io_fromPreMul_roundingMode[0] | N625;
  assign N627 = ~N626;
  assign N628 = io_fromPreMul_highExpC[1] | io_fromPreMul_highExpC[2];
  assign N629 = io_fromPreMul_highExpC[0] | N628;
  assign N630 = ~N629;
  assign { SV2V_UNCONNECTED_32, absSigSumExtraMask_1, T115, T116, T117, T118 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> normTo2ShiftDist;
  assign N631 = T199[10] | T199[11];
  assign N632 = T199[9] | N631;
  assign N633 = T199[8] | N632;
  assign N634 = T199[7] | N633;
  assign N635 = T199[6] | N634;
  assign N636 = T199[5] | N635;
  assign N637 = T199[4] | N636;
  assign N638 = T199[3] | N637;
  assign N639 = T199[2] | N638;
  assign N640 = T199[1] | N639;
  assign { SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, SV2V_UNCONNECTED_49, SV2V_UNCONNECTED_50, SV2V_UNCONNECTED_51, SV2V_UNCONNECTED_52, SV2V_UNCONNECTED_53, SV2V_UNCONNECTED_54, SV2V_UNCONNECTED_55, SV2V_UNCONNECTED_56, SV2V_UNCONNECTED_57, SV2V_UNCONNECTED_58, SV2V_UNCONNECTED_59, SV2V_UNCONNECTED_60, SV2V_UNCONNECTED_61, SV2V_UNCONNECTED_62, SV2V_UNCONNECTED_63, SV2V_UNCONNECTED_64, SV2V_UNCONNECTED_65, SV2V_UNCONNECTED_66, SV2V_UNCONNECTED_67, SV2V_UNCONNECTED_68, SV2V_UNCONNECTED_69, SV2V_UNCONNECTED_70, SV2V_UNCONNECTED_71, SV2V_UNCONNECTED_72, SV2V_UNCONNECTED_73, SV2V_UNCONNECTED_74, SV2V_UNCONNECTED_75, SV2V_UNCONNECTED_76, SV2V_UNCONNECTED_77, SV2V_UNCONNECTED_78, SV2V_UNCONNECTED_79, SV2V_UNCONNECTED_80, SV2V_UNCONNECTED_81, SV2V_UNCONNECTED_82, SV2V_UNCONNECTED_83, SV2V_UNCONNECTED_84, SV2V_UNCONNECTED_85, SV2V_UNCONNECTED_86, SV2V_UNCONNECTED_87, SV2V_UNCONNECTED_88, SV2V_UNCONNECTED_89, SV2V_UNCONNECTED_90, SV2V_UNCONNECTED_91, SV2V_UNCONNECTED_92, SV2V_UNCONNECTED_93, SV2V_UNCONNECTED_94, SV2V_UNCONNECTED_95, SV2V_UNCONNECTED_96, SV2V_UNCONNECTED_97, SV2V_UNCONNECTED_98, SV2V_UNCONNECTED_99, SV2V_UNCONNECTED_100, SV2V_UNCONNECTED_101, SV2V_UNCONNECTED_102, SV2V_UNCONNECTED_103, SV2V_UNCONNECTED_104, SV2V_UNCONNECTED_105, SV2V_UNCONNECTED_106, SV2V_UNCONNECTED_107, SV2V_UNCONNECTED_108, SV2V_UNCONNECTED_109, SV2V_UNCONNECTED_110, SV2V_UNCONNECTED_111, SV2V_UNCONNECTED_112, SV2V_UNCONNECTED_113, SV2V_UNCONNECTED_114, SV2V_UNCONNECTED_115, SV2V_UNCONNECTED_116, SV2V_UNCONNECTED_117, SV2V_UNCONNECTED_118, SV2V_UNCONNECTED_119, SV2V_UNCONNECTED_120, SV2V_UNCONNECTED_121, SV2V_UNCONNECTED_122, SV2V_UNCONNECTED_123, SV2V_UNCONNECTED_124, SV2V_UNCONNECTED_125, SV2V_UNCONNECTED_126, SV2V_UNCONNECTED_127, SV2V_UNCONNECTED_128, SV2V_UNCONNECTED_129, SV2V_UNCONNECTED_130, SV2V_UNCONNECTED_131, SV2V_UNCONNECTED_132, SV2V_UNCONNECTED_133, SV2V_UNCONNECTED_134, SV2V_UNCONNECTED_135, SV2V_UNCONNECTED_136, SV2V_UNCONNECTED_137, SV2V_UNCONNECTED_138, SV2V_UNCONNECTED_139, SV2V_UNCONNECTED_140, SV2V_UNCONNECTED_141, SV2V_UNCONNECTED_142, SV2V_UNCONNECTED_143, SV2V_UNCONNECTED_144, SV2V_UNCONNECTED_145, SV2V_UNCONNECTED_146, SV2V_UNCONNECTED_147, SV2V_UNCONNECTED_148, SV2V_UNCONNECTED_149, SV2V_UNCONNECTED_150, SV2V_UNCONNECTED_151, SV2V_UNCONNECTED_152, SV2V_UNCONNECTED_153, SV2V_UNCONNECTED_154, SV2V_UNCONNECTED_155, SV2V_UNCONNECTED_156, SV2V_UNCONNECTED_157, SV2V_UNCONNECTED_158, SV2V_UNCONNECTED_159, SV2V_UNCONNECTED_160, SV2V_UNCONNECTED_161, SV2V_UNCONNECTED_162, SV2V_UNCONNECTED_163, SV2V_UNCONNECTED_164, SV2V_UNCONNECTED_165, SV2V_UNCONNECTED_166, SV2V_UNCONNECTED_167, SV2V_UNCONNECTED_168, SV2V_UNCONNECTED_169, SV2V_UNCONNECTED_170, SV2V_UNCONNECTED_171, SV2V_UNCONNECTED_172, SV2V_UNCONNECTED_173, SV2V_UNCONNECTED_174, SV2V_UNCONNECTED_175, SV2V_UNCONNECTED_176, SV2V_UNCONNECTED_177, SV2V_UNCONNECTED_178, SV2V_UNCONNECTED_179, SV2V_UNCONNECTED_180, SV2V_UNCONNECTED_181, SV2V_UNCONNECTED_182, SV2V_UNCONNECTED_183, SV2V_UNCONNECTED_184, SV2V_UNCONNECTED_185, SV2V_UNCONNECTED_186, SV2V_UNCONNECTED_187, SV2V_UNCONNECTED_188, SV2V_UNCONNECTED_189, SV2V_UNCONNECTED_190, SV2V_UNCONNECTED_191, SV2V_UNCONNECTED_192, SV2V_UNCONNECTED_193, SV2V_UNCONNECTED_194, SV2V_UNCONNECTED_195, SV2V_UNCONNECTED_196, SV2V_UNCONNECTED_197, SV2V_UNCONNECTED_198, SV2V_UNCONNECTED_199, SV2V_UNCONNECTED_200, SV2V_UNCONNECTED_201, SV2V_UNCONNECTED_202, SV2V_UNCONNECTED_203, SV2V_UNCONNECTED_204, SV2V_UNCONNECTED_205, SV2V_UNCONNECTED_206, SV2V_UNCONNECTED_207, SV2V_UNCONNECTED_208, SV2V_UNCONNECTED_209, SV2V_UNCONNECTED_210, SV2V_UNCONNECTED_211, SV2V_UNCONNECTED_212, SV2V_UNCONNECTED_213, SV2V_UNCONNECTED_214, SV2V_UNCONNECTED_215, SV2V_UNCONNECTED_216, SV2V_UNCONNECTED_217, SV2V_UNCONNECTED_218, SV2V_UNCONNECTED_219, SV2V_UNCONNECTED_220, SV2V_UNCONNECTED_221, SV2V_UNCONNECTED_222, SV2V_UNCONNECTED_223, SV2V_UNCONNECTED_224, SV2V_UNCONNECTED_225, SV2V_UNCONNECTED_226, SV2V_UNCONNECTED_227, SV2V_UNCONNECTED_228, SV2V_UNCONNECTED_229, SV2V_UNCONNECTED_230, SV2V_UNCONNECTED_231, SV2V_UNCONNECTED_232, SV2V_UNCONNECTED_233, SV2V_UNCONNECTED_234, SV2V_UNCONNECTED_235, SV2V_UNCONNECTED_236, SV2V_UNCONNECTED_237, SV2V_UNCONNECTED_238, SV2V_UNCONNECTED_239, SV2V_UNCONNECTED_240, SV2V_UNCONNECTED_241, SV2V_UNCONNECTED_242, SV2V_UNCONNECTED_243, SV2V_UNCONNECTED_244, SV2V_UNCONNECTED_245, SV2V_UNCONNECTED_246, SV2V_UNCONNECTED_247, SV2V_UNCONNECTED_248, SV2V_UNCONNECTED_249, SV2V_UNCONNECTED_250, SV2V_UNCONNECTED_251, SV2V_UNCONNECTED_252, SV2V_UNCONNECTED_253, SV2V_UNCONNECTED_254, SV2V_UNCONNECTED_255, SV2V_UNCONNECTED_256, SV2V_UNCONNECTED_257, SV2V_UNCONNECTED_258, SV2V_UNCONNECTED_259, SV2V_UNCONNECTED_260, SV2V_UNCONNECTED_261, SV2V_UNCONNECTED_262, SV2V_UNCONNECTED_263, SV2V_UNCONNECTED_264, SV2V_UNCONNECTED_265, SV2V_UNCONNECTED_266, SV2V_UNCONNECTED_267, SV2V_UNCONNECTED_268, SV2V_UNCONNECTED_269, SV2V_UNCONNECTED_270, SV2V_UNCONNECTED_271, SV2V_UNCONNECTED_272, SV2V_UNCONNECTED_273, SV2V_UNCONNECTED_274, SV2V_UNCONNECTED_275, SV2V_UNCONNECTED_276, SV2V_UNCONNECTED_277, SV2V_UNCONNECTED_278, SV2V_UNCONNECTED_279, SV2V_UNCONNECTED_280, SV2V_UNCONNECTED_281, SV2V_UNCONNECTED_282, SV2V_UNCONNECTED_283, SV2V_UNCONNECTED_284, SV2V_UNCONNECTED_285, SV2V_UNCONNECTED_286, SV2V_UNCONNECTED_287, SV2V_UNCONNECTED_288, SV2V_UNCONNECTED_289, SV2V_UNCONNECTED_290, SV2V_UNCONNECTED_291, SV2V_UNCONNECTED_292, SV2V_UNCONNECTED_293, SV2V_UNCONNECTED_294, SV2V_UNCONNECTED_295, SV2V_UNCONNECTED_296, SV2V_UNCONNECTED_297, SV2V_UNCONNECTED_298, SV2V_UNCONNECTED_299, SV2V_UNCONNECTED_300, SV2V_UNCONNECTED_301, SV2V_UNCONNECTED_302, SV2V_UNCONNECTED_303, SV2V_UNCONNECTED_304, SV2V_UNCONNECTED_305, SV2V_UNCONNECTED_306, SV2V_UNCONNECTED_307, SV2V_UNCONNECTED_308, SV2V_UNCONNECTED_309, SV2V_UNCONNECTED_310, SV2V_UNCONNECTED_311, SV2V_UNCONNECTED_312, SV2V_UNCONNECTED_313, SV2V_UNCONNECTED_314, SV2V_UNCONNECTED_315, SV2V_UNCONNECTED_316, SV2V_UNCONNECTED_317, SV2V_UNCONNECTED_318, SV2V_UNCONNECTED_319, SV2V_UNCONNECTED_320, SV2V_UNCONNECTED_321, SV2V_UNCONNECTED_322, SV2V_UNCONNECTED_323, SV2V_UNCONNECTED_324, SV2V_UNCONNECTED_325, SV2V_UNCONNECTED_326, SV2V_UNCONNECTED_327, SV2V_UNCONNECTED_328, SV2V_UNCONNECTED_329, SV2V_UNCONNECTED_330, SV2V_UNCONNECTED_331, SV2V_UNCONNECTED_332, SV2V_UNCONNECTED_333, SV2V_UNCONNECTED_334, SV2V_UNCONNECTED_335, SV2V_UNCONNECTED_336, SV2V_UNCONNECTED_337, SV2V_UNCONNECTED_338, SV2V_UNCONNECTED_339, SV2V_UNCONNECTED_340, SV2V_UNCONNECTED_341, SV2V_UNCONNECTED_342, SV2V_UNCONNECTED_343, SV2V_UNCONNECTED_344, SV2V_UNCONNECTED_345, SV2V_UNCONNECTED_346, SV2V_UNCONNECTED_347, SV2V_UNCONNECTED_348, SV2V_UNCONNECTED_349, SV2V_UNCONNECTED_350, SV2V_UNCONNECTED_351, SV2V_UNCONNECTED_352, SV2V_UNCONNECTED_353, SV2V_UNCONNECTED_354, SV2V_UNCONNECTED_355, SV2V_UNCONNECTED_356, SV2V_UNCONNECTED_357, SV2V_UNCONNECTED_358, SV2V_UNCONNECTED_359, SV2V_UNCONNECTED_360, SV2V_UNCONNECTED_361, SV2V_UNCONNECTED_362, SV2V_UNCONNECTED_363, SV2V_UNCONNECTED_364, SV2V_UNCONNECTED_365, SV2V_UNCONNECTED_366, SV2V_UNCONNECTED_367, SV2V_UNCONNECTED_368, SV2V_UNCONNECTED_369, SV2V_UNCONNECTED_370, SV2V_UNCONNECTED_371, SV2V_UNCONNECTED_372, SV2V_UNCONNECTED_373, SV2V_UNCONNECTED_374, SV2V_UNCONNECTED_375, SV2V_UNCONNECTED_376, SV2V_UNCONNECTED_377, SV2V_UNCONNECTED_378, SV2V_UNCONNECTED_379, SV2V_UNCONNECTED_380, SV2V_UNCONNECTED_381, SV2V_UNCONNECTED_382, SV2V_UNCONNECTED_383, SV2V_UNCONNECTED_384, SV2V_UNCONNECTED_385, SV2V_UNCONNECTED_386, SV2V_UNCONNECTED_387, SV2V_UNCONNECTED_388, SV2V_UNCONNECTED_389, SV2V_UNCONNECTED_390, SV2V_UNCONNECTED_391, SV2V_UNCONNECTED_392, SV2V_UNCONNECTED_393, SV2V_UNCONNECTED_394, SV2V_UNCONNECTED_395, SV2V_UNCONNECTED_396, SV2V_UNCONNECTED_397, SV2V_UNCONNECTED_398, SV2V_UNCONNECTED_399, SV2V_UNCONNECTED_400, SV2V_UNCONNECTED_401, SV2V_UNCONNECTED_402, SV2V_UNCONNECTED_403, SV2V_UNCONNECTED_404, SV2V_UNCONNECTED_405, SV2V_UNCONNECTED_406, SV2V_UNCONNECTED_407, SV2V_UNCONNECTED_408, SV2V_UNCONNECTED_409, SV2V_UNCONNECTED_410, SV2V_UNCONNECTED_411, SV2V_UNCONNECTED_412, SV2V_UNCONNECTED_413, SV2V_UNCONNECTED_414, SV2V_UNCONNECTED_415, SV2V_UNCONNECTED_416, SV2V_UNCONNECTED_417, SV2V_UNCONNECTED_418, SV2V_UNCONNECTED_419, SV2V_UNCONNECTED_420, SV2V_UNCONNECTED_421, SV2V_UNCONNECTED_422, SV2V_UNCONNECTED_423, SV2V_UNCONNECTED_424, SV2V_UNCONNECTED_425, SV2V_UNCONNECTED_426, SV2V_UNCONNECTED_427, SV2V_UNCONNECTED_428, SV2V_UNCONNECTED_429, SV2V_UNCONNECTED_430, SV2V_UNCONNECTED_431, SV2V_UNCONNECTED_432, SV2V_UNCONNECTED_433, SV2V_UNCONNECTED_434, SV2V_UNCONNECTED_435, SV2V_UNCONNECTED_436, SV2V_UNCONNECTED_437, SV2V_UNCONNECTED_438, SV2V_UNCONNECTED_439, SV2V_UNCONNECTED_440, SV2V_UNCONNECTED_441, SV2V_UNCONNECTED_442, SV2V_UNCONNECTED_443, SV2V_UNCONNECTED_444, SV2V_UNCONNECTED_445, SV2V_UNCONNECTED_446, SV2V_UNCONNECTED_447, SV2V_UNCONNECTED_448, SV2V_UNCONNECTED_449, SV2V_UNCONNECTED_450, SV2V_UNCONNECTED_451, SV2V_UNCONNECTED_452, SV2V_UNCONNECTED_453, SV2V_UNCONNECTED_454, SV2V_UNCONNECTED_455, SV2V_UNCONNECTED_456, SV2V_UNCONNECTED_457, SV2V_UNCONNECTED_458, SV2V_UNCONNECTED_459, SV2V_UNCONNECTED_460, SV2V_UNCONNECTED_461, SV2V_UNCONNECTED_462, SV2V_UNCONNECTED_463, SV2V_UNCONNECTED_464, SV2V_UNCONNECTED_465, SV2V_UNCONNECTED_466, SV2V_UNCONNECTED_467, SV2V_UNCONNECTED_468, SV2V_UNCONNECTED_469, SV2V_UNCONNECTED_470, SV2V_UNCONNECTED_471, SV2V_UNCONNECTED_472, SV2V_UNCONNECTED_473, SV2V_UNCONNECTED_474, SV2V_UNCONNECTED_475, SV2V_UNCONNECTED_476, SV2V_UNCONNECTED_477, SV2V_UNCONNECTED_478, SV2V_UNCONNECTED_479, SV2V_UNCONNECTED_480, SV2V_UNCONNECTED_481, SV2V_UNCONNECTED_482, SV2V_UNCONNECTED_483, SV2V_UNCONNECTED_484, SV2V_UNCONNECTED_485, SV2V_UNCONNECTED_486, SV2V_UNCONNECTED_487, SV2V_UNCONNECTED_488, SV2V_UNCONNECTED_489, SV2V_UNCONNECTED_490, SV2V_UNCONNECTED_491, SV2V_UNCONNECTED_492, SV2V_UNCONNECTED_493, SV2V_UNCONNECTED_494, SV2V_UNCONNECTED_495, SV2V_UNCONNECTED_496, SV2V_UNCONNECTED_497, SV2V_UNCONNECTED_498, SV2V_UNCONNECTED_499, SV2V_UNCONNECTED_500, SV2V_UNCONNECTED_501, SV2V_UNCONNECTED_502, SV2V_UNCONNECTED_503, SV2V_UNCONNECTED_504, SV2V_UNCONNECTED_505, SV2V_UNCONNECTED_506, SV2V_UNCONNECTED_507, SV2V_UNCONNECTED_508, SV2V_UNCONNECTED_509, SV2V_UNCONNECTED_510, SV2V_UNCONNECTED_511, SV2V_UNCONNECTED_512, SV2V_UNCONNECTED_513, SV2V_UNCONNECTED_514, SV2V_UNCONNECTED_515, SV2V_UNCONNECTED_516, SV2V_UNCONNECTED_517, SV2V_UNCONNECTED_518, SV2V_UNCONNECTED_519, SV2V_UNCONNECTED_520, SV2V_UNCONNECTED_521, SV2V_UNCONNECTED_522, SV2V_UNCONNECTED_523, SV2V_UNCONNECTED_524, SV2V_UNCONNECTED_525, SV2V_UNCONNECTED_526, SV2V_UNCONNECTED_527, SV2V_UNCONNECTED_528, SV2V_UNCONNECTED_529, SV2V_UNCONNECTED_530, SV2V_UNCONNECTED_531, SV2V_UNCONNECTED_532, SV2V_UNCONNECTED_533, SV2V_UNCONNECTED_534, SV2V_UNCONNECTED_535, SV2V_UNCONNECTED_536, SV2V_UNCONNECTED_537, SV2V_UNCONNECTED_538, SV2V_UNCONNECTED_539, SV2V_UNCONNECTED_540, SV2V_UNCONNECTED_541, SV2V_UNCONNECTED_542, SV2V_UNCONNECTED_543, SV2V_UNCONNECTED_544, SV2V_UNCONNECTED_545, SV2V_UNCONNECTED_546, SV2V_UNCONNECTED_547, SV2V_UNCONNECTED_548, SV2V_UNCONNECTED_549, SV2V_UNCONNECTED_550, SV2V_UNCONNECTED_551, SV2V_UNCONNECTED_552, SV2V_UNCONNECTED_553, SV2V_UNCONNECTED_554, SV2V_UNCONNECTED_555, SV2V_UNCONNECTED_556, SV2V_UNCONNECTED_557, SV2V_UNCONNECTED_558, SV2V_UNCONNECTED_559, SV2V_UNCONNECTED_560, SV2V_UNCONNECTED_561, SV2V_UNCONNECTED_562, SV2V_UNCONNECTED_563, SV2V_UNCONNECTED_564, SV2V_UNCONNECTED_565, SV2V_UNCONNECTED_566, SV2V_UNCONNECTED_567, SV2V_UNCONNECTED_568, SV2V_UNCONNECTED_569, SV2V_UNCONNECTED_570, SV2V_UNCONNECTED_571, SV2V_UNCONNECTED_572, SV2V_UNCONNECTED_573, SV2V_UNCONNECTED_574, SV2V_UNCONNECTED_575, SV2V_UNCONNECTED_576, SV2V_UNCONNECTED_577, SV2V_UNCONNECTED_578, SV2V_UNCONNECTED_579, SV2V_UNCONNECTED_580, SV2V_UNCONNECTED_581, SV2V_UNCONNECTED_582, SV2V_UNCONNECTED_583, SV2V_UNCONNECTED_584, SV2V_UNCONNECTED_585, SV2V_UNCONNECTED_586, SV2V_UNCONNECTED_587, SV2V_UNCONNECTED_588, SV2V_UNCONNECTED_589, SV2V_UNCONNECTED_590, SV2V_UNCONNECTED_591, SV2V_UNCONNECTED_592, SV2V_UNCONNECTED_593, SV2V_UNCONNECTED_594, SV2V_UNCONNECTED_595, SV2V_UNCONNECTED_596, SV2V_UNCONNECTED_597, SV2V_UNCONNECTED_598, SV2V_UNCONNECTED_599, SV2V_UNCONNECTED_600, SV2V_UNCONNECTED_601, SV2V_UNCONNECTED_602, SV2V_UNCONNECTED_603, SV2V_UNCONNECTED_604, SV2V_UNCONNECTED_605, SV2V_UNCONNECTED_606, SV2V_UNCONNECTED_607, SV2V_UNCONNECTED_608, SV2V_UNCONNECTED_609, SV2V_UNCONNECTED_610, SV2V_UNCONNECTED_611, SV2V_UNCONNECTED_612, SV2V_UNCONNECTED_613, SV2V_UNCONNECTED_614, SV2V_UNCONNECTED_615, SV2V_UNCONNECTED_616, SV2V_UNCONNECTED_617, SV2V_UNCONNECTED_618, SV2V_UNCONNECTED_619, SV2V_UNCONNECTED_620, SV2V_UNCONNECTED_621, SV2V_UNCONNECTED_622, SV2V_UNCONNECTED_623, SV2V_UNCONNECTED_624, SV2V_UNCONNECTED_625, SV2V_UNCONNECTED_626, SV2V_UNCONNECTED_627, SV2V_UNCONNECTED_628, SV2V_UNCONNECTED_629, SV2V_UNCONNECTED_630, SV2V_UNCONNECTED_631, SV2V_UNCONNECTED_632, SV2V_UNCONNECTED_633, SV2V_UNCONNECTED_634, SV2V_UNCONNECTED_635, SV2V_UNCONNECTED_636, SV2V_UNCONNECTED_637, SV2V_UNCONNECTED_638, SV2V_UNCONNECTED_639, SV2V_UNCONNECTED_640, SV2V_UNCONNECTED_641, SV2V_UNCONNECTED_642, SV2V_UNCONNECTED_643, SV2V_UNCONNECTED_644, SV2V_UNCONNECTED_645, SV2V_UNCONNECTED_646, SV2V_UNCONNECTED_647, SV2V_UNCONNECTED_648, SV2V_UNCONNECTED_649, SV2V_UNCONNECTED_650, SV2V_UNCONNECTED_651, SV2V_UNCONNECTED_652, SV2V_UNCONNECTED_653, SV2V_UNCONNECTED_654, SV2V_UNCONNECTED_655, SV2V_UNCONNECTED_656, SV2V_UNCONNECTED_657, SV2V_UNCONNECTED_658, SV2V_UNCONNECTED_659, SV2V_UNCONNECTED_660, SV2V_UNCONNECTED_661, SV2V_UNCONNECTED_662, SV2V_UNCONNECTED_663, SV2V_UNCONNECTED_664, SV2V_UNCONNECTED_665, SV2V_UNCONNECTED_666, SV2V_UNCONNECTED_667, SV2V_UNCONNECTED_668, SV2V_UNCONNECTED_669, SV2V_UNCONNECTED_670, SV2V_UNCONNECTED_671, SV2V_UNCONNECTED_672, SV2V_UNCONNECTED_673, SV2V_UNCONNECTED_674, SV2V_UNCONNECTED_675, SV2V_UNCONNECTED_676, SV2V_UNCONNECTED_677, SV2V_UNCONNECTED_678, SV2V_UNCONNECTED_679, SV2V_UNCONNECTED_680, SV2V_UNCONNECTED_681, SV2V_UNCONNECTED_682, SV2V_UNCONNECTED_683, SV2V_UNCONNECTED_684, SV2V_UNCONNECTED_685, SV2V_UNCONNECTED_686, SV2V_UNCONNECTED_687, SV2V_UNCONNECTED_688, SV2V_UNCONNECTED_689, SV2V_UNCONNECTED_690, SV2V_UNCONNECTED_691, SV2V_UNCONNECTED_692, SV2V_UNCONNECTED_693, SV2V_UNCONNECTED_694, SV2V_UNCONNECTED_695, SV2V_UNCONNECTED_696, SV2V_UNCONNECTED_697, SV2V_UNCONNECTED_698, SV2V_UNCONNECTED_699, SV2V_UNCONNECTED_700, SV2V_UNCONNECTED_701, SV2V_UNCONNECTED_702, SV2V_UNCONNECTED_703, SV2V_UNCONNECTED_704, SV2V_UNCONNECTED_705, SV2V_UNCONNECTED_706, SV2V_UNCONNECTED_707, SV2V_UNCONNECTED_708, SV2V_UNCONNECTED_709, SV2V_UNCONNECTED_710, SV2V_UNCONNECTED_711, SV2V_UNCONNECTED_712, SV2V_UNCONNECTED_713, SV2V_UNCONNECTED_714, SV2V_UNCONNECTED_715, SV2V_UNCONNECTED_716, SV2V_UNCONNECTED_717, SV2V_UNCONNECTED_718, SV2V_UNCONNECTED_719, SV2V_UNCONNECTED_720, SV2V_UNCONNECTED_721, SV2V_UNCONNECTED_722, SV2V_UNCONNECTED_723, SV2V_UNCONNECTED_724, SV2V_UNCONNECTED_725, SV2V_UNCONNECTED_726, SV2V_UNCONNECTED_727, SV2V_UNCONNECTED_728, SV2V_UNCONNECTED_729, SV2V_UNCONNECTED_730, SV2V_UNCONNECTED_731, SV2V_UNCONNECTED_732, SV2V_UNCONNECTED_733, SV2V_UNCONNECTED_734, SV2V_UNCONNECTED_735, SV2V_UNCONNECTED_736, SV2V_UNCONNECTED_737, SV2V_UNCONNECTED_738, SV2V_UNCONNECTED_739, SV2V_UNCONNECTED_740, SV2V_UNCONNECTED_741, SV2V_UNCONNECTED_742, SV2V_UNCONNECTED_743, SV2V_UNCONNECTED_744, SV2V_UNCONNECTED_745, SV2V_UNCONNECTED_746, SV2V_UNCONNECTED_747, SV2V_UNCONNECTED_748, SV2V_UNCONNECTED_749, SV2V_UNCONNECTED_750, SV2V_UNCONNECTED_751, SV2V_UNCONNECTED_752, SV2V_UNCONNECTED_753, SV2V_UNCONNECTED_754, SV2V_UNCONNECTED_755, SV2V_UNCONNECTED_756, SV2V_UNCONNECTED_757, SV2V_UNCONNECTED_758, SV2V_UNCONNECTED_759, SV2V_UNCONNECTED_760, SV2V_UNCONNECTED_761, SV2V_UNCONNECTED_762, SV2V_UNCONNECTED_763, SV2V_UNCONNECTED_764, SV2V_UNCONNECTED_765, SV2V_UNCONNECTED_766, SV2V_UNCONNECTED_767, SV2V_UNCONNECTED_768, SV2V_UNCONNECTED_769, SV2V_UNCONNECTED_770, SV2V_UNCONNECTED_771, SV2V_UNCONNECTED_772, SV2V_UNCONNECTED_773, SV2V_UNCONNECTED_774, SV2V_UNCONNECTED_775, SV2V_UNCONNECTED_776, SV2V_UNCONNECTED_777, SV2V_UNCONNECTED_778, SV2V_UNCONNECTED_779, SV2V_UNCONNECTED_780, SV2V_UNCONNECTED_781, SV2V_UNCONNECTED_782, SV2V_UNCONNECTED_783, SV2V_UNCONNECTED_784, SV2V_UNCONNECTED_785, SV2V_UNCONNECTED_786, SV2V_UNCONNECTED_787, SV2V_UNCONNECTED_788, SV2V_UNCONNECTED_789, SV2V_UNCONNECTED_790, SV2V_UNCONNECTED_791, SV2V_UNCONNECTED_792, SV2V_UNCONNECTED_793, SV2V_UNCONNECTED_794, SV2V_UNCONNECTED_795, SV2V_UNCONNECTED_796, SV2V_UNCONNECTED_797, SV2V_UNCONNECTED_798, SV2V_UNCONNECTED_799, SV2V_UNCONNECTED_800, SV2V_UNCONNECTED_801, SV2V_UNCONNECTED_802, SV2V_UNCONNECTED_803, SV2V_UNCONNECTED_804, SV2V_UNCONNECTED_805, SV2V_UNCONNECTED_806, SV2V_UNCONNECTED_807, SV2V_UNCONNECTED_808, SV2V_UNCONNECTED_809, SV2V_UNCONNECTED_810, SV2V_UNCONNECTED_811, SV2V_UNCONNECTED_812, SV2V_UNCONNECTED_813, SV2V_UNCONNECTED_814, SV2V_UNCONNECTED_815, SV2V_UNCONNECTED_816, SV2V_UNCONNECTED_817, SV2V_UNCONNECTED_818, SV2V_UNCONNECTED_819, SV2V_UNCONNECTED_820, SV2V_UNCONNECTED_821, SV2V_UNCONNECTED_822, SV2V_UNCONNECTED_823, SV2V_UNCONNECTED_824, SV2V_UNCONNECTED_825, SV2V_UNCONNECTED_826, SV2V_UNCONNECTED_827, SV2V_UNCONNECTED_828, SV2V_UNCONNECTED_829, SV2V_UNCONNECTED_830, SV2V_UNCONNECTED_831, SV2V_UNCONNECTED_832, SV2V_UNCONNECTED_833, SV2V_UNCONNECTED_834, SV2V_UNCONNECTED_835, SV2V_UNCONNECTED_836, SV2V_UNCONNECTED_837, SV2V_UNCONNECTED_838, SV2V_UNCONNECTED_839, SV2V_UNCONNECTED_840, SV2V_UNCONNECTED_841, SV2V_UNCONNECTED_842, SV2V_UNCONNECTED_843, SV2V_UNCONNECTED_844, SV2V_UNCONNECTED_845, SV2V_UNCONNECTED_846, SV2V_UNCONNECTED_847, SV2V_UNCONNECTED_848, SV2V_UNCONNECTED_849, SV2V_UNCONNECTED_850, SV2V_UNCONNECTED_851, SV2V_UNCONNECTED_852, SV2V_UNCONNECTED_853, SV2V_UNCONNECTED_854, SV2V_UNCONNECTED_855, SV2V_UNCONNECTED_856, SV2V_UNCONNECTED_857, SV2V_UNCONNECTED_858, SV2V_UNCONNECTED_859, SV2V_UNCONNECTED_860, SV2V_UNCONNECTED_861, SV2V_UNCONNECTED_862, SV2V_UNCONNECTED_863, SV2V_UNCONNECTED_864, SV2V_UNCONNECTED_865, SV2V_UNCONNECTED_866, SV2V_UNCONNECTED_867, SV2V_UNCONNECTED_868, SV2V_UNCONNECTED_869, SV2V_UNCONNECTED_870, SV2V_UNCONNECTED_871, SV2V_UNCONNECTED_872, SV2V_UNCONNECTED_873, SV2V_UNCONNECTED_874, SV2V_UNCONNECTED_875, SV2V_UNCONNECTED_876, SV2V_UNCONNECTED_877, SV2V_UNCONNECTED_878, SV2V_UNCONNECTED_879, SV2V_UNCONNECTED_880, SV2V_UNCONNECTED_881, SV2V_UNCONNECTED_882, SV2V_UNCONNECTED_883, SV2V_UNCONNECTED_884, SV2V_UNCONNECTED_885, SV2V_UNCONNECTED_886, SV2V_UNCONNECTED_887, SV2V_UNCONNECTED_888, SV2V_UNCONNECTED_889, SV2V_UNCONNECTED_890, SV2V_UNCONNECTED_891, SV2V_UNCONNECTED_892, SV2V_UNCONNECTED_893, SV2V_UNCONNECTED_894, SV2V_UNCONNECTED_895, SV2V_UNCONNECTED_896, SV2V_UNCONNECTED_897, SV2V_UNCONNECTED_898, SV2V_UNCONNECTED_899, SV2V_UNCONNECTED_900, SV2V_UNCONNECTED_901, SV2V_UNCONNECTED_902, SV2V_UNCONNECTED_903, SV2V_UNCONNECTED_904, SV2V_UNCONNECTED_905, SV2V_UNCONNECTED_906, SV2V_UNCONNECTED_907, SV2V_UNCONNECTED_908, SV2V_UNCONNECTED_909, SV2V_UNCONNECTED_910, SV2V_UNCONNECTED_911, SV2V_UNCONNECTED_912, SV2V_UNCONNECTED_913, SV2V_UNCONNECTED_914, SV2V_UNCONNECTED_915, SV2V_UNCONNECTED_916, SV2V_UNCONNECTED_917, SV2V_UNCONNECTED_918, SV2V_UNCONNECTED_919, SV2V_UNCONNECTED_920, SV2V_UNCONNECTED_921, SV2V_UNCONNECTED_922, SV2V_UNCONNECTED_923, SV2V_UNCONNECTED_924, SV2V_UNCONNECTED_925, SV2V_UNCONNECTED_926, SV2V_UNCONNECTED_927, SV2V_UNCONNECTED_928, SV2V_UNCONNECTED_929, SV2V_UNCONNECTED_930, SV2V_UNCONNECTED_931, SV2V_UNCONNECTED_932, SV2V_UNCONNECTED_933, SV2V_UNCONNECTED_934, SV2V_UNCONNECTED_935, SV2V_UNCONNECTED_936, SV2V_UNCONNECTED_937, SV2V_UNCONNECTED_938, SV2V_UNCONNECTED_939, SV2V_UNCONNECTED_940, SV2V_UNCONNECTED_941, SV2V_UNCONNECTED_942, SV2V_UNCONNECTED_943, SV2V_UNCONNECTED_944, SV2V_UNCONNECTED_945, SV2V_UNCONNECTED_946, SV2V_UNCONNECTED_947, SV2V_UNCONNECTED_948, SV2V_UNCONNECTED_949, SV2V_UNCONNECTED_950, SV2V_UNCONNECTED_951, SV2V_UNCONNECTED_952, SV2V_UNCONNECTED_953, SV2V_UNCONNECTED_954, SV2V_UNCONNECTED_955, SV2V_UNCONNECTED_956, SV2V_UNCONNECTED_957, SV2V_UNCONNECTED_958, SV2V_UNCONNECTED_959, SV2V_UNCONNECTED_960, SV2V_UNCONNECTED_961, SV2V_UNCONNECTED_962, SV2V_UNCONNECTED_963, SV2V_UNCONNECTED_964, SV2V_UNCONNECTED_965, SV2V_UNCONNECTED_966, SV2V_UNCONNECTED_967, SV2V_UNCONNECTED_968, SV2V_UNCONNECTED_969, SV2V_UNCONNECTED_970, SV2V_UNCONNECTED_971, SV2V_UNCONNECTED_972, SV2V_UNCONNECTED_973, SV2V_UNCONNECTED_974, SV2V_UNCONNECTED_975, SV2V_UNCONNECTED_976, SV2V_UNCONNECTED_977, SV2V_UNCONNECTED_978, SV2V_UNCONNECTED_979, SV2V_UNCONNECTED_980, SV2V_UNCONNECTED_981, SV2V_UNCONNECTED_982, SV2V_UNCONNECTED_983, SV2V_UNCONNECTED_984, SV2V_UNCONNECTED_985, SV2V_UNCONNECTED_986, SV2V_UNCONNECTED_987, SV2V_UNCONNECTED_988, SV2V_UNCONNECTED_989, SV2V_UNCONNECTED_990, SV2V_UNCONNECTED_991, SV2V_UNCONNECTED_992, SV2V_UNCONNECTED_993, SV2V_UNCONNECTED_994, SV2V_UNCONNECTED_995, SV2V_UNCONNECTED_996, SV2V_UNCONNECTED_997, SV2V_UNCONNECTED_998, SV2V_UNCONNECTED_999, SV2V_UNCONNECTED_1000, SV2V_UNCONNECTED_1001, SV2V_UNCONNECTED_1002, SV2V_UNCONNECTED_1003, SV2V_UNCONNECTED_1004, SV2V_UNCONNECTED_1005, SV2V_UNCONNECTED_1006, SV2V_UNCONNECTED_1007, SV2V_UNCONNECTED_1008, SV2V_UNCONNECTED_1009, SV2V_UNCONNECTED_1010, SV2V_UNCONNECTED_1011, SV2V_UNCONNECTED_1012, SV2V_UNCONNECTED_1013, SV2V_UNCONNECTED_1014, SV2V_UNCONNECTED_1015, SV2V_UNCONNECTED_1016, SV2V_UNCONNECTED_1017, SV2V_UNCONNECTED_1018, SV2V_UNCONNECTED_1019, SV2V_UNCONNECTED_1020, SV2V_UNCONNECTED_1021, SV2V_UNCONNECTED_1022, SV2V_UNCONNECTED_1023, SV2V_UNCONNECTED_1024, SV2V_UNCONNECTED_1025, SV2V_UNCONNECTED_1026, SV2V_UNCONNECTED_1027, SV2V_UNCONNECTED_1028, SV2V_UNCONNECTED_1029, SV2V_UNCONNECTED_1030, SV2V_UNCONNECTED_1031, SV2V_UNCONNECTED_1032, SV2V_UNCONNECTED_1033, SV2V_UNCONNECTED_1034, SV2V_UNCONNECTED_1035, SV2V_UNCONNECTED_1036, SV2V_UNCONNECTED_1037, SV2V_UNCONNECTED_1038, SV2V_UNCONNECTED_1039, SV2V_UNCONNECTED_1040, SV2V_UNCONNECTED_1041, SV2V_UNCONNECTED_1042, SV2V_UNCONNECTED_1043, SV2V_UNCONNECTED_1044, SV2V_UNCONNECTED_1045, SV2V_UNCONNECTED_1046, SV2V_UNCONNECTED_1047, SV2V_UNCONNECTED_1048, SV2V_UNCONNECTED_1049, SV2V_UNCONNECTED_1050, SV2V_UNCONNECTED_1051, SV2V_UNCONNECTED_1052, SV2V_UNCONNECTED_1053, SV2V_UNCONNECTED_1054, SV2V_UNCONNECTED_1055, SV2V_UNCONNECTED_1056, SV2V_UNCONNECTED_1057, SV2V_UNCONNECTED_1058, SV2V_UNCONNECTED_1059, SV2V_UNCONNECTED_1060, SV2V_UNCONNECTED_1061, SV2V_UNCONNECTED_1062, SV2V_UNCONNECTED_1063, SV2V_UNCONNECTED_1064, SV2V_UNCONNECTED_1065, SV2V_UNCONNECTED_1066, SV2V_UNCONNECTED_1067, SV2V_UNCONNECTED_1068, SV2V_UNCONNECTED_1069, SV2V_UNCONNECTED_1070, SV2V_UNCONNECTED_1071, SV2V_UNCONNECTED_1072, SV2V_UNCONNECTED_1073, SV2V_UNCONNECTED_1074, SV2V_UNCONNECTED_1075, SV2V_UNCONNECTED_1076, SV2V_UNCONNECTED_1077, SV2V_UNCONNECTED_1078, SV2V_UNCONNECTED_1079, SV2V_UNCONNECTED_1080, SV2V_UNCONNECTED_1081, SV2V_UNCONNECTED_1082, SV2V_UNCONNECTED_1083, SV2V_UNCONNECTED_1084, SV2V_UNCONNECTED_1085, SV2V_UNCONNECTED_1086, SV2V_UNCONNECTED_1087, SV2V_UNCONNECTED_1088, SV2V_UNCONNECTED_1089, SV2V_UNCONNECTED_1090, SV2V_UNCONNECTED_1091, SV2V_UNCONNECTED_1092, SV2V_UNCONNECTED_1093, SV2V_UNCONNECTED_1094, SV2V_UNCONNECTED_1095, SV2V_UNCONNECTED_1096, SV2V_UNCONNECTED_1097, SV2V_UNCONNECTED_1098, SV2V_UNCONNECTED_1099, SV2V_UNCONNECTED_1100, SV2V_UNCONNECTED_1101, SV2V_UNCONNECTED_1102, SV2V_UNCONNECTED_1103, SV2V_UNCONNECTED_1104, SV2V_UNCONNECTED_1105, SV2V_UNCONNECTED_1106, SV2V_UNCONNECTED_1107, SV2V_UNCONNECTED_1108, SV2V_UNCONNECTED_1109, SV2V_UNCONNECTED_1110, SV2V_UNCONNECTED_1111, SV2V_UNCONNECTED_1112, SV2V_UNCONNECTED_1113, SV2V_UNCONNECTED_1114, SV2V_UNCONNECTED_1115, SV2V_UNCONNECTED_1116, SV2V_UNCONNECTED_1117, SV2V_UNCONNECTED_1118, SV2V_UNCONNECTED_1119, SV2V_UNCONNECTED_1120, SV2V_UNCONNECTED_1121, SV2V_UNCONNECTED_1122, SV2V_UNCONNECTED_1123, SV2V_UNCONNECTED_1124, SV2V_UNCONNECTED_1125, SV2V_UNCONNECTED_1126, SV2V_UNCONNECTED_1127, SV2V_UNCONNECTED_1128, SV2V_UNCONNECTED_1129, SV2V_UNCONNECTED_1130, SV2V_UNCONNECTED_1131, SV2V_UNCONNECTED_1132, SV2V_UNCONNECTED_1133, SV2V_UNCONNECTED_1134, SV2V_UNCONNECTED_1135, SV2V_UNCONNECTED_1136, SV2V_UNCONNECTED_1137, SV2V_UNCONNECTED_1138, SV2V_UNCONNECTED_1139, SV2V_UNCONNECTED_1140, SV2V_UNCONNECTED_1141, SV2V_UNCONNECTED_1142, SV2V_UNCONNECTED_1143, SV2V_UNCONNECTED_1144, SV2V_UNCONNECTED_1145, SV2V_UNCONNECTED_1146, SV2V_UNCONNECTED_1147, SV2V_UNCONNECTED_1148, SV2V_UNCONNECTED_1149, SV2V_UNCONNECTED_1150, SV2V_UNCONNECTED_1151, SV2V_UNCONNECTED_1152, SV2V_UNCONNECTED_1153, SV2V_UNCONNECTED_1154, SV2V_UNCONNECTED_1155, SV2V_UNCONNECTED_1156, SV2V_UNCONNECTED_1157, SV2V_UNCONNECTED_1158, SV2V_UNCONNECTED_1159, SV2V_UNCONNECTED_1160, SV2V_UNCONNECTED_1161, SV2V_UNCONNECTED_1162, SV2V_UNCONNECTED_1163, SV2V_UNCONNECTED_1164, SV2V_UNCONNECTED_1165, SV2V_UNCONNECTED_1166, SV2V_UNCONNECTED_1167, SV2V_UNCONNECTED_1168, SV2V_UNCONNECTED_1169, SV2V_UNCONNECTED_1170, SV2V_UNCONNECTED_1171, SV2V_UNCONNECTED_1172, SV2V_UNCONNECTED_1173, SV2V_UNCONNECTED_1174, SV2V_UNCONNECTED_1175, SV2V_UNCONNECTED_1176, SV2V_UNCONNECTED_1177, SV2V_UNCONNECTED_1178, SV2V_UNCONNECTED_1179, SV2V_UNCONNECTED_1180, SV2V_UNCONNECTED_1181, SV2V_UNCONNECTED_1182, SV2V_UNCONNECTED_1183, SV2V_UNCONNECTED_1184, SV2V_UNCONNECTED_1185, SV2V_UNCONNECTED_1186, SV2V_UNCONNECTED_1187, SV2V_UNCONNECTED_1188, SV2V_UNCONNECTED_1189, SV2V_UNCONNECTED_1190, SV2V_UNCONNECTED_1191, SV2V_UNCONNECTED_1192, SV2V_UNCONNECTED_1193, SV2V_UNCONNECTED_1194, SV2V_UNCONNECTED_1195, SV2V_UNCONNECTED_1196, SV2V_UNCONNECTED_1197, SV2V_UNCONNECTED_1198, SV2V_UNCONNECTED_1199, SV2V_UNCONNECTED_1200, SV2V_UNCONNECTED_1201, SV2V_UNCONNECTED_1202, SV2V_UNCONNECTED_1203, SV2V_UNCONNECTED_1204, SV2V_UNCONNECTED_1205, SV2V_UNCONNECTED_1206, SV2V_UNCONNECTED_1207, SV2V_UNCONNECTED_1208, SV2V_UNCONNECTED_1209, SV2V_UNCONNECTED_1210, SV2V_UNCONNECTED_1211, SV2V_UNCONNECTED_1212, SV2V_UNCONNECTED_1213, SV2V_UNCONNECTED_1214, SV2V_UNCONNECTED_1215, SV2V_UNCONNECTED_1216, SV2V_UNCONNECTED_1217, SV2V_UNCONNECTED_1218, SV2V_UNCONNECTED_1219, SV2V_UNCONNECTED_1220, SV2V_UNCONNECTED_1221, SV2V_UNCONNECTED_1222, SV2V_UNCONNECTED_1223, SV2V_UNCONNECTED_1224, SV2V_UNCONNECTED_1225, SV2V_UNCONNECTED_1226, SV2V_UNCONNECTED_1227, SV2V_UNCONNECTED_1228, SV2V_UNCONNECTED_1229, SV2V_UNCONNECTED_1230, SV2V_UNCONNECTED_1231, SV2V_UNCONNECTED_1232, SV2V_UNCONNECTED_1233, SV2V_UNCONNECTED_1234, SV2V_UNCONNECTED_1235, SV2V_UNCONNECTED_1236, SV2V_UNCONNECTED_1237, SV2V_UNCONNECTED_1238, SV2V_UNCONNECTED_1239, SV2V_UNCONNECTED_1240, SV2V_UNCONNECTED_1241, SV2V_UNCONNECTED_1242, SV2V_UNCONNECTED_1243, SV2V_UNCONNECTED_1244, SV2V_UNCONNECTED_1245, SV2V_UNCONNECTED_1246, SV2V_UNCONNECTED_1247, SV2V_UNCONNECTED_1248, SV2V_UNCONNECTED_1249, SV2V_UNCONNECTED_1250, SV2V_UNCONNECTED_1251, SV2V_UNCONNECTED_1252, SV2V_UNCONNECTED_1253, SV2V_UNCONNECTED_1254, SV2V_UNCONNECTED_1255, SV2V_UNCONNECTED_1256, SV2V_UNCONNECTED_1257, SV2V_UNCONNECTED_1258, SV2V_UNCONNECTED_1259, SV2V_UNCONNECTED_1260, SV2V_UNCONNECTED_1261, SV2V_UNCONNECTED_1262, SV2V_UNCONNECTED_1263, SV2V_UNCONNECTED_1264, SV2V_UNCONNECTED_1265, SV2V_UNCONNECTED_1266, SV2V_UNCONNECTED_1267, SV2V_UNCONNECTED_1268, SV2V_UNCONNECTED_1269, SV2V_UNCONNECTED_1270, SV2V_UNCONNECTED_1271, SV2V_UNCONNECTED_1272, SV2V_UNCONNECTED_1273, SV2V_UNCONNECTED_1274, SV2V_UNCONNECTED_1275, SV2V_UNCONNECTED_1276, SV2V_UNCONNECTED_1277, SV2V_UNCONNECTED_1278, SV2V_UNCONNECTED_1279, SV2V_UNCONNECTED_1280, SV2V_UNCONNECTED_1281, SV2V_UNCONNECTED_1282, SV2V_UNCONNECTED_1283, SV2V_UNCONNECTED_1284, SV2V_UNCONNECTED_1285, SV2V_UNCONNECTED_1286, SV2V_UNCONNECTED_1287, SV2V_UNCONNECTED_1288, SV2V_UNCONNECTED_1289, SV2V_UNCONNECTED_1290, SV2V_UNCONNECTED_1291, SV2V_UNCONNECTED_1292, SV2V_UNCONNECTED_1293, SV2V_UNCONNECTED_1294, SV2V_UNCONNECTED_1295, SV2V_UNCONNECTED_1296, SV2V_UNCONNECTED_1297, SV2V_UNCONNECTED_1298, SV2V_UNCONNECTED_1299, SV2V_UNCONNECTED_1300, SV2V_UNCONNECTED_1301, SV2V_UNCONNECTED_1302, SV2V_UNCONNECTED_1303, SV2V_UNCONNECTED_1304, SV2V_UNCONNECTED_1305, SV2V_UNCONNECTED_1306, SV2V_UNCONNECTED_1307, SV2V_UNCONNECTED_1308, SV2V_UNCONNECTED_1309, SV2V_UNCONNECTED_1310, SV2V_UNCONNECTED_1311, SV2V_UNCONNECTED_1312, SV2V_UNCONNECTED_1313, SV2V_UNCONNECTED_1314, SV2V_UNCONNECTED_1315, SV2V_UNCONNECTED_1316, SV2V_UNCONNECTED_1317, SV2V_UNCONNECTED_1318, SV2V_UNCONNECTED_1319, SV2V_UNCONNECTED_1320, SV2V_UNCONNECTED_1321, SV2V_UNCONNECTED_1322, SV2V_UNCONNECTED_1323, SV2V_UNCONNECTED_1324, SV2V_UNCONNECTED_1325, SV2V_UNCONNECTED_1326, SV2V_UNCONNECTED_1327, SV2V_UNCONNECTED_1328, SV2V_UNCONNECTED_1329, SV2V_UNCONNECTED_1330, SV2V_UNCONNECTED_1331, SV2V_UNCONNECTED_1332, SV2V_UNCONNECTED_1333, SV2V_UNCONNECTED_1334, SV2V_UNCONNECTED_1335, SV2V_UNCONNECTED_1336, SV2V_UNCONNECTED_1337, SV2V_UNCONNECTED_1338, SV2V_UNCONNECTED_1339, SV2V_UNCONNECTED_1340, SV2V_UNCONNECTED_1341, SV2V_UNCONNECTED_1342, SV2V_UNCONNECTED_1343, SV2V_UNCONNECTED_1344, SV2V_UNCONNECTED_1345, SV2V_UNCONNECTED_1346, SV2V_UNCONNECTED_1347, SV2V_UNCONNECTED_1348, SV2V_UNCONNECTED_1349, SV2V_UNCONNECTED_1350, SV2V_UNCONNECTED_1351, SV2V_UNCONNECTED_1352, SV2V_UNCONNECTED_1353, SV2V_UNCONNECTED_1354, SV2V_UNCONNECTED_1355, SV2V_UNCONNECTED_1356, SV2V_UNCONNECTED_1357, SV2V_UNCONNECTED_1358, SV2V_UNCONNECTED_1359, SV2V_UNCONNECTED_1360, SV2V_UNCONNECTED_1361, SV2V_UNCONNECTED_1362, SV2V_UNCONNECTED_1363, SV2V_UNCONNECTED_1364, SV2V_UNCONNECTED_1365, SV2V_UNCONNECTED_1366, SV2V_UNCONNECTED_1367, SV2V_UNCONNECTED_1368, SV2V_UNCONNECTED_1369, SV2V_UNCONNECTED_1370, SV2V_UNCONNECTED_1371, SV2V_UNCONNECTED_1372, SV2V_UNCONNECTED_1373, SV2V_UNCONNECTED_1374, SV2V_UNCONNECTED_1375, SV2V_UNCONNECTED_1376, SV2V_UNCONNECTED_1377, SV2V_UNCONNECTED_1378, SV2V_UNCONNECTED_1379, SV2V_UNCONNECTED_1380, SV2V_UNCONNECTED_1381, SV2V_UNCONNECTED_1382, SV2V_UNCONNECTED_1383, SV2V_UNCONNECTED_1384, SV2V_UNCONNECTED_1385, SV2V_UNCONNECTED_1386, SV2V_UNCONNECTED_1387, SV2V_UNCONNECTED_1388, SV2V_UNCONNECTED_1389, SV2V_UNCONNECTED_1390, SV2V_UNCONNECTED_1391, SV2V_UNCONNECTED_1392, SV2V_UNCONNECTED_1393, SV2V_UNCONNECTED_1394, SV2V_UNCONNECTED_1395, SV2V_UNCONNECTED_1396, SV2V_UNCONNECTED_1397, SV2V_UNCONNECTED_1398, SV2V_UNCONNECTED_1399, SV2V_UNCONNECTED_1400, SV2V_UNCONNECTED_1401, SV2V_UNCONNECTED_1402, SV2V_UNCONNECTED_1403, SV2V_UNCONNECTED_1404, SV2V_UNCONNECTED_1405, SV2V_UNCONNECTED_1406, SV2V_UNCONNECTED_1407, SV2V_UNCONNECTED_1408, SV2V_UNCONNECTED_1409, SV2V_UNCONNECTED_1410, SV2V_UNCONNECTED_1411, SV2V_UNCONNECTED_1412, SV2V_UNCONNECTED_1413, SV2V_UNCONNECTED_1414, SV2V_UNCONNECTED_1415, SV2V_UNCONNECTED_1416, SV2V_UNCONNECTED_1417, SV2V_UNCONNECTED_1418, SV2V_UNCONNECTED_1419, SV2V_UNCONNECTED_1420, SV2V_UNCONNECTED_1421, SV2V_UNCONNECTED_1422, SV2V_UNCONNECTED_1423, SV2V_UNCONNECTED_1424, SV2V_UNCONNECTED_1425, SV2V_UNCONNECTED_1426, SV2V_UNCONNECTED_1427, SV2V_UNCONNECTED_1428, SV2V_UNCONNECTED_1429, SV2V_UNCONNECTED_1430, SV2V_UNCONNECTED_1431, SV2V_UNCONNECTED_1432, SV2V_UNCONNECTED_1433, SV2V_UNCONNECTED_1434, SV2V_UNCONNECTED_1435, SV2V_UNCONNECTED_1436, SV2V_UNCONNECTED_1437, SV2V_UNCONNECTED_1438, SV2V_UNCONNECTED_1439, SV2V_UNCONNECTED_1440, SV2V_UNCONNECTED_1441, SV2V_UNCONNECTED_1442, SV2V_UNCONNECTED_1443, SV2V_UNCONNECTED_1444, SV2V_UNCONNECTED_1445, SV2V_UNCONNECTED_1446, SV2V_UNCONNECTED_1447, SV2V_UNCONNECTED_1448, SV2V_UNCONNECTED_1449, SV2V_UNCONNECTED_1450, SV2V_UNCONNECTED_1451, SV2V_UNCONNECTED_1452, SV2V_UNCONNECTED_1453, SV2V_UNCONNECTED_1454, SV2V_UNCONNECTED_1455, SV2V_UNCONNECTED_1456, SV2V_UNCONNECTED_1457, SV2V_UNCONNECTED_1458, SV2V_UNCONNECTED_1459, SV2V_UNCONNECTED_1460, SV2V_UNCONNECTED_1461, SV2V_UNCONNECTED_1462, SV2V_UNCONNECTED_1463, SV2V_UNCONNECTED_1464, SV2V_UNCONNECTED_1465, SV2V_UNCONNECTED_1466, SV2V_UNCONNECTED_1467, SV2V_UNCONNECTED_1468, SV2V_UNCONNECTED_1469, SV2V_UNCONNECTED_1470, SV2V_UNCONNECTED_1471, SV2V_UNCONNECTED_1472, SV2V_UNCONNECTED_1473, SV2V_UNCONNECTED_1474, SV2V_UNCONNECTED_1475, SV2V_UNCONNECTED_1476, SV2V_UNCONNECTED_1477, SV2V_UNCONNECTED_1478, SV2V_UNCONNECTED_1479, SV2V_UNCONNECTED_1480, SV2V_UNCONNECTED_1481, SV2V_UNCONNECTED_1482, SV2V_UNCONNECTED_1483, SV2V_UNCONNECTED_1484, SV2V_UNCONNECTED_1485, SV2V_UNCONNECTED_1486, SV2V_UNCONNECTED_1487, SV2V_UNCONNECTED_1488, SV2V_UNCONNECTED_1489, SV2V_UNCONNECTED_1490, SV2V_UNCONNECTED_1491, SV2V_UNCONNECTED_1492, SV2V_UNCONNECTED_1493, SV2V_UNCONNECTED_1494, SV2V_UNCONNECTED_1495, SV2V_UNCONNECTED_1496, SV2V_UNCONNECTED_1497, SV2V_UNCONNECTED_1498, SV2V_UNCONNECTED_1499, SV2V_UNCONNECTED_1500, SV2V_UNCONNECTED_1501, SV2V_UNCONNECTED_1502, SV2V_UNCONNECTED_1503, SV2V_UNCONNECTED_1504, SV2V_UNCONNECTED_1505, SV2V_UNCONNECTED_1506, SV2V_UNCONNECTED_1507, SV2V_UNCONNECTED_1508, SV2V_UNCONNECTED_1509, SV2V_UNCONNECTED_1510, SV2V_UNCONNECTED_1511, SV2V_UNCONNECTED_1512, SV2V_UNCONNECTED_1513, SV2V_UNCONNECTED_1514, SV2V_UNCONNECTED_1515, SV2V_UNCONNECTED_1516, SV2V_UNCONNECTED_1517, SV2V_UNCONNECTED_1518, SV2V_UNCONNECTED_1519, SV2V_UNCONNECTED_1520, SV2V_UNCONNECTED_1521, SV2V_UNCONNECTED_1522, SV2V_UNCONNECTED_1523, SV2V_UNCONNECTED_1524, SV2V_UNCONNECTED_1525, SV2V_UNCONNECTED_1526, SV2V_UNCONNECTED_1527, SV2V_UNCONNECTED_1528, SV2V_UNCONNECTED_1529, SV2V_UNCONNECTED_1530, SV2V_UNCONNECTED_1531, SV2V_UNCONNECTED_1532, SV2V_UNCONNECTED_1533, SV2V_UNCONNECTED_1534, SV2V_UNCONNECTED_1535, SV2V_UNCONNECTED_1536, SV2V_UNCONNECTED_1537, SV2V_UNCONNECTED_1538, SV2V_UNCONNECTED_1539, SV2V_UNCONNECTED_1540, SV2V_UNCONNECTED_1541, SV2V_UNCONNECTED_1542, SV2V_UNCONNECTED_1543, SV2V_UNCONNECTED_1544, SV2V_UNCONNECTED_1545, SV2V_UNCONNECTED_1546, SV2V_UNCONNECTED_1547, SV2V_UNCONNECTED_1548, SV2V_UNCONNECTED_1549, SV2V_UNCONNECTED_1550, SV2V_UNCONNECTED_1551, SV2V_UNCONNECTED_1552, SV2V_UNCONNECTED_1553, SV2V_UNCONNECTED_1554, SV2V_UNCONNECTED_1555, SV2V_UNCONNECTED_1556, SV2V_UNCONNECTED_1557, SV2V_UNCONNECTED_1558, SV2V_UNCONNECTED_1559, SV2V_UNCONNECTED_1560, SV2V_UNCONNECTED_1561, SV2V_UNCONNECTED_1562, SV2V_UNCONNECTED_1563, SV2V_UNCONNECTED_1564, SV2V_UNCONNECTED_1565, SV2V_UNCONNECTED_1566, SV2V_UNCONNECTED_1567, SV2V_UNCONNECTED_1568, SV2V_UNCONNECTED_1569, SV2V_UNCONNECTED_1570, SV2V_UNCONNECTED_1571, SV2V_UNCONNECTED_1572, SV2V_UNCONNECTED_1573, SV2V_UNCONNECTED_1574, SV2V_UNCONNECTED_1575, SV2V_UNCONNECTED_1576, SV2V_UNCONNECTED_1577, SV2V_UNCONNECTED_1578, SV2V_UNCONNECTED_1579, SV2V_UNCONNECTED_1580, SV2V_UNCONNECTED_1581, SV2V_UNCONNECTED_1582, SV2V_UNCONNECTED_1583, SV2V_UNCONNECTED_1584, SV2V_UNCONNECTED_1585, SV2V_UNCONNECTED_1586, SV2V_UNCONNECTED_1587, SV2V_UNCONNECTED_1588, SV2V_UNCONNECTED_1589, SV2V_UNCONNECTED_1590, SV2V_UNCONNECTED_1591, SV2V_UNCONNECTED_1592, SV2V_UNCONNECTED_1593, SV2V_UNCONNECTED_1594, SV2V_UNCONNECTED_1595, SV2V_UNCONNECTED_1596, SV2V_UNCONNECTED_1597, SV2V_UNCONNECTED_1598, SV2V_UNCONNECTED_1599, SV2V_UNCONNECTED_1600, SV2V_UNCONNECTED_1601, SV2V_UNCONNECTED_1602, SV2V_UNCONNECTED_1603, SV2V_UNCONNECTED_1604, SV2V_UNCONNECTED_1605, SV2V_UNCONNECTED_1606, SV2V_UNCONNECTED_1607, SV2V_UNCONNECTED_1608, SV2V_UNCONNECTED_1609, SV2V_UNCONNECTED_1610, SV2V_UNCONNECTED_1611, SV2V_UNCONNECTED_1612, SV2V_UNCONNECTED_1613, SV2V_UNCONNECTED_1614, SV2V_UNCONNECTED_1615, SV2V_UNCONNECTED_1616, SV2V_UNCONNECTED_1617, SV2V_UNCONNECTED_1618, SV2V_UNCONNECTED_1619, SV2V_UNCONNECTED_1620, SV2V_UNCONNECTED_1621, SV2V_UNCONNECTED_1622, SV2V_UNCONNECTED_1623, SV2V_UNCONNECTED_1624, SV2V_UNCONNECTED_1625, SV2V_UNCONNECTED_1626, SV2V_UNCONNECTED_1627, SV2V_UNCONNECTED_1628, SV2V_UNCONNECTED_1629, SV2V_UNCONNECTED_1630, SV2V_UNCONNECTED_1631, SV2V_UNCONNECTED_1632, SV2V_UNCONNECTED_1633, SV2V_UNCONNECTED_1634, SV2V_UNCONNECTED_1635, SV2V_UNCONNECTED_1636, SV2V_UNCONNECTED_1637, SV2V_UNCONNECTED_1638, SV2V_UNCONNECTED_1639, SV2V_UNCONNECTED_1640, SV2V_UNCONNECTED_1641, SV2V_UNCONNECTED_1642, SV2V_UNCONNECTED_1643, SV2V_UNCONNECTED_1644, SV2V_UNCONNECTED_1645, SV2V_UNCONNECTED_1646, SV2V_UNCONNECTED_1647, SV2V_UNCONNECTED_1648, SV2V_UNCONNECTED_1649, SV2V_UNCONNECTED_1650, SV2V_UNCONNECTED_1651, SV2V_UNCONNECTED_1652, SV2V_UNCONNECTED_1653, SV2V_UNCONNECTED_1654, SV2V_UNCONNECTED_1655, SV2V_UNCONNECTED_1656, SV2V_UNCONNECTED_1657, SV2V_UNCONNECTED_1658, SV2V_UNCONNECTED_1659, SV2V_UNCONNECTED_1660, SV2V_UNCONNECTED_1661, SV2V_UNCONNECTED_1662, SV2V_UNCONNECTED_1663, SV2V_UNCONNECTED_1664, SV2V_UNCONNECTED_1665, SV2V_UNCONNECTED_1666, SV2V_UNCONNECTED_1667, SV2V_UNCONNECTED_1668, SV2V_UNCONNECTED_1669, SV2V_UNCONNECTED_1670, SV2V_UNCONNECTED_1671, SV2V_UNCONNECTED_1672, SV2V_UNCONNECTED_1673, SV2V_UNCONNECTED_1674, SV2V_UNCONNECTED_1675, SV2V_UNCONNECTED_1676, SV2V_UNCONNECTED_1677, SV2V_UNCONNECTED_1678, SV2V_UNCONNECTED_1679, SV2V_UNCONNECTED_1680, SV2V_UNCONNECTED_1681, SV2V_UNCONNECTED_1682, SV2V_UNCONNECTED_1683, SV2V_UNCONNECTED_1684, SV2V_UNCONNECTED_1685, SV2V_UNCONNECTED_1686, SV2V_UNCONNECTED_1687, SV2V_UNCONNECTED_1688, SV2V_UNCONNECTED_1689, SV2V_UNCONNECTED_1690, SV2V_UNCONNECTED_1691, SV2V_UNCONNECTED_1692, SV2V_UNCONNECTED_1693, SV2V_UNCONNECTED_1694, SV2V_UNCONNECTED_1695, SV2V_UNCONNECTED_1696, SV2V_UNCONNECTED_1697, SV2V_UNCONNECTED_1698, SV2V_UNCONNECTED_1699, SV2V_UNCONNECTED_1700, SV2V_UNCONNECTED_1701, SV2V_UNCONNECTED_1702, SV2V_UNCONNECTED_1703, SV2V_UNCONNECTED_1704, SV2V_UNCONNECTED_1705, SV2V_UNCONNECTED_1706, SV2V_UNCONNECTED_1707, SV2V_UNCONNECTED_1708, SV2V_UNCONNECTED_1709, SV2V_UNCONNECTED_1710, SV2V_UNCONNECTED_1711, SV2V_UNCONNECTED_1712, SV2V_UNCONNECTED_1713, SV2V_UNCONNECTED_1714, SV2V_UNCONNECTED_1715, SV2V_UNCONNECTED_1716, SV2V_UNCONNECTED_1717, SV2V_UNCONNECTED_1718, SV2V_UNCONNECTED_1719, SV2V_UNCONNECTED_1720, SV2V_UNCONNECTED_1721, SV2V_UNCONNECTED_1722, SV2V_UNCONNECTED_1723, SV2V_UNCONNECTED_1724, SV2V_UNCONNECTED_1725, SV2V_UNCONNECTED_1726, SV2V_UNCONNECTED_1727, SV2V_UNCONNECTED_1728, SV2V_UNCONNECTED_1729, SV2V_UNCONNECTED_1730, SV2V_UNCONNECTED_1731, SV2V_UNCONNECTED_1732, SV2V_UNCONNECTED_1733, SV2V_UNCONNECTED_1734, SV2V_UNCONNECTED_1735, SV2V_UNCONNECTED_1736, SV2V_UNCONNECTED_1737, SV2V_UNCONNECTED_1738, SV2V_UNCONNECTED_1739, SV2V_UNCONNECTED_1740, SV2V_UNCONNECTED_1741, SV2V_UNCONNECTED_1742, SV2V_UNCONNECTED_1743, SV2V_UNCONNECTED_1744, SV2V_UNCONNECTED_1745, SV2V_UNCONNECTED_1746, SV2V_UNCONNECTED_1747, SV2V_UNCONNECTED_1748, SV2V_UNCONNECTED_1749, SV2V_UNCONNECTED_1750, SV2V_UNCONNECTED_1751, SV2V_UNCONNECTED_1752, SV2V_UNCONNECTED_1753, SV2V_UNCONNECTED_1754, SV2V_UNCONNECTED_1755, SV2V_UNCONNECTED_1756, SV2V_UNCONNECTED_1757, SV2V_UNCONNECTED_1758, SV2V_UNCONNECTED_1759, SV2V_UNCONNECTED_1760, SV2V_UNCONNECTED_1761, SV2V_UNCONNECTED_1762, SV2V_UNCONNECTED_1763, SV2V_UNCONNECTED_1764, SV2V_UNCONNECTED_1765, SV2V_UNCONNECTED_1766, SV2V_UNCONNECTED_1767, SV2V_UNCONNECTED_1768, SV2V_UNCONNECTED_1769, SV2V_UNCONNECTED_1770, SV2V_UNCONNECTED_1771, SV2V_UNCONNECTED_1772, SV2V_UNCONNECTED_1773, SV2V_UNCONNECTED_1774, SV2V_UNCONNECTED_1775, SV2V_UNCONNECTED_1776, SV2V_UNCONNECTED_1777, SV2V_UNCONNECTED_1778, SV2V_UNCONNECTED_1779, SV2V_UNCONNECTED_1780, SV2V_UNCONNECTED_1781, SV2V_UNCONNECTED_1782, SV2V_UNCONNECTED_1783, SV2V_UNCONNECTED_1784, SV2V_UNCONNECTED_1785, SV2V_UNCONNECTED_1786, SV2V_UNCONNECTED_1787, SV2V_UNCONNECTED_1788, SV2V_UNCONNECTED_1789, SV2V_UNCONNECTED_1790, SV2V_UNCONNECTED_1791, SV2V_UNCONNECTED_1792, SV2V_UNCONNECTED_1793, SV2V_UNCONNECTED_1794, SV2V_UNCONNECTED_1795, SV2V_UNCONNECTED_1796, SV2V_UNCONNECTED_1797, SV2V_UNCONNECTED_1798, SV2V_UNCONNECTED_1799, SV2V_UNCONNECTED_1800, SV2V_UNCONNECTED_1801, SV2V_UNCONNECTED_1802, SV2V_UNCONNECTED_1803, SV2V_UNCONNECTED_1804, SV2V_UNCONNECTED_1805, SV2V_UNCONNECTED_1806, SV2V_UNCONNECTED_1807, SV2V_UNCONNECTED_1808, SV2V_UNCONNECTED_1809, SV2V_UNCONNECTED_1810, SV2V_UNCONNECTED_1811, SV2V_UNCONNECTED_1812, SV2V_UNCONNECTED_1813, SV2V_UNCONNECTED_1814, SV2V_UNCONNECTED_1815, SV2V_UNCONNECTED_1816, SV2V_UNCONNECTED_1817, SV2V_UNCONNECTED_1818, SV2V_UNCONNECTED_1819, SV2V_UNCONNECTED_1820, SV2V_UNCONNECTED_1821, SV2V_UNCONNECTED_1822, SV2V_UNCONNECTED_1823, SV2V_UNCONNECTED_1824, SV2V_UNCONNECTED_1825, SV2V_UNCONNECTED_1826, SV2V_UNCONNECTED_1827, SV2V_UNCONNECTED_1828, SV2V_UNCONNECTED_1829, SV2V_UNCONNECTED_1830, SV2V_UNCONNECTED_1831, SV2V_UNCONNECTED_1832, SV2V_UNCONNECTED_1833, SV2V_UNCONNECTED_1834, SV2V_UNCONNECTED_1835, SV2V_UNCONNECTED_1836, SV2V_UNCONNECTED_1837, SV2V_UNCONNECTED_1838, SV2V_UNCONNECTED_1839, SV2V_UNCONNECTED_1840, SV2V_UNCONNECTED_1841, SV2V_UNCONNECTED_1842, SV2V_UNCONNECTED_1843, SV2V_UNCONNECTED_1844, SV2V_UNCONNECTED_1845, SV2V_UNCONNECTED_1846, SV2V_UNCONNECTED_1847, SV2V_UNCONNECTED_1848, SV2V_UNCONNECTED_1849, SV2V_UNCONNECTED_1850, SV2V_UNCONNECTED_1851, SV2V_UNCONNECTED_1852, SV2V_UNCONNECTED_1853, SV2V_UNCONNECTED_1854, SV2V_UNCONNECTED_1855, SV2V_UNCONNECTED_1856, SV2V_UNCONNECTED_1857, SV2V_UNCONNECTED_1858, SV2V_UNCONNECTED_1859, SV2V_UNCONNECTED_1860, SV2V_UNCONNECTED_1861, SV2V_UNCONNECTED_1862, SV2V_UNCONNECTED_1863, SV2V_UNCONNECTED_1864, SV2V_UNCONNECTED_1865, SV2V_UNCONNECTED_1866, SV2V_UNCONNECTED_1867, SV2V_UNCONNECTED_1868, SV2V_UNCONNECTED_1869, SV2V_UNCONNECTED_1870, SV2V_UNCONNECTED_1871, SV2V_UNCONNECTED_1872, SV2V_UNCONNECTED_1873, SV2V_UNCONNECTED_1874, SV2V_UNCONNECTED_1875, SV2V_UNCONNECTED_1876, SV2V_UNCONNECTED_1877, SV2V_UNCONNECTED_1878, SV2V_UNCONNECTED_1879, SV2V_UNCONNECTED_1880, SV2V_UNCONNECTED_1881, SV2V_UNCONNECTED_1882, SV2V_UNCONNECTED_1883, SV2V_UNCONNECTED_1884, SV2V_UNCONNECTED_1885, SV2V_UNCONNECTED_1886, SV2V_UNCONNECTED_1887, SV2V_UNCONNECTED_1888, SV2V_UNCONNECTED_1889, SV2V_UNCONNECTED_1890, SV2V_UNCONNECTED_1891, SV2V_UNCONNECTED_1892, SV2V_UNCONNECTED_1893, SV2V_UNCONNECTED_1894, SV2V_UNCONNECTED_1895, SV2V_UNCONNECTED_1896, SV2V_UNCONNECTED_1897, SV2V_UNCONNECTED_1898, SV2V_UNCONNECTED_1899, SV2V_UNCONNECTED_1900, SV2V_UNCONNECTED_1901, SV2V_UNCONNECTED_1902, SV2V_UNCONNECTED_1903, SV2V_UNCONNECTED_1904, SV2V_UNCONNECTED_1905, SV2V_UNCONNECTED_1906, SV2V_UNCONNECTED_1907, SV2V_UNCONNECTED_1908, SV2V_UNCONNECTED_1909, SV2V_UNCONNECTED_1910, SV2V_UNCONNECTED_1911, SV2V_UNCONNECTED_1912, SV2V_UNCONNECTED_1913, SV2V_UNCONNECTED_1914, SV2V_UNCONNECTED_1915, SV2V_UNCONNECTED_1916, SV2V_UNCONNECTED_1917, SV2V_UNCONNECTED_1918, SV2V_UNCONNECTED_1919, SV2V_UNCONNECTED_1920, SV2V_UNCONNECTED_1921, SV2V_UNCONNECTED_1922, SV2V_UNCONNECTED_1923, SV2V_UNCONNECTED_1924, SV2V_UNCONNECTED_1925, SV2V_UNCONNECTED_1926, SV2V_UNCONNECTED_1927, SV2V_UNCONNECTED_1928, SV2V_UNCONNECTED_1929, SV2V_UNCONNECTED_1930, SV2V_UNCONNECTED_1931, SV2V_UNCONNECTED_1932, SV2V_UNCONNECTED_1933, SV2V_UNCONNECTED_1934, SV2V_UNCONNECTED_1935, SV2V_UNCONNECTED_1936, SV2V_UNCONNECTED_1937, SV2V_UNCONNECTED_1938, SV2V_UNCONNECTED_1939, SV2V_UNCONNECTED_1940, SV2V_UNCONNECTED_1941, SV2V_UNCONNECTED_1942, SV2V_UNCONNECTED_1943, SV2V_UNCONNECTED_1944, SV2V_UNCONNECTED_1945, SV2V_UNCONNECTED_1946, SV2V_UNCONNECTED_1947, SV2V_UNCONNECTED_1948, SV2V_UNCONNECTED_1949, SV2V_UNCONNECTED_1950, SV2V_UNCONNECTED_1951, SV2V_UNCONNECTED_1952, SV2V_UNCONNECTED_1953, SV2V_UNCONNECTED_1954, SV2V_UNCONNECTED_1955, SV2V_UNCONNECTED_1956, SV2V_UNCONNECTED_1957, SV2V_UNCONNECTED_1958, SV2V_UNCONNECTED_1959, SV2V_UNCONNECTED_1960, SV2V_UNCONNECTED_1961, SV2V_UNCONNECTED_1962, SV2V_UNCONNECTED_1963, SV2V_UNCONNECTED_1964, SV2V_UNCONNECTED_1965, SV2V_UNCONNECTED_1966, SV2V_UNCONNECTED_1967, SV2V_UNCONNECTED_1968, SV2V_UNCONNECTED_1969, SV2V_UNCONNECTED_1970, SV2V_UNCONNECTED_1971, SV2V_UNCONNECTED_1972, SV2V_UNCONNECTED_1973, SV2V_UNCONNECTED_1974, SV2V_UNCONNECTED_1975, SV2V_UNCONNECTED_1976, SV2V_UNCONNECTED_1977, SV2V_UNCONNECTED_1978, SV2V_UNCONNECTED_1979, SV2V_UNCONNECTED_1980, SV2V_UNCONNECTED_1981, SV2V_UNCONNECTED_1982, SV2V_UNCONNECTED_1983, SV2V_UNCONNECTED_1984, SV2V_UNCONNECTED_1985, SV2V_UNCONNECTED_1986, SV2V_UNCONNECTED_1987, SV2V_UNCONNECTED_1988, SV2V_UNCONNECTED_1989, SV2V_UNCONNECTED_1990, SV2V_UNCONNECTED_1991, SV2V_UNCONNECTED_1992, SV2V_UNCONNECTED_1993, SV2V_UNCONNECTED_1994, SV2V_UNCONNECTED_1995, SV2V_UNCONNECTED_1996, SV2V_UNCONNECTED_1997, SV2V_UNCONNECTED_1998, SV2V_UNCONNECTED_1999, SV2V_UNCONNECTED_2000, SV2V_UNCONNECTED_2001, SV2V_UNCONNECTED_2002, SV2V_UNCONNECTED_2003, SV2V_UNCONNECTED_2004, SV2V_UNCONNECTED_2005, SV2V_UNCONNECTED_2006, SV2V_UNCONNECTED_2007, SV2V_UNCONNECTED_2008, SV2V_UNCONNECTED_2009, SV2V_UNCONNECTED_2010, SV2V_UNCONNECTED_2011, SV2V_UNCONNECTED_2012, SV2V_UNCONNECTED_2013, SV2V_UNCONNECTED_2014, SV2V_UNCONNECTED_2015, SV2V_UNCONNECTED_2016, SV2V_UNCONNECTED_2017, SV2V_UNCONNECTED_2018, SV2V_UNCONNECTED_2019, SV2V_UNCONNECTED_2020, SV2V_UNCONNECTED_2021, SV2V_UNCONNECTED_2022, SV2V_UNCONNECTED_2023, SV2V_UNCONNECTED_2024, SV2V_UNCONNECTED_2025, SV2V_UNCONNECTED_2026, SV2V_UNCONNECTED_2027, SV2V_UNCONNECTED_2028, SV2V_UNCONNECTED_2029, SV2V_UNCONNECTED_2030, SV2V_UNCONNECTED_2031, SV2V_UNCONNECTED_2032, SV2V_UNCONNECTED_2033, SV2V_UNCONNECTED_2034, SV2V_UNCONNECTED_2035, SV2V_UNCONNECTED_2036, SV2V_UNCONNECTED_2037, SV2V_UNCONNECTED_2038, SV2V_UNCONNECTED_2039, SV2V_UNCONNECTED_2040, SV2V_UNCONNECTED_2041, SV2V_UNCONNECTED_2042, SV2V_UNCONNECTED_2043, SV2V_UNCONNECTED_2044, SV2V_UNCONNECTED_2045, SV2V_UNCONNECTED_2046, SV2V_UNCONNECTED_2047, SV2V_UNCONNECTED_2048, SV2V_UNCONNECTED_2049, SV2V_UNCONNECTED_2050, SV2V_UNCONNECTED_2051, SV2V_UNCONNECTED_2052, SV2V_UNCONNECTED_2053, SV2V_UNCONNECTED_2054, SV2V_UNCONNECTED_2055, SV2V_UNCONNECTED_2056, SV2V_UNCONNECTED_2057, SV2V_UNCONNECTED_2058, SV2V_UNCONNECTED_2059, SV2V_UNCONNECTED_2060, SV2V_UNCONNECTED_2061, SV2V_UNCONNECTED_2062, SV2V_UNCONNECTED_2063, SV2V_UNCONNECTED_2064, SV2V_UNCONNECTED_2065, SV2V_UNCONNECTED_2066, SV2V_UNCONNECTED_2067, SV2V_UNCONNECTED_2068, SV2V_UNCONNECTED_2069, SV2V_UNCONNECTED_2070, SV2V_UNCONNECTED_2071, SV2V_UNCONNECTED_2072, SV2V_UNCONNECTED_2073, SV2V_UNCONNECTED_2074, SV2V_UNCONNECTED_2075, SV2V_UNCONNECTED_2076, SV2V_UNCONNECTED_2077, SV2V_UNCONNECTED_2078, SV2V_UNCONNECTED_2079, SV2V_UNCONNECTED_2080, SV2V_UNCONNECTED_2081, SV2V_UNCONNECTED_2082, SV2V_UNCONNECTED_2083, SV2V_UNCONNECTED_2084, SV2V_UNCONNECTED_2085, SV2V_UNCONNECTED_2086, SV2V_UNCONNECTED_2087, SV2V_UNCONNECTED_2088, SV2V_UNCONNECTED_2089, SV2V_UNCONNECTED_2090, SV2V_UNCONNECTED_2091, SV2V_UNCONNECTED_2092, SV2V_UNCONNECTED_2093, SV2V_UNCONNECTED_2094, SV2V_UNCONNECTED_2095, SV2V_UNCONNECTED_2096, SV2V_UNCONNECTED_2097, SV2V_UNCONNECTED_2098, SV2V_UNCONNECTED_2099, SV2V_UNCONNECTED_2100, SV2V_UNCONNECTED_2101, SV2V_UNCONNECTED_2102, SV2V_UNCONNECTED_2103, SV2V_UNCONNECTED_2104, SV2V_UNCONNECTED_2105, SV2V_UNCONNECTED_2106, SV2V_UNCONNECTED_2107, SV2V_UNCONNECTED_2108, SV2V_UNCONNECTED_2109, SV2V_UNCONNECTED_2110, SV2V_UNCONNECTED_2111, SV2V_UNCONNECTED_2112, SV2V_UNCONNECTED_2113, SV2V_UNCONNECTED_2114, SV2V_UNCONNECTED_2115, SV2V_UNCONNECTED_2116, SV2V_UNCONNECTED_2117, SV2V_UNCONNECTED_2118, SV2V_UNCONNECTED_2119, SV2V_UNCONNECTED_2120, SV2V_UNCONNECTED_2121, SV2V_UNCONNECTED_2122, SV2V_UNCONNECTED_2123, SV2V_UNCONNECTED_2124, SV2V_UNCONNECTED_2125, SV2V_UNCONNECTED_2126, SV2V_UNCONNECTED_2127, SV2V_UNCONNECTED_2128, SV2V_UNCONNECTED_2129, SV2V_UNCONNECTED_2130, SV2V_UNCONNECTED_2131, SV2V_UNCONNECTED_2132, SV2V_UNCONNECTED_2133, SV2V_UNCONNECTED_2134, SV2V_UNCONNECTED_2135, SV2V_UNCONNECTED_2136, SV2V_UNCONNECTED_2137, SV2V_UNCONNECTED_2138, SV2V_UNCONNECTED_2139, SV2V_UNCONNECTED_2140, SV2V_UNCONNECTED_2141, SV2V_UNCONNECTED_2142, SV2V_UNCONNECTED_2143, SV2V_UNCONNECTED_2144, SV2V_UNCONNECTED_2145, SV2V_UNCONNECTED_2146, SV2V_UNCONNECTED_2147, SV2V_UNCONNECTED_2148, SV2V_UNCONNECTED_2149, SV2V_UNCONNECTED_2150, SV2V_UNCONNECTED_2151, SV2V_UNCONNECTED_2152, SV2V_UNCONNECTED_2153, SV2V_UNCONNECTED_2154, SV2V_UNCONNECTED_2155, SV2V_UNCONNECTED_2156, SV2V_UNCONNECTED_2157, SV2V_UNCONNECTED_2158, SV2V_UNCONNECTED_2159, SV2V_UNCONNECTED_2160, SV2V_UNCONNECTED_2161, SV2V_UNCONNECTED_2162, SV2V_UNCONNECTED_2163, SV2V_UNCONNECTED_2164, SV2V_UNCONNECTED_2165, SV2V_UNCONNECTED_2166, SV2V_UNCONNECTED_2167, SV2V_UNCONNECTED_2168, SV2V_UNCONNECTED_2169, SV2V_UNCONNECTED_2170, SV2V_UNCONNECTED_2171, SV2V_UNCONNECTED_2172, SV2V_UNCONNECTED_2173, SV2V_UNCONNECTED_2174, SV2V_UNCONNECTED_2175, SV2V_UNCONNECTED_2176, SV2V_UNCONNECTED_2177, SV2V_UNCONNECTED_2178, SV2V_UNCONNECTED_2179, SV2V_UNCONNECTED_2180, SV2V_UNCONNECTED_2181, SV2V_UNCONNECTED_2182, SV2V_UNCONNECTED_2183, SV2V_UNCONNECTED_2184, SV2V_UNCONNECTED_2185, SV2V_UNCONNECTED_2186, SV2V_UNCONNECTED_2187, SV2V_UNCONNECTED_2188, SV2V_UNCONNECTED_2189, SV2V_UNCONNECTED_2190, SV2V_UNCONNECTED_2191, SV2V_UNCONNECTED_2192, SV2V_UNCONNECTED_2193, SV2V_UNCONNECTED_2194, SV2V_UNCONNECTED_2195, SV2V_UNCONNECTED_2196, SV2V_UNCONNECTED_2197, SV2V_UNCONNECTED_2198, SV2V_UNCONNECTED_2199, SV2V_UNCONNECTED_2200, SV2V_UNCONNECTED_2201, SV2V_UNCONNECTED_2202, SV2V_UNCONNECTED_2203, SV2V_UNCONNECTED_2204, SV2V_UNCONNECTED_2205, SV2V_UNCONNECTED_2206, SV2V_UNCONNECTED_2207, SV2V_UNCONNECTED_2208, SV2V_UNCONNECTED_2209, SV2V_UNCONNECTED_2210, SV2V_UNCONNECTED_2211, SV2V_UNCONNECTED_2212, SV2V_UNCONNECTED_2213, SV2V_UNCONNECTED_2214, SV2V_UNCONNECTED_2215, SV2V_UNCONNECTED_2216, SV2V_UNCONNECTED_2217, SV2V_UNCONNECTED_2218, SV2V_UNCONNECTED_2219, SV2V_UNCONNECTED_2220, SV2V_UNCONNECTED_2221, SV2V_UNCONNECTED_2222, SV2V_UNCONNECTED_2223, SV2V_UNCONNECTED_2224, SV2V_UNCONNECTED_2225, SV2V_UNCONNECTED_2226, SV2V_UNCONNECTED_2227, SV2V_UNCONNECTED_2228, SV2V_UNCONNECTED_2229, SV2V_UNCONNECTED_2230, SV2V_UNCONNECTED_2231, SV2V_UNCONNECTED_2232, SV2V_UNCONNECTED_2233, SV2V_UNCONNECTED_2234, SV2V_UNCONNECTED_2235, SV2V_UNCONNECTED_2236, SV2V_UNCONNECTED_2237, SV2V_UNCONNECTED_2238, SV2V_UNCONNECTED_2239, SV2V_UNCONNECTED_2240, SV2V_UNCONNECTED_2241, SV2V_UNCONNECTED_2242, SV2V_UNCONNECTED_2243, SV2V_UNCONNECTED_2244, SV2V_UNCONNECTED_2245, SV2V_UNCONNECTED_2246, SV2V_UNCONNECTED_2247, SV2V_UNCONNECTED_2248, SV2V_UNCONNECTED_2249, SV2V_UNCONNECTED_2250, SV2V_UNCONNECTED_2251, SV2V_UNCONNECTED_2252, SV2V_UNCONNECTED_2253, SV2V_UNCONNECTED_2254, SV2V_UNCONNECTED_2255, SV2V_UNCONNECTED_2256, SV2V_UNCONNECTED_2257, SV2V_UNCONNECTED_2258, SV2V_UNCONNECTED_2259, SV2V_UNCONNECTED_2260, SV2V_UNCONNECTED_2261, SV2V_UNCONNECTED_2262, SV2V_UNCONNECTED_2263, SV2V_UNCONNECTED_2264, SV2V_UNCONNECTED_2265, SV2V_UNCONNECTED_2266, SV2V_UNCONNECTED_2267, SV2V_UNCONNECTED_2268, SV2V_UNCONNECTED_2269, SV2V_UNCONNECTED_2270, SV2V_UNCONNECTED_2271, SV2V_UNCONNECTED_2272, SV2V_UNCONNECTED_2273, SV2V_UNCONNECTED_2274, SV2V_UNCONNECTED_2275, SV2V_UNCONNECTED_2276, SV2V_UNCONNECTED_2277, SV2V_UNCONNECTED_2278, SV2V_UNCONNECTED_2279, SV2V_UNCONNECTED_2280, SV2V_UNCONNECTED_2281, SV2V_UNCONNECTED_2282, SV2V_UNCONNECTED_2283, SV2V_UNCONNECTED_2284, SV2V_UNCONNECTED_2285, SV2V_UNCONNECTED_2286, SV2V_UNCONNECTED_2287, SV2V_UNCONNECTED_2288, SV2V_UNCONNECTED_2289, SV2V_UNCONNECTED_2290, SV2V_UNCONNECTED_2291, SV2V_UNCONNECTED_2292, SV2V_UNCONNECTED_2293, SV2V_UNCONNECTED_2294, SV2V_UNCONNECTED_2295, SV2V_UNCONNECTED_2296, SV2V_UNCONNECTED_2297, SV2V_UNCONNECTED_2298, SV2V_UNCONNECTED_2299, SV2V_UNCONNECTED_2300, SV2V_UNCONNECTED_2301, SV2V_UNCONNECTED_2302, SV2V_UNCONNECTED_2303, SV2V_UNCONNECTED_2304, SV2V_UNCONNECTED_2305, SV2V_UNCONNECTED_2306, SV2V_UNCONNECTED_2307, SV2V_UNCONNECTED_2308, SV2V_UNCONNECTED_2309, SV2V_UNCONNECTED_2310, SV2V_UNCONNECTED_2311, SV2V_UNCONNECTED_2312, SV2V_UNCONNECTED_2313, SV2V_UNCONNECTED_2314, SV2V_UNCONNECTED_2315, SV2V_UNCONNECTED_2316, SV2V_UNCONNECTED_2317, SV2V_UNCONNECTED_2318, SV2V_UNCONNECTED_2319, SV2V_UNCONNECTED_2320, SV2V_UNCONNECTED_2321, SV2V_UNCONNECTED_2322, SV2V_UNCONNECTED_2323, SV2V_UNCONNECTED_2324, SV2V_UNCONNECTED_2325, SV2V_UNCONNECTED_2326, SV2V_UNCONNECTED_2327, SV2V_UNCONNECTED_2328, SV2V_UNCONNECTED_2329, SV2V_UNCONNECTED_2330, SV2V_UNCONNECTED_2331, SV2V_UNCONNECTED_2332, SV2V_UNCONNECTED_2333, SV2V_UNCONNECTED_2334, SV2V_UNCONNECTED_2335, SV2V_UNCONNECTED_2336, SV2V_UNCONNECTED_2337, SV2V_UNCONNECTED_2338, SV2V_UNCONNECTED_2339, SV2V_UNCONNECTED_2340, SV2V_UNCONNECTED_2341, SV2V_UNCONNECTED_2342, SV2V_UNCONNECTED_2343, SV2V_UNCONNECTED_2344, SV2V_UNCONNECTED_2345, SV2V_UNCONNECTED_2346, SV2V_UNCONNECTED_2347, SV2V_UNCONNECTED_2348, SV2V_UNCONNECTED_2349, SV2V_UNCONNECTED_2350, SV2V_UNCONNECTED_2351, SV2V_UNCONNECTED_2352, SV2V_UNCONNECTED_2353, SV2V_UNCONNECTED_2354, SV2V_UNCONNECTED_2355, SV2V_UNCONNECTED_2356, SV2V_UNCONNECTED_2357, SV2V_UNCONNECTED_2358, SV2V_UNCONNECTED_2359, SV2V_UNCONNECTED_2360, SV2V_UNCONNECTED_2361, SV2V_UNCONNECTED_2362, SV2V_UNCONNECTED_2363, SV2V_UNCONNECTED_2364, SV2V_UNCONNECTED_2365, SV2V_UNCONNECTED_2366, SV2V_UNCONNECTED_2367, SV2V_UNCONNECTED_2368, SV2V_UNCONNECTED_2369, SV2V_UNCONNECTED_2370, SV2V_UNCONNECTED_2371, SV2V_UNCONNECTED_2372, SV2V_UNCONNECTED_2373, SV2V_UNCONNECTED_2374, SV2V_UNCONNECTED_2375, SV2V_UNCONNECTED_2376, SV2V_UNCONNECTED_2377, SV2V_UNCONNECTED_2378, SV2V_UNCONNECTED_2379, SV2V_UNCONNECTED_2380, SV2V_UNCONNECTED_2381, SV2V_UNCONNECTED_2382, SV2V_UNCONNECTED_2383, SV2V_UNCONNECTED_2384, SV2V_UNCONNECTED_2385, SV2V_UNCONNECTED_2386, SV2V_UNCONNECTED_2387, SV2V_UNCONNECTED_2388, SV2V_UNCONNECTED_2389, SV2V_UNCONNECTED_2390, SV2V_UNCONNECTED_2391, SV2V_UNCONNECTED_2392, SV2V_UNCONNECTED_2393, SV2V_UNCONNECTED_2394, SV2V_UNCONNECTED_2395, SV2V_UNCONNECTED_2396, SV2V_UNCONNECTED_2397, SV2V_UNCONNECTED_2398, SV2V_UNCONNECTED_2399, SV2V_UNCONNECTED_2400, SV2V_UNCONNECTED_2401, SV2V_UNCONNECTED_2402, SV2V_UNCONNECTED_2403, SV2V_UNCONNECTED_2404, SV2V_UNCONNECTED_2405, SV2V_UNCONNECTED_2406, SV2V_UNCONNECTED_2407, SV2V_UNCONNECTED_2408, SV2V_UNCONNECTED_2409, SV2V_UNCONNECTED_2410, SV2V_UNCONNECTED_2411, SV2V_UNCONNECTED_2412, SV2V_UNCONNECTED_2413, SV2V_UNCONNECTED_2414, SV2V_UNCONNECTED_2415, SV2V_UNCONNECTED_2416, SV2V_UNCONNECTED_2417, SV2V_UNCONNECTED_2418, SV2V_UNCONNECTED_2419, SV2V_UNCONNECTED_2420, SV2V_UNCONNECTED_2421, SV2V_UNCONNECTED_2422, SV2V_UNCONNECTED_2423, SV2V_UNCONNECTED_2424, SV2V_UNCONNECTED_2425, SV2V_UNCONNECTED_2426, SV2V_UNCONNECTED_2427, SV2V_UNCONNECTED_2428, SV2V_UNCONNECTED_2429, SV2V_UNCONNECTED_2430, SV2V_UNCONNECTED_2431, SV2V_UNCONNECTED_2432, SV2V_UNCONNECTED_2433, SV2V_UNCONNECTED_2434, SV2V_UNCONNECTED_2435, SV2V_UNCONNECTED_2436, SV2V_UNCONNECTED_2437, SV2V_UNCONNECTED_2438, SV2V_UNCONNECTED_2439, SV2V_UNCONNECTED_2440, SV2V_UNCONNECTED_2441, SV2V_UNCONNECTED_2442, SV2V_UNCONNECTED_2443, SV2V_UNCONNECTED_2444, SV2V_UNCONNECTED_2445, SV2V_UNCONNECTED_2446, SV2V_UNCONNECTED_2447, SV2V_UNCONNECTED_2448, SV2V_UNCONNECTED_2449, SV2V_UNCONNECTED_2450, SV2V_UNCONNECTED_2451, SV2V_UNCONNECTED_2452, SV2V_UNCONNECTED_2453, SV2V_UNCONNECTED_2454, SV2V_UNCONNECTED_2455, SV2V_UNCONNECTED_2456, SV2V_UNCONNECTED_2457, SV2V_UNCONNECTED_2458, SV2V_UNCONNECTED_2459, SV2V_UNCONNECTED_2460, SV2V_UNCONNECTED_2461, SV2V_UNCONNECTED_2462, SV2V_UNCONNECTED_2463, SV2V_UNCONNECTED_2464, SV2V_UNCONNECTED_2465, SV2V_UNCONNECTED_2466, SV2V_UNCONNECTED_2467, SV2V_UNCONNECTED_2468, SV2V_UNCONNECTED_2469, SV2V_UNCONNECTED_2470, SV2V_UNCONNECTED_2471, SV2V_UNCONNECTED_2472, SV2V_UNCONNECTED_2473, SV2V_UNCONNECTED_2474, SV2V_UNCONNECTED_2475, SV2V_UNCONNECTED_2476, SV2V_UNCONNECTED_2477, SV2V_UNCONNECTED_2478, SV2V_UNCONNECTED_2479, SV2V_UNCONNECTED_2480, SV2V_UNCONNECTED_2481, SV2V_UNCONNECTED_2482, SV2V_UNCONNECTED_2483, SV2V_UNCONNECTED_2484, SV2V_UNCONNECTED_2485, SV2V_UNCONNECTED_2486, SV2V_UNCONNECTED_2487, SV2V_UNCONNECTED_2488, SV2V_UNCONNECTED_2489, SV2V_UNCONNECTED_2490, SV2V_UNCONNECTED_2491, SV2V_UNCONNECTED_2492, SV2V_UNCONNECTED_2493, SV2V_UNCONNECTED_2494, SV2V_UNCONNECTED_2495, SV2V_UNCONNECTED_2496, SV2V_UNCONNECTED_2497, SV2V_UNCONNECTED_2498, SV2V_UNCONNECTED_2499, SV2V_UNCONNECTED_2500, SV2V_UNCONNECTED_2501, SV2V_UNCONNECTED_2502, SV2V_UNCONNECTED_2503, SV2V_UNCONNECTED_2504, SV2V_UNCONNECTED_2505, SV2V_UNCONNECTED_2506, SV2V_UNCONNECTED_2507, SV2V_UNCONNECTED_2508, SV2V_UNCONNECTED_2509, SV2V_UNCONNECTED_2510, SV2V_UNCONNECTED_2511, SV2V_UNCONNECTED_2512, SV2V_UNCONNECTED_2513, SV2V_UNCONNECTED_2514, SV2V_UNCONNECTED_2515, SV2V_UNCONNECTED_2516, SV2V_UNCONNECTED_2517, SV2V_UNCONNECTED_2518, SV2V_UNCONNECTED_2519, SV2V_UNCONNECTED_2520, SV2V_UNCONNECTED_2521, SV2V_UNCONNECTED_2522, SV2V_UNCONNECTED_2523, SV2V_UNCONNECTED_2524, SV2V_UNCONNECTED_2525, SV2V_UNCONNECTED_2526, SV2V_UNCONNECTED_2527, SV2V_UNCONNECTED_2528, SV2V_UNCONNECTED_2529, SV2V_UNCONNECTED_2530, SV2V_UNCONNECTED_2531, SV2V_UNCONNECTED_2532, SV2V_UNCONNECTED_2533, SV2V_UNCONNECTED_2534, SV2V_UNCONNECTED_2535, SV2V_UNCONNECTED_2536, SV2V_UNCONNECTED_2537, SV2V_UNCONNECTED_2538, SV2V_UNCONNECTED_2539, SV2V_UNCONNECTED_2540, SV2V_UNCONNECTED_2541, SV2V_UNCONNECTED_2542, SV2V_UNCONNECTED_2543, SV2V_UNCONNECTED_2544, SV2V_UNCONNECTED_2545, SV2V_UNCONNECTED_2546, SV2V_UNCONNECTED_2547, SV2V_UNCONNECTED_2548, SV2V_UNCONNECTED_2549, SV2V_UNCONNECTED_2550, SV2V_UNCONNECTED_2551, SV2V_UNCONNECTED_2552, SV2V_UNCONNECTED_2553, SV2V_UNCONNECTED_2554, SV2V_UNCONNECTED_2555, SV2V_UNCONNECTED_2556, SV2V_UNCONNECTED_2557, SV2V_UNCONNECTED_2558, SV2V_UNCONNECTED_2559, SV2V_UNCONNECTED_2560, SV2V_UNCONNECTED_2561, SV2V_UNCONNECTED_2562, SV2V_UNCONNECTED_2563, SV2V_UNCONNECTED_2564, SV2V_UNCONNECTED_2565, SV2V_UNCONNECTED_2566, SV2V_UNCONNECTED_2567, SV2V_UNCONNECTED_2568, SV2V_UNCONNECTED_2569, SV2V_UNCONNECTED_2570, SV2V_UNCONNECTED_2571, SV2V_UNCONNECTED_2572, SV2V_UNCONNECTED_2573, SV2V_UNCONNECTED_2574, SV2V_UNCONNECTED_2575, SV2V_UNCONNECTED_2576, SV2V_UNCONNECTED_2577, SV2V_UNCONNECTED_2578, SV2V_UNCONNECTED_2579, SV2V_UNCONNECTED_2580, SV2V_UNCONNECTED_2581, SV2V_UNCONNECTED_2582, SV2V_UNCONNECTED_2583, SV2V_UNCONNECTED_2584, SV2V_UNCONNECTED_2585, SV2V_UNCONNECTED_2586, SV2V_UNCONNECTED_2587, SV2V_UNCONNECTED_2588, SV2V_UNCONNECTED_2589, SV2V_UNCONNECTED_2590, SV2V_UNCONNECTED_2591, SV2V_UNCONNECTED_2592, SV2V_UNCONNECTED_2593, SV2V_UNCONNECTED_2594, SV2V_UNCONNECTED_2595, SV2V_UNCONNECTED_2596, SV2V_UNCONNECTED_2597, SV2V_UNCONNECTED_2598, SV2V_UNCONNECTED_2599, SV2V_UNCONNECTED_2600, SV2V_UNCONNECTED_2601, SV2V_UNCONNECTED_2602, SV2V_UNCONNECTED_2603, SV2V_UNCONNECTED_2604, SV2V_UNCONNECTED_2605, SV2V_UNCONNECTED_2606, SV2V_UNCONNECTED_2607, SV2V_UNCONNECTED_2608, SV2V_UNCONNECTED_2609, SV2V_UNCONNECTED_2610, SV2V_UNCONNECTED_2611, SV2V_UNCONNECTED_2612, SV2V_UNCONNECTED_2613, SV2V_UNCONNECTED_2614, SV2V_UNCONNECTED_2615, SV2V_UNCONNECTED_2616, SV2V_UNCONNECTED_2617, SV2V_UNCONNECTED_2618, SV2V_UNCONNECTED_2619, SV2V_UNCONNECTED_2620, SV2V_UNCONNECTED_2621, SV2V_UNCONNECTED_2622, SV2V_UNCONNECTED_2623, SV2V_UNCONNECTED_2624, SV2V_UNCONNECTED_2625, SV2V_UNCONNECTED_2626, SV2V_UNCONNECTED_2627, SV2V_UNCONNECTED_2628, SV2V_UNCONNECTED_2629, SV2V_UNCONNECTED_2630, SV2V_UNCONNECTED_2631, SV2V_UNCONNECTED_2632, SV2V_UNCONNECTED_2633, SV2V_UNCONNECTED_2634, SV2V_UNCONNECTED_2635, SV2V_UNCONNECTED_2636, SV2V_UNCONNECTED_2637, SV2V_UNCONNECTED_2638, SV2V_UNCONNECTED_2639, SV2V_UNCONNECTED_2640, SV2V_UNCONNECTED_2641, SV2V_UNCONNECTED_2642, SV2V_UNCONNECTED_2643, SV2V_UNCONNECTED_2644, SV2V_UNCONNECTED_2645, SV2V_UNCONNECTED_2646, SV2V_UNCONNECTED_2647, SV2V_UNCONNECTED_2648, SV2V_UNCONNECTED_2649, SV2V_UNCONNECTED_2650, SV2V_UNCONNECTED_2651, SV2V_UNCONNECTED_2652, SV2V_UNCONNECTED_2653, SV2V_UNCONNECTED_2654, SV2V_UNCONNECTED_2655, SV2V_UNCONNECTED_2656, SV2V_UNCONNECTED_2657, SV2V_UNCONNECTED_2658, SV2V_UNCONNECTED_2659, SV2V_UNCONNECTED_2660, SV2V_UNCONNECTED_2661, SV2V_UNCONNECTED_2662, SV2V_UNCONNECTED_2663, SV2V_UNCONNECTED_2664, SV2V_UNCONNECTED_2665, SV2V_UNCONNECTED_2666, SV2V_UNCONNECTED_2667, SV2V_UNCONNECTED_2668, SV2V_UNCONNECTED_2669, SV2V_UNCONNECTED_2670, SV2V_UNCONNECTED_2671, SV2V_UNCONNECTED_2672, SV2V_UNCONNECTED_2673, SV2V_UNCONNECTED_2674, SV2V_UNCONNECTED_2675, SV2V_UNCONNECTED_2676, SV2V_UNCONNECTED_2677, SV2V_UNCONNECTED_2678, SV2V_UNCONNECTED_2679, SV2V_UNCONNECTED_2680, SV2V_UNCONNECTED_2681, SV2V_UNCONNECTED_2682, SV2V_UNCONNECTED_2683, SV2V_UNCONNECTED_2684, SV2V_UNCONNECTED_2685, SV2V_UNCONNECTED_2686, SV2V_UNCONNECTED_2687, SV2V_UNCONNECTED_2688, SV2V_UNCONNECTED_2689, SV2V_UNCONNECTED_2690, SV2V_UNCONNECTED_2691, SV2V_UNCONNECTED_2692, SV2V_UNCONNECTED_2693, SV2V_UNCONNECTED_2694, SV2V_UNCONNECTED_2695, SV2V_UNCONNECTED_2696, SV2V_UNCONNECTED_2697, SV2V_UNCONNECTED_2698, SV2V_UNCONNECTED_2699, SV2V_UNCONNECTED_2700, SV2V_UNCONNECTED_2701, SV2V_UNCONNECTED_2702, SV2V_UNCONNECTED_2703, SV2V_UNCONNECTED_2704, SV2V_UNCONNECTED_2705, SV2V_UNCONNECTED_2706, SV2V_UNCONNECTED_2707, SV2V_UNCONNECTED_2708, SV2V_UNCONNECTED_2709, SV2V_UNCONNECTED_2710, SV2V_UNCONNECTED_2711, SV2V_UNCONNECTED_2712, SV2V_UNCONNECTED_2713, SV2V_UNCONNECTED_2714, SV2V_UNCONNECTED_2715, SV2V_UNCONNECTED_2716, SV2V_UNCONNECTED_2717, SV2V_UNCONNECTED_2718, SV2V_UNCONNECTED_2719, SV2V_UNCONNECTED_2720, SV2V_UNCONNECTED_2721, SV2V_UNCONNECTED_2722, SV2V_UNCONNECTED_2723, SV2V_UNCONNECTED_2724, SV2V_UNCONNECTED_2725, SV2V_UNCONNECTED_2726, SV2V_UNCONNECTED_2727, SV2V_UNCONNECTED_2728, SV2V_UNCONNECTED_2729, SV2V_UNCONNECTED_2730, SV2V_UNCONNECTED_2731, SV2V_UNCONNECTED_2732, SV2V_UNCONNECTED_2733, SV2V_UNCONNECTED_2734, SV2V_UNCONNECTED_2735, SV2V_UNCONNECTED_2736, SV2V_UNCONNECTED_2737, SV2V_UNCONNECTED_2738, SV2V_UNCONNECTED_2739, SV2V_UNCONNECTED_2740, SV2V_UNCONNECTED_2741, SV2V_UNCONNECTED_2742, SV2V_UNCONNECTED_2743, SV2V_UNCONNECTED_2744, SV2V_UNCONNECTED_2745, SV2V_UNCONNECTED_2746, SV2V_UNCONNECTED_2747, SV2V_UNCONNECTED_2748, SV2V_UNCONNECTED_2749, SV2V_UNCONNECTED_2750, SV2V_UNCONNECTED_2751, SV2V_UNCONNECTED_2752, SV2V_UNCONNECTED_2753, SV2V_UNCONNECTED_2754, SV2V_UNCONNECTED_2755, SV2V_UNCONNECTED_2756, SV2V_UNCONNECTED_2757, SV2V_UNCONNECTED_2758, SV2V_UNCONNECTED_2759, SV2V_UNCONNECTED_2760, SV2V_UNCONNECTED_2761, SV2V_UNCONNECTED_2762, SV2V_UNCONNECTED_2763, SV2V_UNCONNECTED_2764, SV2V_UNCONNECTED_2765, SV2V_UNCONNECTED_2766, SV2V_UNCONNECTED_2767, SV2V_UNCONNECTED_2768, SV2V_UNCONNECTED_2769, SV2V_UNCONNECTED_2770, SV2V_UNCONNECTED_2771, SV2V_UNCONNECTED_2772, SV2V_UNCONNECTED_2773, SV2V_UNCONNECTED_2774, SV2V_UNCONNECTED_2775, SV2V_UNCONNECTED_2776, SV2V_UNCONNECTED_2777, SV2V_UNCONNECTED_2778, SV2V_UNCONNECTED_2779, SV2V_UNCONNECTED_2780, SV2V_UNCONNECTED_2781, SV2V_UNCONNECTED_2782, SV2V_UNCONNECTED_2783, SV2V_UNCONNECTED_2784, SV2V_UNCONNECTED_2785, SV2V_UNCONNECTED_2786, SV2V_UNCONNECTED_2787, SV2V_UNCONNECTED_2788, SV2V_UNCONNECTED_2789, SV2V_UNCONNECTED_2790, SV2V_UNCONNECTED_2791, SV2V_UNCONNECTED_2792, SV2V_UNCONNECTED_2793, SV2V_UNCONNECTED_2794, SV2V_UNCONNECTED_2795, SV2V_UNCONNECTED_2796, SV2V_UNCONNECTED_2797, SV2V_UNCONNECTED_2798, SV2V_UNCONNECTED_2799, SV2V_UNCONNECTED_2800, SV2V_UNCONNECTED_2801, SV2V_UNCONNECTED_2802, SV2V_UNCONNECTED_2803, SV2V_UNCONNECTED_2804, SV2V_UNCONNECTED_2805, SV2V_UNCONNECTED_2806, SV2V_UNCONNECTED_2807, SV2V_UNCONNECTED_2808, SV2V_UNCONNECTED_2809, SV2V_UNCONNECTED_2810, SV2V_UNCONNECTED_2811, SV2V_UNCONNECTED_2812, SV2V_UNCONNECTED_2813, SV2V_UNCONNECTED_2814, SV2V_UNCONNECTED_2815, SV2V_UNCONNECTED_2816, SV2V_UNCONNECTED_2817, SV2V_UNCONNECTED_2818, SV2V_UNCONNECTED_2819, SV2V_UNCONNECTED_2820, SV2V_UNCONNECTED_2821, SV2V_UNCONNECTED_2822, SV2V_UNCONNECTED_2823, SV2V_UNCONNECTED_2824, SV2V_UNCONNECTED_2825, SV2V_UNCONNECTED_2826, SV2V_UNCONNECTED_2827, SV2V_UNCONNECTED_2828, SV2V_UNCONNECTED_2829, SV2V_UNCONNECTED_2830, SV2V_UNCONNECTED_2831, SV2V_UNCONNECTED_2832, SV2V_UNCONNECTED_2833, SV2V_UNCONNECTED_2834, SV2V_UNCONNECTED_2835, SV2V_UNCONNECTED_2836, SV2V_UNCONNECTED_2837, SV2V_UNCONNECTED_2838, SV2V_UNCONNECTED_2839, SV2V_UNCONNECTED_2840, SV2V_UNCONNECTED_2841, SV2V_UNCONNECTED_2842, SV2V_UNCONNECTED_2843, SV2V_UNCONNECTED_2844, SV2V_UNCONNECTED_2845, SV2V_UNCONNECTED_2846, SV2V_UNCONNECTED_2847, SV2V_UNCONNECTED_2848, SV2V_UNCONNECTED_2849, SV2V_UNCONNECTED_2850, SV2V_UNCONNECTED_2851, SV2V_UNCONNECTED_2852, SV2V_UNCONNECTED_2853, SV2V_UNCONNECTED_2854, SV2V_UNCONNECTED_2855, SV2V_UNCONNECTED_2856, SV2V_UNCONNECTED_2857, SV2V_UNCONNECTED_2858, SV2V_UNCONNECTED_2859, SV2V_UNCONNECTED_2860, SV2V_UNCONNECTED_2861, SV2V_UNCONNECTED_2862, SV2V_UNCONNECTED_2863, SV2V_UNCONNECTED_2864, SV2V_UNCONNECTED_2865, SV2V_UNCONNECTED_2866, SV2V_UNCONNECTED_2867, SV2V_UNCONNECTED_2868, SV2V_UNCONNECTED_2869, SV2V_UNCONNECTED_2870, SV2V_UNCONNECTED_2871, SV2V_UNCONNECTED_2872, SV2V_UNCONNECTED_2873, SV2V_UNCONNECTED_2874, SV2V_UNCONNECTED_2875, SV2V_UNCONNECTED_2876, SV2V_UNCONNECTED_2877, SV2V_UNCONNECTED_2878, SV2V_UNCONNECTED_2879, SV2V_UNCONNECTED_2880, SV2V_UNCONNECTED_2881, SV2V_UNCONNECTED_2882, SV2V_UNCONNECTED_2883, SV2V_UNCONNECTED_2884, SV2V_UNCONNECTED_2885, SV2V_UNCONNECTED_2886, SV2V_UNCONNECTED_2887, SV2V_UNCONNECTED_2888, SV2V_UNCONNECTED_2889, SV2V_UNCONNECTED_2890, SV2V_UNCONNECTED_2891, SV2V_UNCONNECTED_2892, SV2V_UNCONNECTED_2893, SV2V_UNCONNECTED_2894, SV2V_UNCONNECTED_2895, SV2V_UNCONNECTED_2896, SV2V_UNCONNECTED_2897, SV2V_UNCONNECTED_2898, SV2V_UNCONNECTED_2899, SV2V_UNCONNECTED_2900, SV2V_UNCONNECTED_2901, SV2V_UNCONNECTED_2902, SV2V_UNCONNECTED_2903, SV2V_UNCONNECTED_2904, SV2V_UNCONNECTED_2905, SV2V_UNCONNECTED_2906, SV2V_UNCONNECTED_2907, SV2V_UNCONNECTED_2908, SV2V_UNCONNECTED_2909, SV2V_UNCONNECTED_2910, SV2V_UNCONNECTED_2911, SV2V_UNCONNECTED_2912, SV2V_UNCONNECTED_2913, SV2V_UNCONNECTED_2914, SV2V_UNCONNECTED_2915, SV2V_UNCONNECTED_2916, SV2V_UNCONNECTED_2917, SV2V_UNCONNECTED_2918, SV2V_UNCONNECTED_2919, SV2V_UNCONNECTED_2920, SV2V_UNCONNECTED_2921, SV2V_UNCONNECTED_2922, SV2V_UNCONNECTED_2923, SV2V_UNCONNECTED_2924, SV2V_UNCONNECTED_2925, SV2V_UNCONNECTED_2926, SV2V_UNCONNECTED_2927, SV2V_UNCONNECTED_2928, SV2V_UNCONNECTED_2929, SV2V_UNCONNECTED_2930, SV2V_UNCONNECTED_2931, SV2V_UNCONNECTED_2932, SV2V_UNCONNECTED_2933, SV2V_UNCONNECTED_2934, SV2V_UNCONNECTED_2935, SV2V_UNCONNECTED_2936, SV2V_UNCONNECTED_2937, SV2V_UNCONNECTED_2938, SV2V_UNCONNECTED_2939, SV2V_UNCONNECTED_2940, SV2V_UNCONNECTED_2941, SV2V_UNCONNECTED_2942, SV2V_UNCONNECTED_2943, SV2V_UNCONNECTED_2944, SV2V_UNCONNECTED_2945, SV2V_UNCONNECTED_2946, SV2V_UNCONNECTED_2947, SV2V_UNCONNECTED_2948, SV2V_UNCONNECTED_2949, SV2V_UNCONNECTED_2950, SV2V_UNCONNECTED_2951, SV2V_UNCONNECTED_2952, SV2V_UNCONNECTED_2953, SV2V_UNCONNECTED_2954, SV2V_UNCONNECTED_2955, SV2V_UNCONNECTED_2956, SV2V_UNCONNECTED_2957, SV2V_UNCONNECTED_2958, SV2V_UNCONNECTED_2959, SV2V_UNCONNECTED_2960, SV2V_UNCONNECTED_2961, SV2V_UNCONNECTED_2962, SV2V_UNCONNECTED_2963, SV2V_UNCONNECTED_2964, SV2V_UNCONNECTED_2965, SV2V_UNCONNECTED_2966, SV2V_UNCONNECTED_2967, SV2V_UNCONNECTED_2968, SV2V_UNCONNECTED_2969, SV2V_UNCONNECTED_2970, SV2V_UNCONNECTED_2971, SV2V_UNCONNECTED_2972, SV2V_UNCONNECTED_2973, SV2V_UNCONNECTED_2974, SV2V_UNCONNECTED_2975, SV2V_UNCONNECTED_2976, SV2V_UNCONNECTED_2977, SV2V_UNCONNECTED_2978, SV2V_UNCONNECTED_2979, SV2V_UNCONNECTED_2980, SV2V_UNCONNECTED_2981, SV2V_UNCONNECTED_2982, SV2V_UNCONNECTED_2983, SV2V_UNCONNECTED_2984, SV2V_UNCONNECTED_2985, SV2V_UNCONNECTED_2986, SV2V_UNCONNECTED_2987, SV2V_UNCONNECTED_2988, SV2V_UNCONNECTED_2989, SV2V_UNCONNECTED_2990, SV2V_UNCONNECTED_2991, SV2V_UNCONNECTED_2992, SV2V_UNCONNECTED_2993, SV2V_UNCONNECTED_2994, SV2V_UNCONNECTED_2995, SV2V_UNCONNECTED_2996, SV2V_UNCONNECTED_2997, SV2V_UNCONNECTED_2998, SV2V_UNCONNECTED_2999, SV2V_UNCONNECTED_3000, SV2V_UNCONNECTED_3001, SV2V_UNCONNECTED_3002, SV2V_UNCONNECTED_3003, SV2V_UNCONNECTED_3004, SV2V_UNCONNECTED_3005, SV2V_UNCONNECTED_3006, SV2V_UNCONNECTED_3007, SV2V_UNCONNECTED_3008, SV2V_UNCONNECTED_3009, SV2V_UNCONNECTED_3010, SV2V_UNCONNECTED_3011, SV2V_UNCONNECTED_3012, SV2V_UNCONNECTED_3013, SV2V_UNCONNECTED_3014, SV2V_UNCONNECTED_3015, SV2V_UNCONNECTED_3016, SV2V_UNCONNECTED_3017, SV2V_UNCONNECTED_3018, SV2V_UNCONNECTED_3019, SV2V_UNCONNECTED_3020, SV2V_UNCONNECTED_3021, SV2V_UNCONNECTED_3022, SV2V_UNCONNECTED_3023, SV2V_UNCONNECTED_3024, SV2V_UNCONNECTED_3025, SV2V_UNCONNECTED_3026, SV2V_UNCONNECTED_3027, SV2V_UNCONNECTED_3028, SV2V_UNCONNECTED_3029, SV2V_UNCONNECTED_3030, SV2V_UNCONNECTED_3031, SV2V_UNCONNECTED_3032, SV2V_UNCONNECTED_3033, SV2V_UNCONNECTED_3034, SV2V_UNCONNECTED_3035, SV2V_UNCONNECTED_3036, SV2V_UNCONNECTED_3037, SV2V_UNCONNECTED_3038, SV2V_UNCONNECTED_3039, SV2V_UNCONNECTED_3040, SV2V_UNCONNECTED_3041, SV2V_UNCONNECTED_3042, SV2V_UNCONNECTED_3043, SV2V_UNCONNECTED_3044, SV2V_UNCONNECTED_3045, SV2V_UNCONNECTED_3046, SV2V_UNCONNECTED_3047, SV2V_UNCONNECTED_3048, SV2V_UNCONNECTED_3049, SV2V_UNCONNECTED_3050, SV2V_UNCONNECTED_3051, SV2V_UNCONNECTED_3052, SV2V_UNCONNECTED_3053, SV2V_UNCONNECTED_3054, SV2V_UNCONNECTED_3055, SV2V_UNCONNECTED_3056, SV2V_UNCONNECTED_3057, SV2V_UNCONNECTED_3058, SV2V_UNCONNECTED_3059, SV2V_UNCONNECTED_3060, SV2V_UNCONNECTED_3061, SV2V_UNCONNECTED_3062, SV2V_UNCONNECTED_3063, SV2V_UNCONNECTED_3064, SV2V_UNCONNECTED_3065, SV2V_UNCONNECTED_3066, SV2V_UNCONNECTED_3067, SV2V_UNCONNECTED_3068, SV2V_UNCONNECTED_3069, SV2V_UNCONNECTED_3070, SV2V_UNCONNECTED_3071, SV2V_UNCONNECTED_3072, SV2V_UNCONNECTED_3073, SV2V_UNCONNECTED_3074, SV2V_UNCONNECTED_3075, SV2V_UNCONNECTED_3076, SV2V_UNCONNECTED_3077, SV2V_UNCONNECTED_3078, SV2V_UNCONNECTED_3079, SV2V_UNCONNECTED_3080, SV2V_UNCONNECTED_3081, SV2V_UNCONNECTED_3082, SV2V_UNCONNECTED_3083, SV2V_UNCONNECTED_3084, SV2V_UNCONNECTED_3085, SV2V_UNCONNECTED_3086, SV2V_UNCONNECTED_3087, SV2V_UNCONNECTED_3088, SV2V_UNCONNECTED_3089, SV2V_UNCONNECTED_3090, SV2V_UNCONNECTED_3091, SV2V_UNCONNECTED_3092, SV2V_UNCONNECTED_3093, SV2V_UNCONNECTED_3094, SV2V_UNCONNECTED_3095, SV2V_UNCONNECTED_3096, SV2V_UNCONNECTED_3097, SV2V_UNCONNECTED_3098, SV2V_UNCONNECTED_3099, SV2V_UNCONNECTED_3100, SV2V_UNCONNECTED_3101, SV2V_UNCONNECTED_3102, SV2V_UNCONNECTED_3103, SV2V_UNCONNECTED_3104, SV2V_UNCONNECTED_3105, SV2V_UNCONNECTED_3106, SV2V_UNCONNECTED_3107, SV2V_UNCONNECTED_3108, SV2V_UNCONNECTED_3109, SV2V_UNCONNECTED_3110, SV2V_UNCONNECTED_3111, SV2V_UNCONNECTED_3112, SV2V_UNCONNECTED_3113, SV2V_UNCONNECTED_3114, SV2V_UNCONNECTED_3115, SV2V_UNCONNECTED_3116, SV2V_UNCONNECTED_3117, SV2V_UNCONNECTED_3118, SV2V_UNCONNECTED_3119, SV2V_UNCONNECTED_3120, SV2V_UNCONNECTED_3121, SV2V_UNCONNECTED_3122, SV2V_UNCONNECTED_3123, SV2V_UNCONNECTED_3124, SV2V_UNCONNECTED_3125, SV2V_UNCONNECTED_3126, SV2V_UNCONNECTED_3127, SV2V_UNCONNECTED_3128, SV2V_UNCONNECTED_3129, SV2V_UNCONNECTED_3130, SV2V_UNCONNECTED_3131, SV2V_UNCONNECTED_3132, SV2V_UNCONNECTED_3133, SV2V_UNCONNECTED_3134, SV2V_UNCONNECTED_3135, SV2V_UNCONNECTED_3136, SV2V_UNCONNECTED_3137, SV2V_UNCONNECTED_3138, SV2V_UNCONNECTED_3139, SV2V_UNCONNECTED_3140, SV2V_UNCONNECTED_3141, SV2V_UNCONNECTED_3142, SV2V_UNCONNECTED_3143, SV2V_UNCONNECTED_3144, SV2V_UNCONNECTED_3145, SV2V_UNCONNECTED_3146, SV2V_UNCONNECTED_3147, SV2V_UNCONNECTED_3148, SV2V_UNCONNECTED_3149, SV2V_UNCONNECTED_3150, SV2V_UNCONNECTED_3151, SV2V_UNCONNECTED_3152, SV2V_UNCONNECTED_3153, SV2V_UNCONNECTED_3154, SV2V_UNCONNECTED_3155, SV2V_UNCONNECTED_3156, SV2V_UNCONNECTED_3157, SV2V_UNCONNECTED_3158, SV2V_UNCONNECTED_3159, SV2V_UNCONNECTED_3160, SV2V_UNCONNECTED_3161, SV2V_UNCONNECTED_3162, SV2V_UNCONNECTED_3163, SV2V_UNCONNECTED_3164, SV2V_UNCONNECTED_3165, SV2V_UNCONNECTED_3166, SV2V_UNCONNECTED_3167, SV2V_UNCONNECTED_3168, SV2V_UNCONNECTED_3169, SV2V_UNCONNECTED_3170, SV2V_UNCONNECTED_3171, SV2V_UNCONNECTED_3172, SV2V_UNCONNECTED_3173, SV2V_UNCONNECTED_3174, SV2V_UNCONNECTED_3175, SV2V_UNCONNECTED_3176, SV2V_UNCONNECTED_3177, SV2V_UNCONNECTED_3178, SV2V_UNCONNECTED_3179, SV2V_UNCONNECTED_3180, SV2V_UNCONNECTED_3181, SV2V_UNCONNECTED_3182, SV2V_UNCONNECTED_3183, SV2V_UNCONNECTED_3184, SV2V_UNCONNECTED_3185, SV2V_UNCONNECTED_3186, SV2V_UNCONNECTED_3187, SV2V_UNCONNECTED_3188, SV2V_UNCONNECTED_3189, SV2V_UNCONNECTED_3190, SV2V_UNCONNECTED_3191, SV2V_UNCONNECTED_3192, SV2V_UNCONNECTED_3193, SV2V_UNCONNECTED_3194, SV2V_UNCONNECTED_3195, SV2V_UNCONNECTED_3196, SV2V_UNCONNECTED_3197, SV2V_UNCONNECTED_3198, SV2V_UNCONNECTED_3199, SV2V_UNCONNECTED_3200, SV2V_UNCONNECTED_3201, SV2V_UNCONNECTED_3202, SV2V_UNCONNECTED_3203, SV2V_UNCONNECTED_3204, SV2V_UNCONNECTED_3205, SV2V_UNCONNECTED_3206, SV2V_UNCONNECTED_3207, SV2V_UNCONNECTED_3208, SV2V_UNCONNECTED_3209, SV2V_UNCONNECTED_3210, SV2V_UNCONNECTED_3211, SV2V_UNCONNECTED_3212, SV2V_UNCONNECTED_3213, SV2V_UNCONNECTED_3214, SV2V_UNCONNECTED_3215, SV2V_UNCONNECTED_3216, SV2V_UNCONNECTED_3217, SV2V_UNCONNECTED_3218, SV2V_UNCONNECTED_3219, SV2V_UNCONNECTED_3220, SV2V_UNCONNECTED_3221, SV2V_UNCONNECTED_3222, SV2V_UNCONNECTED_3223, SV2V_UNCONNECTED_3224, SV2V_UNCONNECTED_3225, SV2V_UNCONNECTED_3226, SV2V_UNCONNECTED_3227, SV2V_UNCONNECTED_3228, SV2V_UNCONNECTED_3229, SV2V_UNCONNECTED_3230, SV2V_UNCONNECTED_3231, SV2V_UNCONNECTED_3232, SV2V_UNCONNECTED_3233, SV2V_UNCONNECTED_3234, SV2V_UNCONNECTED_3235, SV2V_UNCONNECTED_3236, SV2V_UNCONNECTED_3237, SV2V_UNCONNECTED_3238, SV2V_UNCONNECTED_3239, SV2V_UNCONNECTED_3240, SV2V_UNCONNECTED_3241, SV2V_UNCONNECTED_3242, SV2V_UNCONNECTED_3243, SV2V_UNCONNECTED_3244, SV2V_UNCONNECTED_3245, SV2V_UNCONNECTED_3246, SV2V_UNCONNECTED_3247, SV2V_UNCONNECTED_3248, SV2V_UNCONNECTED_3249, SV2V_UNCONNECTED_3250, SV2V_UNCONNECTED_3251, SV2V_UNCONNECTED_3252, SV2V_UNCONNECTED_3253, SV2V_UNCONNECTED_3254, SV2V_UNCONNECTED_3255, SV2V_UNCONNECTED_3256, SV2V_UNCONNECTED_3257, SV2V_UNCONNECTED_3258, SV2V_UNCONNECTED_3259, SV2V_UNCONNECTED_3260, SV2V_UNCONNECTED_3261, SV2V_UNCONNECTED_3262, SV2V_UNCONNECTED_3263, SV2V_UNCONNECTED_3264, SV2V_UNCONNECTED_3265, SV2V_UNCONNECTED_3266, SV2V_UNCONNECTED_3267, SV2V_UNCONNECTED_3268, SV2V_UNCONNECTED_3269, SV2V_UNCONNECTED_3270, SV2V_UNCONNECTED_3271, SV2V_UNCONNECTED_3272, SV2V_UNCONNECTED_3273, SV2V_UNCONNECTED_3274, SV2V_UNCONNECTED_3275, SV2V_UNCONNECTED_3276, SV2V_UNCONNECTED_3277, SV2V_UNCONNECTED_3278, SV2V_UNCONNECTED_3279, SV2V_UNCONNECTED_3280, SV2V_UNCONNECTED_3281, SV2V_UNCONNECTED_3282, SV2V_UNCONNECTED_3283, SV2V_UNCONNECTED_3284, SV2V_UNCONNECTED_3285, SV2V_UNCONNECTED_3286, SV2V_UNCONNECTED_3287, SV2V_UNCONNECTED_3288, SV2V_UNCONNECTED_3289, SV2V_UNCONNECTED_3290, SV2V_UNCONNECTED_3291, SV2V_UNCONNECTED_3292, SV2V_UNCONNECTED_3293, SV2V_UNCONNECTED_3294, SV2V_UNCONNECTED_3295, SV2V_UNCONNECTED_3296, SV2V_UNCONNECTED_3297, SV2V_UNCONNECTED_3298, SV2V_UNCONNECTED_3299, SV2V_UNCONNECTED_3300, SV2V_UNCONNECTED_3301, SV2V_UNCONNECTED_3302, SV2V_UNCONNECTED_3303, SV2V_UNCONNECTED_3304, SV2V_UNCONNECTED_3305, SV2V_UNCONNECTED_3306, SV2V_UNCONNECTED_3307, SV2V_UNCONNECTED_3308, SV2V_UNCONNECTED_3309, SV2V_UNCONNECTED_3310, SV2V_UNCONNECTED_3311, SV2V_UNCONNECTED_3312, SV2V_UNCONNECTED_3313, SV2V_UNCONNECTED_3314, SV2V_UNCONNECTED_3315, SV2V_UNCONNECTED_3316, SV2V_UNCONNECTED_3317, SV2V_UNCONNECTED_3318, SV2V_UNCONNECTED_3319, SV2V_UNCONNECTED_3320, SV2V_UNCONNECTED_3321, SV2V_UNCONNECTED_3322, SV2V_UNCONNECTED_3323, SV2V_UNCONNECTED_3324, SV2V_UNCONNECTED_3325, SV2V_UNCONNECTED_3326, SV2V_UNCONNECTED_3327, SV2V_UNCONNECTED_3328, SV2V_UNCONNECTED_3329, SV2V_UNCONNECTED_3330, SV2V_UNCONNECTED_3331, SV2V_UNCONNECTED_3332, SV2V_UNCONNECTED_3333, SV2V_UNCONNECTED_3334, SV2V_UNCONNECTED_3335, SV2V_UNCONNECTED_3336, SV2V_UNCONNECTED_3337, SV2V_UNCONNECTED_3338, SV2V_UNCONNECTED_3339, SV2V_UNCONNECTED_3340, SV2V_UNCONNECTED_3341, SV2V_UNCONNECTED_3342, SV2V_UNCONNECTED_3343, SV2V_UNCONNECTED_3344, SV2V_UNCONNECTED_3345, SV2V_UNCONNECTED_3346, SV2V_UNCONNECTED_3347, SV2V_UNCONNECTED_3348, SV2V_UNCONNECTED_3349, SV2V_UNCONNECTED_3350, SV2V_UNCONNECTED_3351, SV2V_UNCONNECTED_3352, SV2V_UNCONNECTED_3353, SV2V_UNCONNECTED_3354, SV2V_UNCONNECTED_3355, SV2V_UNCONNECTED_3356, SV2V_UNCONNECTED_3357, SV2V_UNCONNECTED_3358, SV2V_UNCONNECTED_3359, SV2V_UNCONNECTED_3360, SV2V_UNCONNECTED_3361, SV2V_UNCONNECTED_3362, SV2V_UNCONNECTED_3363, SV2V_UNCONNECTED_3364, SV2V_UNCONNECTED_3365, SV2V_UNCONNECTED_3366, SV2V_UNCONNECTED_3367, SV2V_UNCONNECTED_3368, SV2V_UNCONNECTED_3369, SV2V_UNCONNECTED_3370, SV2V_UNCONNECTED_3371, SV2V_UNCONNECTED_3372, SV2V_UNCONNECTED_3373, SV2V_UNCONNECTED_3374, SV2V_UNCONNECTED_3375, SV2V_UNCONNECTED_3376, SV2V_UNCONNECTED_3377, SV2V_UNCONNECTED_3378, SV2V_UNCONNECTED_3379, SV2V_UNCONNECTED_3380, SV2V_UNCONNECTED_3381, SV2V_UNCONNECTED_3382, SV2V_UNCONNECTED_3383, SV2V_UNCONNECTED_3384, SV2V_UNCONNECTED_3385, SV2V_UNCONNECTED_3386, SV2V_UNCONNECTED_3387, SV2V_UNCONNECTED_3388, SV2V_UNCONNECTED_3389, SV2V_UNCONNECTED_3390, SV2V_UNCONNECTED_3391, SV2V_UNCONNECTED_3392, SV2V_UNCONNECTED_3393, SV2V_UNCONNECTED_3394, SV2V_UNCONNECTED_3395, SV2V_UNCONNECTED_3396, SV2V_UNCONNECTED_3397, SV2V_UNCONNECTED_3398, SV2V_UNCONNECTED_3399, SV2V_UNCONNECTED_3400, SV2V_UNCONNECTED_3401, SV2V_UNCONNECTED_3402, SV2V_UNCONNECTED_3403, SV2V_UNCONNECTED_3404, SV2V_UNCONNECTED_3405, SV2V_UNCONNECTED_3406, SV2V_UNCONNECTED_3407, SV2V_UNCONNECTED_3408, SV2V_UNCONNECTED_3409, SV2V_UNCONNECTED_3410, SV2V_UNCONNECTED_3411, SV2V_UNCONNECTED_3412, SV2V_UNCONNECTED_3413, SV2V_UNCONNECTED_3414, SV2V_UNCONNECTED_3415, SV2V_UNCONNECTED_3416, SV2V_UNCONNECTED_3417, SV2V_UNCONNECTED_3418, SV2V_UNCONNECTED_3419, SV2V_UNCONNECTED_3420, SV2V_UNCONNECTED_3421, SV2V_UNCONNECTED_3422, SV2V_UNCONNECTED_3423, SV2V_UNCONNECTED_3424, SV2V_UNCONNECTED_3425, SV2V_UNCONNECTED_3426, SV2V_UNCONNECTED_3427, SV2V_UNCONNECTED_3428, SV2V_UNCONNECTED_3429, SV2V_UNCONNECTED_3430, SV2V_UNCONNECTED_3431, SV2V_UNCONNECTED_3432, SV2V_UNCONNECTED_3433, SV2V_UNCONNECTED_3434, SV2V_UNCONNECTED_3435, SV2V_UNCONNECTED_3436, SV2V_UNCONNECTED_3437, SV2V_UNCONNECTED_3438, SV2V_UNCONNECTED_3439, SV2V_UNCONNECTED_3440, SV2V_UNCONNECTED_3441, SV2V_UNCONNECTED_3442, SV2V_UNCONNECTED_3443, SV2V_UNCONNECTED_3444, SV2V_UNCONNECTED_3445, SV2V_UNCONNECTED_3446, SV2V_UNCONNECTED_3447, SV2V_UNCONNECTED_3448, SV2V_UNCONNECTED_3449, SV2V_UNCONNECTED_3450, SV2V_UNCONNECTED_3451, SV2V_UNCONNECTED_3452, SV2V_UNCONNECTED_3453, SV2V_UNCONNECTED_3454, SV2V_UNCONNECTED_3455, SV2V_UNCONNECTED_3456, SV2V_UNCONNECTED_3457, SV2V_UNCONNECTED_3458, SV2V_UNCONNECTED_3459, SV2V_UNCONNECTED_3460, SV2V_UNCONNECTED_3461, SV2V_UNCONNECTED_3462, SV2V_UNCONNECTED_3463, SV2V_UNCONNECTED_3464, SV2V_UNCONNECTED_3465, SV2V_UNCONNECTED_3466, SV2V_UNCONNECTED_3467, SV2V_UNCONNECTED_3468, SV2V_UNCONNECTED_3469, SV2V_UNCONNECTED_3470, SV2V_UNCONNECTED_3471, SV2V_UNCONNECTED_3472, SV2V_UNCONNECTED_3473, SV2V_UNCONNECTED_3474, SV2V_UNCONNECTED_3475, SV2V_UNCONNECTED_3476, SV2V_UNCONNECTED_3477, SV2V_UNCONNECTED_3478, SV2V_UNCONNECTED_3479, SV2V_UNCONNECTED_3480, SV2V_UNCONNECTED_3481, SV2V_UNCONNECTED_3482, SV2V_UNCONNECTED_3483, SV2V_UNCONNECTED_3484, SV2V_UNCONNECTED_3485, SV2V_UNCONNECTED_3486, SV2V_UNCONNECTED_3487, SV2V_UNCONNECTED_3488, SV2V_UNCONNECTED_3489, SV2V_UNCONNECTED_3490, SV2V_UNCONNECTED_3491, SV2V_UNCONNECTED_3492, SV2V_UNCONNECTED_3493, SV2V_UNCONNECTED_3494, SV2V_UNCONNECTED_3495, SV2V_UNCONNECTED_3496, SV2V_UNCONNECTED_3497, SV2V_UNCONNECTED_3498, SV2V_UNCONNECTED_3499, SV2V_UNCONNECTED_3500, SV2V_UNCONNECTED_3501, SV2V_UNCONNECTED_3502, SV2V_UNCONNECTED_3503, SV2V_UNCONNECTED_3504, SV2V_UNCONNECTED_3505, SV2V_UNCONNECTED_3506, SV2V_UNCONNECTED_3507, SV2V_UNCONNECTED_3508, SV2V_UNCONNECTED_3509, SV2V_UNCONNECTED_3510, SV2V_UNCONNECTED_3511, SV2V_UNCONNECTED_3512, SV2V_UNCONNECTED_3513, SV2V_UNCONNECTED_3514, SV2V_UNCONNECTED_3515, SV2V_UNCONNECTED_3516, SV2V_UNCONNECTED_3517, SV2V_UNCONNECTED_3518, SV2V_UNCONNECTED_3519, SV2V_UNCONNECTED_3520, SV2V_UNCONNECTED_3521, SV2V_UNCONNECTED_3522, SV2V_UNCONNECTED_3523, SV2V_UNCONNECTED_3524, SV2V_UNCONNECTED_3525, SV2V_UNCONNECTED_3526, SV2V_UNCONNECTED_3527, SV2V_UNCONNECTED_3528, SV2V_UNCONNECTED_3529, SV2V_UNCONNECTED_3530, SV2V_UNCONNECTED_3531, SV2V_UNCONNECTED_3532, SV2V_UNCONNECTED_3533, SV2V_UNCONNECTED_3534, SV2V_UNCONNECTED_3535, SV2V_UNCONNECTED_3536, SV2V_UNCONNECTED_3537, SV2V_UNCONNECTED_3538, SV2V_UNCONNECTED_3539, SV2V_UNCONNECTED_3540, SV2V_UNCONNECTED_3541, SV2V_UNCONNECTED_3542, SV2V_UNCONNECTED_3543, SV2V_UNCONNECTED_3544, SV2V_UNCONNECTED_3545, SV2V_UNCONNECTED_3546, SV2V_UNCONNECTED_3547, SV2V_UNCONNECTED_3548, SV2V_UNCONNECTED_3549, SV2V_UNCONNECTED_3550, SV2V_UNCONNECTED_3551, SV2V_UNCONNECTED_3552, SV2V_UNCONNECTED_3553, SV2V_UNCONNECTED_3554, SV2V_UNCONNECTED_3555, SV2V_UNCONNECTED_3556, SV2V_UNCONNECTED_3557, SV2V_UNCONNECTED_3558, SV2V_UNCONNECTED_3559, SV2V_UNCONNECTED_3560, SV2V_UNCONNECTED_3561, SV2V_UNCONNECTED_3562, SV2V_UNCONNECTED_3563, SV2V_UNCONNECTED_3564, SV2V_UNCONNECTED_3565, SV2V_UNCONNECTED_3566, SV2V_UNCONNECTED_3567, SV2V_UNCONNECTED_3568, SV2V_UNCONNECTED_3569, SV2V_UNCONNECTED_3570, SV2V_UNCONNECTED_3571, SV2V_UNCONNECTED_3572, SV2V_UNCONNECTED_3573, SV2V_UNCONNECTED_3574, SV2V_UNCONNECTED_3575, SV2V_UNCONNECTED_3576, SV2V_UNCONNECTED_3577, SV2V_UNCONNECTED_3578, SV2V_UNCONNECTED_3579, SV2V_UNCONNECTED_3580, SV2V_UNCONNECTED_3581, SV2V_UNCONNECTED_3582, SV2V_UNCONNECTED_3583, SV2V_UNCONNECTED_3584, SV2V_UNCONNECTED_3585, SV2V_UNCONNECTED_3586, SV2V_UNCONNECTED_3587, SV2V_UNCONNECTED_3588, SV2V_UNCONNECTED_3589, SV2V_UNCONNECTED_3590, SV2V_UNCONNECTED_3591, SV2V_UNCONNECTED_3592, SV2V_UNCONNECTED_3593, SV2V_UNCONNECTED_3594, SV2V_UNCONNECTED_3595, SV2V_UNCONNECTED_3596, SV2V_UNCONNECTED_3597, SV2V_UNCONNECTED_3598, SV2V_UNCONNECTED_3599, SV2V_UNCONNECTED_3600, SV2V_UNCONNECTED_3601, SV2V_UNCONNECTED_3602, SV2V_UNCONNECTED_3603, SV2V_UNCONNECTED_3604, SV2V_UNCONNECTED_3605, SV2V_UNCONNECTED_3606, SV2V_UNCONNECTED_3607, SV2V_UNCONNECTED_3608, SV2V_UNCONNECTED_3609, SV2V_UNCONNECTED_3610, SV2V_UNCONNECTED_3611, SV2V_UNCONNECTED_3612, SV2V_UNCONNECTED_3613, SV2V_UNCONNECTED_3614, SV2V_UNCONNECTED_3615, SV2V_UNCONNECTED_3616, SV2V_UNCONNECTED_3617, SV2V_UNCONNECTED_3618, SV2V_UNCONNECTED_3619, SV2V_UNCONNECTED_3620, SV2V_UNCONNECTED_3621, SV2V_UNCONNECTED_3622, SV2V_UNCONNECTED_3623, SV2V_UNCONNECTED_3624, SV2V_UNCONNECTED_3625, SV2V_UNCONNECTED_3626, SV2V_UNCONNECTED_3627, SV2V_UNCONNECTED_3628, SV2V_UNCONNECTED_3629, SV2V_UNCONNECTED_3630, SV2V_UNCONNECTED_3631, SV2V_UNCONNECTED_3632, SV2V_UNCONNECTED_3633, SV2V_UNCONNECTED_3634, SV2V_UNCONNECTED_3635, SV2V_UNCONNECTED_3636, SV2V_UNCONNECTED_3637, SV2V_UNCONNECTED_3638, SV2V_UNCONNECTED_3639, SV2V_UNCONNECTED_3640, SV2V_UNCONNECTED_3641, SV2V_UNCONNECTED_3642, SV2V_UNCONNECTED_3643, SV2V_UNCONNECTED_3644, SV2V_UNCONNECTED_3645, SV2V_UNCONNECTED_3646, SV2V_UNCONNECTED_3647, SV2V_UNCONNECTED_3648, SV2V_UNCONNECTED_3649, SV2V_UNCONNECTED_3650, SV2V_UNCONNECTED_3651, SV2V_UNCONNECTED_3652, SV2V_UNCONNECTED_3653, SV2V_UNCONNECTED_3654, SV2V_UNCONNECTED_3655, SV2V_UNCONNECTED_3656, SV2V_UNCONNECTED_3657, SV2V_UNCONNECTED_3658, SV2V_UNCONNECTED_3659, SV2V_UNCONNECTED_3660, SV2V_UNCONNECTED_3661, SV2V_UNCONNECTED_3662, SV2V_UNCONNECTED_3663, SV2V_UNCONNECTED_3664, SV2V_UNCONNECTED_3665, SV2V_UNCONNECTED_3666, SV2V_UNCONNECTED_3667, SV2V_UNCONNECTED_3668, SV2V_UNCONNECTED_3669, SV2V_UNCONNECTED_3670, SV2V_UNCONNECTED_3671, SV2V_UNCONNECTED_3672, SV2V_UNCONNECTED_3673, SV2V_UNCONNECTED_3674, SV2V_UNCONNECTED_3675, SV2V_UNCONNECTED_3676, SV2V_UNCONNECTED_3677, SV2V_UNCONNECTED_3678, SV2V_UNCONNECTED_3679, SV2V_UNCONNECTED_3680, SV2V_UNCONNECTED_3681, SV2V_UNCONNECTED_3682, SV2V_UNCONNECTED_3683, SV2V_UNCONNECTED_3684, SV2V_UNCONNECTED_3685, SV2V_UNCONNECTED_3686, SV2V_UNCONNECTED_3687, SV2V_UNCONNECTED_3688, SV2V_UNCONNECTED_3689, SV2V_UNCONNECTED_3690, SV2V_UNCONNECTED_3691, SV2V_UNCONNECTED_3692, SV2V_UNCONNECTED_3693, SV2V_UNCONNECTED_3694, SV2V_UNCONNECTED_3695, SV2V_UNCONNECTED_3696, SV2V_UNCONNECTED_3697, SV2V_UNCONNECTED_3698, SV2V_UNCONNECTED_3699, SV2V_UNCONNECTED_3700, SV2V_UNCONNECTED_3701, SV2V_UNCONNECTED_3702, SV2V_UNCONNECTED_3703, SV2V_UNCONNECTED_3704, SV2V_UNCONNECTED_3705, SV2V_UNCONNECTED_3706, SV2V_UNCONNECTED_3707, SV2V_UNCONNECTED_3708, SV2V_UNCONNECTED_3709, SV2V_UNCONNECTED_3710, SV2V_UNCONNECTED_3711, SV2V_UNCONNECTED_3712, SV2V_UNCONNECTED_3713, SV2V_UNCONNECTED_3714, SV2V_UNCONNECTED_3715, SV2V_UNCONNECTED_3716, SV2V_UNCONNECTED_3717, SV2V_UNCONNECTED_3718, SV2V_UNCONNECTED_3719, SV2V_UNCONNECTED_3720, SV2V_UNCONNECTED_3721, SV2V_UNCONNECTED_3722, SV2V_UNCONNECTED_3723, SV2V_UNCONNECTED_3724, SV2V_UNCONNECTED_3725, SV2V_UNCONNECTED_3726, SV2V_UNCONNECTED_3727, SV2V_UNCONNECTED_3728, SV2V_UNCONNECTED_3729, SV2V_UNCONNECTED_3730, SV2V_UNCONNECTED_3731, SV2V_UNCONNECTED_3732, SV2V_UNCONNECTED_3733, SV2V_UNCONNECTED_3734, SV2V_UNCONNECTED_3735, SV2V_UNCONNECTED_3736, SV2V_UNCONNECTED_3737, SV2V_UNCONNECTED_3738, SV2V_UNCONNECTED_3739, SV2V_UNCONNECTED_3740, SV2V_UNCONNECTED_3741, SV2V_UNCONNECTED_3742, SV2V_UNCONNECTED_3743, SV2V_UNCONNECTED_3744, SV2V_UNCONNECTED_3745, SV2V_UNCONNECTED_3746, SV2V_UNCONNECTED_3747, SV2V_UNCONNECTED_3748, SV2V_UNCONNECTED_3749, SV2V_UNCONNECTED_3750, SV2V_UNCONNECTED_3751, SV2V_UNCONNECTED_3752, SV2V_UNCONNECTED_3753, SV2V_UNCONNECTED_3754, SV2V_UNCONNECTED_3755, SV2V_UNCONNECTED_3756, SV2V_UNCONNECTED_3757, SV2V_UNCONNECTED_3758, SV2V_UNCONNECTED_3759, SV2V_UNCONNECTED_3760, SV2V_UNCONNECTED_3761, SV2V_UNCONNECTED_3762, SV2V_UNCONNECTED_3763, SV2V_UNCONNECTED_3764, SV2V_UNCONNECTED_3765, SV2V_UNCONNECTED_3766, SV2V_UNCONNECTED_3767, SV2V_UNCONNECTED_3768, SV2V_UNCONNECTED_3769, SV2V_UNCONNECTED_3770, SV2V_UNCONNECTED_3771, SV2V_UNCONNECTED_3772, SV2V_UNCONNECTED_3773, SV2V_UNCONNECTED_3774, SV2V_UNCONNECTED_3775, SV2V_UNCONNECTED_3776, SV2V_UNCONNECTED_3777, SV2V_UNCONNECTED_3778, SV2V_UNCONNECTED_3779, SV2V_UNCONNECTED_3780, SV2V_UNCONNECTED_3781, SV2V_UNCONNECTED_3782, SV2V_UNCONNECTED_3783, SV2V_UNCONNECTED_3784, SV2V_UNCONNECTED_3785, SV2V_UNCONNECTED_3786, SV2V_UNCONNECTED_3787, SV2V_UNCONNECTED_3788, SV2V_UNCONNECTED_3789, SV2V_UNCONNECTED_3790, SV2V_UNCONNECTED_3791, SV2V_UNCONNECTED_3792, SV2V_UNCONNECTED_3793, SV2V_UNCONNECTED_3794, SV2V_UNCONNECTED_3795, SV2V_UNCONNECTED_3796, SV2V_UNCONNECTED_3797, SV2V_UNCONNECTED_3798, SV2V_UNCONNECTED_3799, SV2V_UNCONNECTED_3800, SV2V_UNCONNECTED_3801, SV2V_UNCONNECTED_3802, SV2V_UNCONNECTED_3803, SV2V_UNCONNECTED_3804, SV2V_UNCONNECTED_3805, SV2V_UNCONNECTED_3806, SV2V_UNCONNECTED_3807, SV2V_UNCONNECTED_3808, SV2V_UNCONNECTED_3809, SV2V_UNCONNECTED_3810, SV2V_UNCONNECTED_3811, SV2V_UNCONNECTED_3812, SV2V_UNCONNECTED_3813, SV2V_UNCONNECTED_3814, SV2V_UNCONNECTED_3815, SV2V_UNCONNECTED_3816, SV2V_UNCONNECTED_3817, SV2V_UNCONNECTED_3818, SV2V_UNCONNECTED_3819, SV2V_UNCONNECTED_3820, SV2V_UNCONNECTED_3821, SV2V_UNCONNECTED_3822, SV2V_UNCONNECTED_3823, SV2V_UNCONNECTED_3824, SV2V_UNCONNECTED_3825, SV2V_UNCONNECTED_3826, SV2V_UNCONNECTED_3827, SV2V_UNCONNECTED_3828, SV2V_UNCONNECTED_3829, SV2V_UNCONNECTED_3830, SV2V_UNCONNECTED_3831, SV2V_UNCONNECTED_3832, SV2V_UNCONNECTED_3833, SV2V_UNCONNECTED_3834, SV2V_UNCONNECTED_3835, SV2V_UNCONNECTED_3836, SV2V_UNCONNECTED_3837, SV2V_UNCONNECTED_3838, SV2V_UNCONNECTED_3839, SV2V_UNCONNECTED_3840, SV2V_UNCONNECTED_3841, SV2V_UNCONNECTED_3842, SV2V_UNCONNECTED_3843, SV2V_UNCONNECTED_3844, SV2V_UNCONNECTED_3845, SV2V_UNCONNECTED_3846, SV2V_UNCONNECTED_3847, SV2V_UNCONNECTED_3848, SV2V_UNCONNECTED_3849, SV2V_UNCONNECTED_3850, SV2V_UNCONNECTED_3851, SV2V_UNCONNECTED_3852, SV2V_UNCONNECTED_3853, SV2V_UNCONNECTED_3854, SV2V_UNCONNECTED_3855, SV2V_UNCONNECTED_3856, SV2V_UNCONNECTED_3857, SV2V_UNCONNECTED_3858, SV2V_UNCONNECTED_3859, SV2V_UNCONNECTED_3860, SV2V_UNCONNECTED_3861, SV2V_UNCONNECTED_3862, SV2V_UNCONNECTED_3863, SV2V_UNCONNECTED_3864, SV2V_UNCONNECTED_3865, SV2V_UNCONNECTED_3866, SV2V_UNCONNECTED_3867, SV2V_UNCONNECTED_3868, SV2V_UNCONNECTED_3869, SV2V_UNCONNECTED_3870, SV2V_UNCONNECTED_3871, SV2V_UNCONNECTED_3872, SV2V_UNCONNECTED_3873, SV2V_UNCONNECTED_3874, SV2V_UNCONNECTED_3875, SV2V_UNCONNECTED_3876, SV2V_UNCONNECTED_3877, SV2V_UNCONNECTED_3878, SV2V_UNCONNECTED_3879, SV2V_UNCONNECTED_3880, SV2V_UNCONNECTED_3881, SV2V_UNCONNECTED_3882, SV2V_UNCONNECTED_3883, SV2V_UNCONNECTED_3884, SV2V_UNCONNECTED_3885, SV2V_UNCONNECTED_3886, SV2V_UNCONNECTED_3887, SV2V_UNCONNECTED_3888, SV2V_UNCONNECTED_3889, SV2V_UNCONNECTED_3890, SV2V_UNCONNECTED_3891, SV2V_UNCONNECTED_3892, SV2V_UNCONNECTED_3893, SV2V_UNCONNECTED_3894, SV2V_UNCONNECTED_3895, SV2V_UNCONNECTED_3896, SV2V_UNCONNECTED_3897, SV2V_UNCONNECTED_3898, SV2V_UNCONNECTED_3899, SV2V_UNCONNECTED_3900, SV2V_UNCONNECTED_3901, SV2V_UNCONNECTED_3902, SV2V_UNCONNECTED_3903, SV2V_UNCONNECTED_3904, SV2V_UNCONNECTED_3905, SV2V_UNCONNECTED_3906, SV2V_UNCONNECTED_3907, SV2V_UNCONNECTED_3908, SV2V_UNCONNECTED_3909, SV2V_UNCONNECTED_3910, SV2V_UNCONNECTED_3911, SV2V_UNCONNECTED_3912, SV2V_UNCONNECTED_3913, SV2V_UNCONNECTED_3914, SV2V_UNCONNECTED_3915, SV2V_UNCONNECTED_3916, SV2V_UNCONNECTED_3917, SV2V_UNCONNECTED_3918, SV2V_UNCONNECTED_3919, SV2V_UNCONNECTED_3920, SV2V_UNCONNECTED_3921, SV2V_UNCONNECTED_3922, SV2V_UNCONNECTED_3923, SV2V_UNCONNECTED_3924, SV2V_UNCONNECTED_3925, SV2V_UNCONNECTED_3926, SV2V_UNCONNECTED_3927, SV2V_UNCONNECTED_3928, SV2V_UNCONNECTED_3929, SV2V_UNCONNECTED_3930, SV2V_UNCONNECTED_3931, SV2V_UNCONNECTED_3932, SV2V_UNCONNECTED_3933, SV2V_UNCONNECTED_3934, SV2V_UNCONNECTED_3935, SV2V_UNCONNECTED_3936, SV2V_UNCONNECTED_3937, SV2V_UNCONNECTED_3938, SV2V_UNCONNECTED_3939, SV2V_UNCONNECTED_3940, SV2V_UNCONNECTED_3941, SV2V_UNCONNECTED_3942, SV2V_UNCONNECTED_3943, SV2V_UNCONNECTED_3944, SV2V_UNCONNECTED_3945, SV2V_UNCONNECTED_3946, SV2V_UNCONNECTED_3947, SV2V_UNCONNECTED_3948, SV2V_UNCONNECTED_3949, SV2V_UNCONNECTED_3950, SV2V_UNCONNECTED_3951, SV2V_UNCONNECTED_3952, SV2V_UNCONNECTED_3953, SV2V_UNCONNECTED_3954, SV2V_UNCONNECTED_3955, SV2V_UNCONNECTED_3956, SV2V_UNCONNECTED_3957, SV2V_UNCONNECTED_3958, SV2V_UNCONNECTED_3959, SV2V_UNCONNECTED_3960, SV2V_UNCONNECTED_3961, SV2V_UNCONNECTED_3962, SV2V_UNCONNECTED_3963, SV2V_UNCONNECTED_3964, SV2V_UNCONNECTED_3965, SV2V_UNCONNECTED_3966, SV2V_UNCONNECTED_3967, SV2V_UNCONNECTED_3968, SV2V_UNCONNECTED_3969, SV2V_UNCONNECTED_3970, SV2V_UNCONNECTED_3971, SV2V_UNCONNECTED_3972, SV2V_UNCONNECTED_3973, SV2V_UNCONNECTED_3974, SV2V_UNCONNECTED_3975, SV2V_UNCONNECTED_3976, SV2V_UNCONNECTED_3977, SV2V_UNCONNECTED_3978, SV2V_UNCONNECTED_3979, SV2V_UNCONNECTED_3980, SV2V_UNCONNECTED_3981, SV2V_UNCONNECTED_3982, SV2V_UNCONNECTED_3983, SV2V_UNCONNECTED_3984, SV2V_UNCONNECTED_3985, SV2V_UNCONNECTED_3986, SV2V_UNCONNECTED_3987, SV2V_UNCONNECTED_3988, SV2V_UNCONNECTED_3989, SV2V_UNCONNECTED_3990, SV2V_UNCONNECTED_3991, SV2V_UNCONNECTED_3992, SV2V_UNCONNECTED_3993, SV2V_UNCONNECTED_3994, SV2V_UNCONNECTED_3995, SV2V_UNCONNECTED_3996, SV2V_UNCONNECTED_3997, SV2V_UNCONNECTED_3998, SV2V_UNCONNECTED_3999, SV2V_UNCONNECTED_4000, SV2V_UNCONNECTED_4001, SV2V_UNCONNECTED_4002, SV2V_UNCONNECTED_4003, SV2V_UNCONNECTED_4004, SV2V_UNCONNECTED_4005, SV2V_UNCONNECTED_4006, SV2V_UNCONNECTED_4007, SV2V_UNCONNECTED_4008, SV2V_UNCONNECTED_4009, SV2V_UNCONNECTED_4010, SV2V_UNCONNECTED_4011, SV2V_UNCONNECTED_4012, SV2V_UNCONNECTED_4013, SV2V_UNCONNECTED_4014, SV2V_UNCONNECTED_4015, SV2V_UNCONNECTED_4016, SV2V_UNCONNECTED_4017, SV2V_UNCONNECTED_4018, SV2V_UNCONNECTED_4019, SV2V_UNCONNECTED_4020, SV2V_UNCONNECTED_4021, SV2V_UNCONNECTED_4022, SV2V_UNCONNECTED_4023, SV2V_UNCONNECTED_4024, SV2V_UNCONNECTED_4025, SV2V_UNCONNECTED_4026, SV2V_UNCONNECTED_4027, SV2V_UNCONNECTED_4028, SV2V_UNCONNECTED_4029, SV2V_UNCONNECTED_4030, SV2V_UNCONNECTED_4031, SV2V_UNCONNECTED_4032, SV2V_UNCONNECTED_4033, SV2V_UNCONNECTED_4034, SV2V_UNCONNECTED_4035, SV2V_UNCONNECTED_4036, SV2V_UNCONNECTED_4037, SV2V_UNCONNECTED_4038, SV2V_UNCONNECTED_4039, SV2V_UNCONNECTED_4040, SV2V_UNCONNECTED_4041, SV2V_UNCONNECTED_4042, SV2V_UNCONNECTED_4043, SV2V_UNCONNECTED_4044, SV2V_UNCONNECTED_4045, SV2V_UNCONNECTED_4046, SV2V_UNCONNECTED_4047, SV2V_UNCONNECTED_4048, SV2V_UNCONNECTED_4049, SV2V_UNCONNECTED_4050, SV2V_UNCONNECTED_4051, SV2V_UNCONNECTED_4052, SV2V_UNCONNECTED_4053, SV2V_UNCONNECTED_4054, SV2V_UNCONNECTED_4055, SV2V_UNCONNECTED_4056, SV2V_UNCONNECTED_4057, SV2V_UNCONNECTED_4058, SV2V_UNCONNECTED_4059, SV2V_UNCONNECTED_4060, SV2V_UNCONNECTED_4061, SV2V_UNCONNECTED_4062, SV2V_UNCONNECTED_4063, SV2V_UNCONNECTED_4064, SV2V_UNCONNECTED_4065, SV2V_UNCONNECTED_4066, SV2V_UNCONNECTED_4067, SV2V_UNCONNECTED_4068, SV2V_UNCONNECTED_4069, SV2V_UNCONNECTED_4070, SV2V_UNCONNECTED_4071, SV2V_UNCONNECTED_4072, SV2V_UNCONNECTED_4073, SV2V_UNCONNECTED_4074, SV2V_UNCONNECTED_4075, SV2V_UNCONNECTED_4076, SV2V_UNCONNECTED_4077, SV2V_UNCONNECTED_4078, SV2V_UNCONNECTED_4079, SV2V_UNCONNECTED_4080, SV2V_UNCONNECTED_4081, SV2V_UNCONNECTED_4082, SV2V_UNCONNECTED_4083, SV2V_UNCONNECTED_4084, SV2V_UNCONNECTED_4085, SV2V_UNCONNECTED_4086, SV2V_UNCONNECTED_4087, SV2V_UNCONNECTED_4088, SV2V_UNCONNECTED_4089, SV2V_UNCONNECTED_4090, SV2V_UNCONNECTED_4091, SV2V_UNCONNECTED_4092, SV2V_UNCONNECTED_4093, SV2V_UNCONNECTED_4094, SV2V_UNCONNECTED_4095, SV2V_UNCONNECTED_4096, SV2V_UNCONNECTED_4097, SV2V_UNCONNECTED_4098, SV2V_UNCONNECTED_4099, SV2V_UNCONNECTED_4100, SV2V_UNCONNECTED_4101, SV2V_UNCONNECTED_4102, SV2V_UNCONNECTED_4103, SV2V_UNCONNECTED_4104, SV2V_UNCONNECTED_4105, SV2V_UNCONNECTED_4106, SV2V_UNCONNECTED_4107, SV2V_UNCONNECTED_4108, SV2V_UNCONNECTED_4109, SV2V_UNCONNECTED_4110, SV2V_UNCONNECTED_4111, SV2V_UNCONNECTED_4112, SV2V_UNCONNECTED_4113, SV2V_UNCONNECTED_4114, SV2V_UNCONNECTED_4115, SV2V_UNCONNECTED_4116, SV2V_UNCONNECTED_4117, SV2V_UNCONNECTED_4118, SV2V_UNCONNECTED_4119, SV2V_UNCONNECTED_4120, SV2V_UNCONNECTED_4121, SV2V_UNCONNECTED_4122, SV2V_UNCONNECTED_4123, SV2V_UNCONNECTED_4124, SV2V_UNCONNECTED_4125, SV2V_UNCONNECTED_4126, SV2V_UNCONNECTED_4127, SV2V_UNCONNECTED_4128, SV2V_UNCONNECTED_4129, SV2V_UNCONNECTED_4130, SV2V_UNCONNECTED_4131, SV2V_UNCONNECTED_4132, SV2V_UNCONNECTED_4133, SV2V_UNCONNECTED_4134, SV2V_UNCONNECTED_4135, SV2V_UNCONNECTED_4136, SV2V_UNCONNECTED_4137, SV2V_UNCONNECTED_4138, SV2V_UNCONNECTED_4139, SV2V_UNCONNECTED_4140, SV2V_UNCONNECTED_4141, SV2V_UNCONNECTED_4142, SV2V_UNCONNECTED_4143, SV2V_UNCONNECTED_4144, SV2V_UNCONNECTED_4145, SV2V_UNCONNECTED_4146, SV2V_UNCONNECTED_4147, SV2V_UNCONNECTED_4148, SV2V_UNCONNECTED_4149, SV2V_UNCONNECTED_4150, SV2V_UNCONNECTED_4151, SV2V_UNCONNECTED_4152, SV2V_UNCONNECTED_4153, SV2V_UNCONNECTED_4154, SV2V_UNCONNECTED_4155, SV2V_UNCONNECTED_4156, SV2V_UNCONNECTED_4157, SV2V_UNCONNECTED_4158, SV2V_UNCONNECTED_4159, SV2V_UNCONNECTED_4160, SV2V_UNCONNECTED_4161, SV2V_UNCONNECTED_4162, SV2V_UNCONNECTED_4163, SV2V_UNCONNECTED_4164, SV2V_UNCONNECTED_4165, SV2V_UNCONNECTED_4166, SV2V_UNCONNECTED_4167, SV2V_UNCONNECTED_4168, SV2V_UNCONNECTED_4169, SV2V_UNCONNECTED_4170, SV2V_UNCONNECTED_4171, SV2V_UNCONNECTED_4172, SV2V_UNCONNECTED_4173, SV2V_UNCONNECTED_4174, SV2V_UNCONNECTED_4175, SV2V_UNCONNECTED_4176, SV2V_UNCONNECTED_4177, SV2V_UNCONNECTED_4178, SV2V_UNCONNECTED_4179, SV2V_UNCONNECTED_4180, SV2V_UNCONNECTED_4181, SV2V_UNCONNECTED_4182, SV2V_UNCONNECTED_4183, SV2V_UNCONNECTED_4184, SV2V_UNCONNECTED_4185, SV2V_UNCONNECTED_4186, SV2V_UNCONNECTED_4187, SV2V_UNCONNECTED_4188, SV2V_UNCONNECTED_4189, SV2V_UNCONNECTED_4190, SV2V_UNCONNECTED_4191, SV2V_UNCONNECTED_4192, SV2V_UNCONNECTED_4193, SV2V_UNCONNECTED_4194, SV2V_UNCONNECTED_4195, SV2V_UNCONNECTED_4196, SV2V_UNCONNECTED_4197, SV2V_UNCONNECTED_4198, SV2V_UNCONNECTED_4199, SV2V_UNCONNECTED_4200, SV2V_UNCONNECTED_4201, SV2V_UNCONNECTED_4202, SV2V_UNCONNECTED_4203, SV2V_UNCONNECTED_4204, SV2V_UNCONNECTED_4205, SV2V_UNCONNECTED_4206, SV2V_UNCONNECTED_4207, SV2V_UNCONNECTED_4208, SV2V_UNCONNECTED_4209, SV2V_UNCONNECTED_4210, SV2V_UNCONNECTED_4211, SV2V_UNCONNECTED_4212, SV2V_UNCONNECTED_4213, SV2V_UNCONNECTED_4214, SV2V_UNCONNECTED_4215, SV2V_UNCONNECTED_4216, SV2V_UNCONNECTED_4217, SV2V_UNCONNECTED_4218, SV2V_UNCONNECTED_4219, SV2V_UNCONNECTED_4220, SV2V_UNCONNECTED_4221, SV2V_UNCONNECTED_4222, SV2V_UNCONNECTED_4223, SV2V_UNCONNECTED_4224, SV2V_UNCONNECTED_4225, SV2V_UNCONNECTED_4226, SV2V_UNCONNECTED_4227, SV2V_UNCONNECTED_4228, SV2V_UNCONNECTED_4229, SV2V_UNCONNECTED_4230, SV2V_UNCONNECTED_4231, SV2V_UNCONNECTED_4232, SV2V_UNCONNECTED_4233, SV2V_UNCONNECTED_4234, SV2V_UNCONNECTED_4235, SV2V_UNCONNECTED_4236, SV2V_UNCONNECTED_4237, SV2V_UNCONNECTED_4238, SV2V_UNCONNECTED_4239, SV2V_UNCONNECTED_4240, SV2V_UNCONNECTED_4241, SV2V_UNCONNECTED_4242, SV2V_UNCONNECTED_4243, SV2V_UNCONNECTED_4244, SV2V_UNCONNECTED_4245, SV2V_UNCONNECTED_4246, SV2V_UNCONNECTED_4247, SV2V_UNCONNECTED_4248, SV2V_UNCONNECTED_4249, SV2V_UNCONNECTED_4250, SV2V_UNCONNECTED_4251, SV2V_UNCONNECTED_4252, SV2V_UNCONNECTED_4253, SV2V_UNCONNECTED_4254, SV2V_UNCONNECTED_4255, SV2V_UNCONNECTED_4256, SV2V_UNCONNECTED_4257, SV2V_UNCONNECTED_4258, SV2V_UNCONNECTED_4259, SV2V_UNCONNECTED_4260, SV2V_UNCONNECTED_4261, SV2V_UNCONNECTED_4262, SV2V_UNCONNECTED_4263, SV2V_UNCONNECTED_4264, SV2V_UNCONNECTED_4265, SV2V_UNCONNECTED_4266, SV2V_UNCONNECTED_4267, SV2V_UNCONNECTED_4268, SV2V_UNCONNECTED_4269, SV2V_UNCONNECTED_4270, SV2V_UNCONNECTED_4271, SV2V_UNCONNECTED_4272, SV2V_UNCONNECTED_4273, SV2V_UNCONNECTED_4274, SV2V_UNCONNECTED_4275, SV2V_UNCONNECTED_4276, SV2V_UNCONNECTED_4277, SV2V_UNCONNECTED_4278, SV2V_UNCONNECTED_4279, SV2V_UNCONNECTED_4280, SV2V_UNCONNECTED_4281, SV2V_UNCONNECTED_4282, SV2V_UNCONNECTED_4283, SV2V_UNCONNECTED_4284, SV2V_UNCONNECTED_4285, SV2V_UNCONNECTED_4286, SV2V_UNCONNECTED_4287, SV2V_UNCONNECTED_4288, SV2V_UNCONNECTED_4289, SV2V_UNCONNECTED_4290, SV2V_UNCONNECTED_4291, SV2V_UNCONNECTED_4292, SV2V_UNCONNECTED_4293, SV2V_UNCONNECTED_4294, SV2V_UNCONNECTED_4295, SV2V_UNCONNECTED_4296, SV2V_UNCONNECTED_4297, SV2V_UNCONNECTED_4298, SV2V_UNCONNECTED_4299, SV2V_UNCONNECTED_4300, SV2V_UNCONNECTED_4301, SV2V_UNCONNECTED_4302, SV2V_UNCONNECTED_4303, SV2V_UNCONNECTED_4304, SV2V_UNCONNECTED_4305, SV2V_UNCONNECTED_4306, SV2V_UNCONNECTED_4307, SV2V_UNCONNECTED_4308, SV2V_UNCONNECTED_4309, SV2V_UNCONNECTED_4310, SV2V_UNCONNECTED_4311, SV2V_UNCONNECTED_4312, SV2V_UNCONNECTED_4313, SV2V_UNCONNECTED_4314, SV2V_UNCONNECTED_4315, SV2V_UNCONNECTED_4316, SV2V_UNCONNECTED_4317, SV2V_UNCONNECTED_4318, SV2V_UNCONNECTED_4319, SV2V_UNCONNECTED_4320, SV2V_UNCONNECTED_4321, SV2V_UNCONNECTED_4322, SV2V_UNCONNECTED_4323, SV2V_UNCONNECTED_4324, SV2V_UNCONNECTED_4325, SV2V_UNCONNECTED_4326, SV2V_UNCONNECTED_4327, SV2V_UNCONNECTED_4328, SV2V_UNCONNECTED_4329, SV2V_UNCONNECTED_4330, SV2V_UNCONNECTED_4331, SV2V_UNCONNECTED_4332, SV2V_UNCONNECTED_4333, SV2V_UNCONNECTED_4334, SV2V_UNCONNECTED_4335, SV2V_UNCONNECTED_4336, SV2V_UNCONNECTED_4337, SV2V_UNCONNECTED_4338, SV2V_UNCONNECTED_4339, SV2V_UNCONNECTED_4340, SV2V_UNCONNECTED_4341, SV2V_UNCONNECTED_4342, SV2V_UNCONNECTED_4343, SV2V_UNCONNECTED_4344, SV2V_UNCONNECTED_4345, SV2V_UNCONNECTED_4346, SV2V_UNCONNECTED_4347, SV2V_UNCONNECTED_4348, SV2V_UNCONNECTED_4349, SV2V_UNCONNECTED_4350, SV2V_UNCONNECTED_4351, SV2V_UNCONNECTED_4352, SV2V_UNCONNECTED_4353, SV2V_UNCONNECTED_4354, SV2V_UNCONNECTED_4355, SV2V_UNCONNECTED_4356, SV2V_UNCONNECTED_4357, SV2V_UNCONNECTED_4358, SV2V_UNCONNECTED_4359, SV2V_UNCONNECTED_4360, SV2V_UNCONNECTED_4361, SV2V_UNCONNECTED_4362, SV2V_UNCONNECTED_4363, SV2V_UNCONNECTED_4364, SV2V_UNCONNECTED_4365, SV2V_UNCONNECTED_4366, SV2V_UNCONNECTED_4367, SV2V_UNCONNECTED_4368, SV2V_UNCONNECTED_4369, SV2V_UNCONNECTED_4370, SV2V_UNCONNECTED_4371, SV2V_UNCONNECTED_4372, SV2V_UNCONNECTED_4373, SV2V_UNCONNECTED_4374, SV2V_UNCONNECTED_4375, SV2V_UNCONNECTED_4376, SV2V_UNCONNECTED_4377, SV2V_UNCONNECTED_4378, SV2V_UNCONNECTED_4379, SV2V_UNCONNECTED_4380, SV2V_UNCONNECTED_4381, SV2V_UNCONNECTED_4382, SV2V_UNCONNECTED_4383, SV2V_UNCONNECTED_4384, SV2V_UNCONNECTED_4385, SV2V_UNCONNECTED_4386, SV2V_UNCONNECTED_4387, SV2V_UNCONNECTED_4388, SV2V_UNCONNECTED_4389, SV2V_UNCONNECTED_4390, SV2V_UNCONNECTED_4391, SV2V_UNCONNECTED_4392, SV2V_UNCONNECTED_4393, SV2V_UNCONNECTED_4394, SV2V_UNCONNECTED_4395, SV2V_UNCONNECTED_4396, SV2V_UNCONNECTED_4397, SV2V_UNCONNECTED_4398, SV2V_UNCONNECTED_4399, SV2V_UNCONNECTED_4400, SV2V_UNCONNECTED_4401, SV2V_UNCONNECTED_4402, SV2V_UNCONNECTED_4403, SV2V_UNCONNECTED_4404, SV2V_UNCONNECTED_4405, SV2V_UNCONNECTED_4406, SV2V_UNCONNECTED_4407, SV2V_UNCONNECTED_4408, SV2V_UNCONNECTED_4409, SV2V_UNCONNECTED_4410, SV2V_UNCONNECTED_4411, SV2V_UNCONNECTED_4412, SV2V_UNCONNECTED_4413, SV2V_UNCONNECTED_4414, SV2V_UNCONNECTED_4415, SV2V_UNCONNECTED_4416, SV2V_UNCONNECTED_4417, SV2V_UNCONNECTED_4418, SV2V_UNCONNECTED_4419, SV2V_UNCONNECTED_4420, SV2V_UNCONNECTED_4421, SV2V_UNCONNECTED_4422, SV2V_UNCONNECTED_4423, SV2V_UNCONNECTED_4424, SV2V_UNCONNECTED_4425, SV2V_UNCONNECTED_4426, SV2V_UNCONNECTED_4427, SV2V_UNCONNECTED_4428, SV2V_UNCONNECTED_4429, SV2V_UNCONNECTED_4430, SV2V_UNCONNECTED_4431, SV2V_UNCONNECTED_4432, SV2V_UNCONNECTED_4433, SV2V_UNCONNECTED_4434, SV2V_UNCONNECTED_4435, SV2V_UNCONNECTED_4436, SV2V_UNCONNECTED_4437, SV2V_UNCONNECTED_4438, SV2V_UNCONNECTED_4439, SV2V_UNCONNECTED_4440, SV2V_UNCONNECTED_4441, SV2V_UNCONNECTED_4442, SV2V_UNCONNECTED_4443, SV2V_UNCONNECTED_4444, SV2V_UNCONNECTED_4445, SV2V_UNCONNECTED_4446, SV2V_UNCONNECTED_4447, SV2V_UNCONNECTED_4448, SV2V_UNCONNECTED_4449, SV2V_UNCONNECTED_4450, SV2V_UNCONNECTED_4451, SV2V_UNCONNECTED_4452, SV2V_UNCONNECTED_4453, SV2V_UNCONNECTED_4454, SV2V_UNCONNECTED_4455, SV2V_UNCONNECTED_4456, SV2V_UNCONNECTED_4457, SV2V_UNCONNECTED_4458, SV2V_UNCONNECTED_4459, SV2V_UNCONNECTED_4460, SV2V_UNCONNECTED_4461, SV2V_UNCONNECTED_4462, SV2V_UNCONNECTED_4463, SV2V_UNCONNECTED_4464, SV2V_UNCONNECTED_4465, SV2V_UNCONNECTED_4466, SV2V_UNCONNECTED_4467, SV2V_UNCONNECTED_4468, SV2V_UNCONNECTED_4469, SV2V_UNCONNECTED_4470, SV2V_UNCONNECTED_4471, SV2V_UNCONNECTED_4472, SV2V_UNCONNECTED_4473, SV2V_UNCONNECTED_4474, SV2V_UNCONNECTED_4475, SV2V_UNCONNECTED_4476, SV2V_UNCONNECTED_4477, SV2V_UNCONNECTED_4478, SV2V_UNCONNECTED_4479, SV2V_UNCONNECTED_4480, SV2V_UNCONNECTED_4481, SV2V_UNCONNECTED_4482, SV2V_UNCONNECTED_4483, SV2V_UNCONNECTED_4484, SV2V_UNCONNECTED_4485, SV2V_UNCONNECTED_4486, SV2V_UNCONNECTED_4487, SV2V_UNCONNECTED_4488, SV2V_UNCONNECTED_4489, SV2V_UNCONNECTED_4490, SV2V_UNCONNECTED_4491, SV2V_UNCONNECTED_4492, SV2V_UNCONNECTED_4493, SV2V_UNCONNECTED_4494, SV2V_UNCONNECTED_4495, SV2V_UNCONNECTED_4496, SV2V_UNCONNECTED_4497, SV2V_UNCONNECTED_4498, SV2V_UNCONNECTED_4499, SV2V_UNCONNECTED_4500, SV2V_UNCONNECTED_4501, SV2V_UNCONNECTED_4502, SV2V_UNCONNECTED_4503, SV2V_UNCONNECTED_4504, SV2V_UNCONNECTED_4505, SV2V_UNCONNECTED_4506, SV2V_UNCONNECTED_4507, SV2V_UNCONNECTED_4508, SV2V_UNCONNECTED_4509, SV2V_UNCONNECTED_4510, SV2V_UNCONNECTED_4511, SV2V_UNCONNECTED_4512, SV2V_UNCONNECTED_4513, SV2V_UNCONNECTED_4514, SV2V_UNCONNECTED_4515, SV2V_UNCONNECTED_4516, SV2V_UNCONNECTED_4517, SV2V_UNCONNECTED_4518, SV2V_UNCONNECTED_4519, SV2V_UNCONNECTED_4520, SV2V_UNCONNECTED_4521, SV2V_UNCONNECTED_4522, SV2V_UNCONNECTED_4523, SV2V_UNCONNECTED_4524, SV2V_UNCONNECTED_4525, SV2V_UNCONNECTED_4526, SV2V_UNCONNECTED_4527, SV2V_UNCONNECTED_4528, SV2V_UNCONNECTED_4529, SV2V_UNCONNECTED_4530, SV2V_UNCONNECTED_4531, SV2V_UNCONNECTED_4532, SV2V_UNCONNECTED_4533, SV2V_UNCONNECTED_4534, SV2V_UNCONNECTED_4535, SV2V_UNCONNECTED_4536, SV2V_UNCONNECTED_4537, SV2V_UNCONNECTED_4538, SV2V_UNCONNECTED_4539, SV2V_UNCONNECTED_4540, SV2V_UNCONNECTED_4541, SV2V_UNCONNECTED_4542, SV2V_UNCONNECTED_4543, SV2V_UNCONNECTED_4544, SV2V_UNCONNECTED_4545, SV2V_UNCONNECTED_4546, SV2V_UNCONNECTED_4547, SV2V_UNCONNECTED_4548, SV2V_UNCONNECTED_4549, SV2V_UNCONNECTED_4550, SV2V_UNCONNECTED_4551, SV2V_UNCONNECTED_4552, SV2V_UNCONNECTED_4553, SV2V_UNCONNECTED_4554, SV2V_UNCONNECTED_4555, SV2V_UNCONNECTED_4556, SV2V_UNCONNECTED_4557, SV2V_UNCONNECTED_4558, SV2V_UNCONNECTED_4559, SV2V_UNCONNECTED_4560, SV2V_UNCONNECTED_4561, SV2V_UNCONNECTED_4562, SV2V_UNCONNECTED_4563, SV2V_UNCONNECTED_4564, SV2V_UNCONNECTED_4565, SV2V_UNCONNECTED_4566, SV2V_UNCONNECTED_4567, SV2V_UNCONNECTED_4568, SV2V_UNCONNECTED_4569, SV2V_UNCONNECTED_4570, SV2V_UNCONNECTED_4571, SV2V_UNCONNECTED_4572, SV2V_UNCONNECTED_4573, SV2V_UNCONNECTED_4574, SV2V_UNCONNECTED_4575, SV2V_UNCONNECTED_4576, SV2V_UNCONNECTED_4577, SV2V_UNCONNECTED_4578, SV2V_UNCONNECTED_4579, SV2V_UNCONNECTED_4580, SV2V_UNCONNECTED_4581, SV2V_UNCONNECTED_4582, SV2V_UNCONNECTED_4583, SV2V_UNCONNECTED_4584, SV2V_UNCONNECTED_4585, SV2V_UNCONNECTED_4586, SV2V_UNCONNECTED_4587, SV2V_UNCONNECTED_4588, SV2V_UNCONNECTED_4589, SV2V_UNCONNECTED_4590, SV2V_UNCONNECTED_4591, SV2V_UNCONNECTED_4592, SV2V_UNCONNECTED_4593, SV2V_UNCONNECTED_4594, SV2V_UNCONNECTED_4595, SV2V_UNCONNECTED_4596, SV2V_UNCONNECTED_4597, SV2V_UNCONNECTED_4598, SV2V_UNCONNECTED_4599, SV2V_UNCONNECTED_4600, SV2V_UNCONNECTED_4601, SV2V_UNCONNECTED_4602, SV2V_UNCONNECTED_4603, SV2V_UNCONNECTED_4604, SV2V_UNCONNECTED_4605, SV2V_UNCONNECTED_4606, SV2V_UNCONNECTED_4607, SV2V_UNCONNECTED_4608, SV2V_UNCONNECTED_4609, SV2V_UNCONNECTED_4610, SV2V_UNCONNECTED_4611, SV2V_UNCONNECTED_4612, SV2V_UNCONNECTED_4613, SV2V_UNCONNECTED_4614, SV2V_UNCONNECTED_4615, SV2V_UNCONNECTED_4616, SV2V_UNCONNECTED_4617, SV2V_UNCONNECTED_4618, SV2V_UNCONNECTED_4619, SV2V_UNCONNECTED_4620, SV2V_UNCONNECTED_4621, SV2V_UNCONNECTED_4622, SV2V_UNCONNECTED_4623, SV2V_UNCONNECTED_4624, SV2V_UNCONNECTED_4625, SV2V_UNCONNECTED_4626, SV2V_UNCONNECTED_4627, SV2V_UNCONNECTED_4628, SV2V_UNCONNECTED_4629, SV2V_UNCONNECTED_4630, SV2V_UNCONNECTED_4631, SV2V_UNCONNECTED_4632, SV2V_UNCONNECTED_4633, SV2V_UNCONNECTED_4634, SV2V_UNCONNECTED_4635, SV2V_UNCONNECTED_4636, SV2V_UNCONNECTED_4637, SV2V_UNCONNECTED_4638, SV2V_UNCONNECTED_4639, SV2V_UNCONNECTED_4640, SV2V_UNCONNECTED_4641, SV2V_UNCONNECTED_4642, SV2V_UNCONNECTED_4643, SV2V_UNCONNECTED_4644, SV2V_UNCONNECTED_4645, SV2V_UNCONNECTED_4646, SV2V_UNCONNECTED_4647, SV2V_UNCONNECTED_4648, SV2V_UNCONNECTED_4649, SV2V_UNCONNECTED_4650, SV2V_UNCONNECTED_4651, SV2V_UNCONNECTED_4652, SV2V_UNCONNECTED_4653, SV2V_UNCONNECTED_4654, SV2V_UNCONNECTED_4655, SV2V_UNCONNECTED_4656, SV2V_UNCONNECTED_4657, SV2V_UNCONNECTED_4658, SV2V_UNCONNECTED_4659, SV2V_UNCONNECTED_4660, SV2V_UNCONNECTED_4661, SV2V_UNCONNECTED_4662, SV2V_UNCONNECTED_4663, SV2V_UNCONNECTED_4664, SV2V_UNCONNECTED_4665, SV2V_UNCONNECTED_4666, SV2V_UNCONNECTED_4667, SV2V_UNCONNECTED_4668, SV2V_UNCONNECTED_4669, SV2V_UNCONNECTED_4670, SV2V_UNCONNECTED_4671, SV2V_UNCONNECTED_4672, SV2V_UNCONNECTED_4673, SV2V_UNCONNECTED_4674, SV2V_UNCONNECTED_4675, SV2V_UNCONNECTED_4676, SV2V_UNCONNECTED_4677, SV2V_UNCONNECTED_4678, SV2V_UNCONNECTED_4679, SV2V_UNCONNECTED_4680, SV2V_UNCONNECTED_4681, SV2V_UNCONNECTED_4682, SV2V_UNCONNECTED_4683, SV2V_UNCONNECTED_4684, SV2V_UNCONNECTED_4685, SV2V_UNCONNECTED_4686, SV2V_UNCONNECTED_4687, SV2V_UNCONNECTED_4688, SV2V_UNCONNECTED_4689, SV2V_UNCONNECTED_4690, SV2V_UNCONNECTED_4691, SV2V_UNCONNECTED_4692, SV2V_UNCONNECTED_4693, SV2V_UNCONNECTED_4694, SV2V_UNCONNECTED_4695, SV2V_UNCONNECTED_4696, SV2V_UNCONNECTED_4697, SV2V_UNCONNECTED_4698, SV2V_UNCONNECTED_4699, SV2V_UNCONNECTED_4700, SV2V_UNCONNECTED_4701, SV2V_UNCONNECTED_4702, SV2V_UNCONNECTED_4703, SV2V_UNCONNECTED_4704, SV2V_UNCONNECTED_4705, SV2V_UNCONNECTED_4706, SV2V_UNCONNECTED_4707, SV2V_UNCONNECTED_4708, SV2V_UNCONNECTED_4709, SV2V_UNCONNECTED_4710, SV2V_UNCONNECTED_4711, SV2V_UNCONNECTED_4712, SV2V_UNCONNECTED_4713, SV2V_UNCONNECTED_4714, SV2V_UNCONNECTED_4715, SV2V_UNCONNECTED_4716, SV2V_UNCONNECTED_4717, SV2V_UNCONNECTED_4718, SV2V_UNCONNECTED_4719, SV2V_UNCONNECTED_4720, SV2V_UNCONNECTED_4721, SV2V_UNCONNECTED_4722, SV2V_UNCONNECTED_4723, SV2V_UNCONNECTED_4724, SV2V_UNCONNECTED_4725, SV2V_UNCONNECTED_4726, SV2V_UNCONNECTED_4727, SV2V_UNCONNECTED_4728, SV2V_UNCONNECTED_4729, SV2V_UNCONNECTED_4730, SV2V_UNCONNECTED_4731, SV2V_UNCONNECTED_4732, SV2V_UNCONNECTED_4733, SV2V_UNCONNECTED_4734, SV2V_UNCONNECTED_4735, SV2V_UNCONNECTED_4736, SV2V_UNCONNECTED_4737, SV2V_UNCONNECTED_4738, SV2V_UNCONNECTED_4739, SV2V_UNCONNECTED_4740, SV2V_UNCONNECTED_4741, SV2V_UNCONNECTED_4742, SV2V_UNCONNECTED_4743, SV2V_UNCONNECTED_4744, SV2V_UNCONNECTED_4745, SV2V_UNCONNECTED_4746, SV2V_UNCONNECTED_4747, SV2V_UNCONNECTED_4748, SV2V_UNCONNECTED_4749, SV2V_UNCONNECTED_4750, SV2V_UNCONNECTED_4751, SV2V_UNCONNECTED_4752, SV2V_UNCONNECTED_4753, SV2V_UNCONNECTED_4754, SV2V_UNCONNECTED_4755, SV2V_UNCONNECTED_4756, SV2V_UNCONNECTED_4757, SV2V_UNCONNECTED_4758, SV2V_UNCONNECTED_4759, SV2V_UNCONNECTED_4760, SV2V_UNCONNECTED_4761, SV2V_UNCONNECTED_4762, SV2V_UNCONNECTED_4763, SV2V_UNCONNECTED_4764, SV2V_UNCONNECTED_4765, SV2V_UNCONNECTED_4766, SV2V_UNCONNECTED_4767, SV2V_UNCONNECTED_4768, SV2V_UNCONNECTED_4769, SV2V_UNCONNECTED_4770, SV2V_UNCONNECTED_4771, SV2V_UNCONNECTED_4772, SV2V_UNCONNECTED_4773, SV2V_UNCONNECTED_4774, SV2V_UNCONNECTED_4775, SV2V_UNCONNECTED_4776, SV2V_UNCONNECTED_4777, SV2V_UNCONNECTED_4778, SV2V_UNCONNECTED_4779, SV2V_UNCONNECTED_4780, SV2V_UNCONNECTED_4781, SV2V_UNCONNECTED_4782, SV2V_UNCONNECTED_4783, SV2V_UNCONNECTED_4784, SV2V_UNCONNECTED_4785, SV2V_UNCONNECTED_4786, SV2V_UNCONNECTED_4787, SV2V_UNCONNECTED_4788, SV2V_UNCONNECTED_4789, SV2V_UNCONNECTED_4790, SV2V_UNCONNECTED_4791, SV2V_UNCONNECTED_4792, SV2V_UNCONNECTED_4793, SV2V_UNCONNECTED_4794, SV2V_UNCONNECTED_4795, SV2V_UNCONNECTED_4796, SV2V_UNCONNECTED_4797, SV2V_UNCONNECTED_4798, SV2V_UNCONNECTED_4799, SV2V_UNCONNECTED_4800, SV2V_UNCONNECTED_4801, SV2V_UNCONNECTED_4802, SV2V_UNCONNECTED_4803, SV2V_UNCONNECTED_4804, SV2V_UNCONNECTED_4805, SV2V_UNCONNECTED_4806, SV2V_UNCONNECTED_4807, SV2V_UNCONNECTED_4808, SV2V_UNCONNECTED_4809, SV2V_UNCONNECTED_4810, SV2V_UNCONNECTED_4811, SV2V_UNCONNECTED_4812, SV2V_UNCONNECTED_4813, SV2V_UNCONNECTED_4814, SV2V_UNCONNECTED_4815, SV2V_UNCONNECTED_4816, SV2V_UNCONNECTED_4817, SV2V_UNCONNECTED_4818, SV2V_UNCONNECTED_4819, SV2V_UNCONNECTED_4820, SV2V_UNCONNECTED_4821, SV2V_UNCONNECTED_4822, SV2V_UNCONNECTED_4823, SV2V_UNCONNECTED_4824, SV2V_UNCONNECTED_4825, SV2V_UNCONNECTED_4826, SV2V_UNCONNECTED_4827, SV2V_UNCONNECTED_4828, SV2V_UNCONNECTED_4829, SV2V_UNCONNECTED_4830, SV2V_UNCONNECTED_4831, SV2V_UNCONNECTED_4832, SV2V_UNCONNECTED_4833, SV2V_UNCONNECTED_4834, SV2V_UNCONNECTED_4835, SV2V_UNCONNECTED_4836, SV2V_UNCONNECTED_4837, SV2V_UNCONNECTED_4838, SV2V_UNCONNECTED_4839, SV2V_UNCONNECTED_4840, SV2V_UNCONNECTED_4841, SV2V_UNCONNECTED_4842, SV2V_UNCONNECTED_4843, SV2V_UNCONNECTED_4844, SV2V_UNCONNECTED_4845, SV2V_UNCONNECTED_4846, SV2V_UNCONNECTED_4847, SV2V_UNCONNECTED_4848, SV2V_UNCONNECTED_4849, SV2V_UNCONNECTED_4850, SV2V_UNCONNECTED_4851, SV2V_UNCONNECTED_4852, SV2V_UNCONNECTED_4853, SV2V_UNCONNECTED_4854, SV2V_UNCONNECTED_4855, SV2V_UNCONNECTED_4856, SV2V_UNCONNECTED_4857, SV2V_UNCONNECTED_4858, SV2V_UNCONNECTED_4859, SV2V_UNCONNECTED_4860, SV2V_UNCONNECTED_4861, SV2V_UNCONNECTED_4862, SV2V_UNCONNECTED_4863, SV2V_UNCONNECTED_4864, SV2V_UNCONNECTED_4865, SV2V_UNCONNECTED_4866, SV2V_UNCONNECTED_4867, SV2V_UNCONNECTED_4868, SV2V_UNCONNECTED_4869, SV2V_UNCONNECTED_4870, SV2V_UNCONNECTED_4871, SV2V_UNCONNECTED_4872, SV2V_UNCONNECTED_4873, SV2V_UNCONNECTED_4874, SV2V_UNCONNECTED_4875, SV2V_UNCONNECTED_4876, SV2V_UNCONNECTED_4877, SV2V_UNCONNECTED_4878, SV2V_UNCONNECTED_4879, SV2V_UNCONNECTED_4880, SV2V_UNCONNECTED_4881, SV2V_UNCONNECTED_4882, SV2V_UNCONNECTED_4883, SV2V_UNCONNECTED_4884, SV2V_UNCONNECTED_4885, SV2V_UNCONNECTED_4886, SV2V_UNCONNECTED_4887, SV2V_UNCONNECTED_4888, SV2V_UNCONNECTED_4889, SV2V_UNCONNECTED_4890, SV2V_UNCONNECTED_4891, SV2V_UNCONNECTED_4892, SV2V_UNCONNECTED_4893, SV2V_UNCONNECTED_4894, SV2V_UNCONNECTED_4895, SV2V_UNCONNECTED_4896, SV2V_UNCONNECTED_4897, SV2V_UNCONNECTED_4898, SV2V_UNCONNECTED_4899, SV2V_UNCONNECTED_4900, SV2V_UNCONNECTED_4901, SV2V_UNCONNECTED_4902, SV2V_UNCONNECTED_4903, SV2V_UNCONNECTED_4904, SV2V_UNCONNECTED_4905, SV2V_UNCONNECTED_4906, SV2V_UNCONNECTED_4907, SV2V_UNCONNECTED_4908, SV2V_UNCONNECTED_4909, SV2V_UNCONNECTED_4910, SV2V_UNCONNECTED_4911, SV2V_UNCONNECTED_4912, SV2V_UNCONNECTED_4913, SV2V_UNCONNECTED_4914, SV2V_UNCONNECTED_4915, SV2V_UNCONNECTED_4916, SV2V_UNCONNECTED_4917, SV2V_UNCONNECTED_4918, SV2V_UNCONNECTED_4919, SV2V_UNCONNECTED_4920, SV2V_UNCONNECTED_4921, SV2V_UNCONNECTED_4922, SV2V_UNCONNECTED_4923, SV2V_UNCONNECTED_4924, SV2V_UNCONNECTED_4925, SV2V_UNCONNECTED_4926, SV2V_UNCONNECTED_4927, SV2V_UNCONNECTED_4928, SV2V_UNCONNECTED_4929, SV2V_UNCONNECTED_4930, SV2V_UNCONNECTED_4931, SV2V_UNCONNECTED_4932, SV2V_UNCONNECTED_4933, SV2V_UNCONNECTED_4934, SV2V_UNCONNECTED_4935, SV2V_UNCONNECTED_4936, SV2V_UNCONNECTED_4937, SV2V_UNCONNECTED_4938, SV2V_UNCONNECTED_4939, SV2V_UNCONNECTED_4940, SV2V_UNCONNECTED_4941, SV2V_UNCONNECTED_4942, SV2V_UNCONNECTED_4943, SV2V_UNCONNECTED_4944, SV2V_UNCONNECTED_4945, SV2V_UNCONNECTED_4946, SV2V_UNCONNECTED_4947, SV2V_UNCONNECTED_4948, SV2V_UNCONNECTED_4949, SV2V_UNCONNECTED_4950, SV2V_UNCONNECTED_4951, SV2V_UNCONNECTED_4952, SV2V_UNCONNECTED_4953, SV2V_UNCONNECTED_4954, SV2V_UNCONNECTED_4955, SV2V_UNCONNECTED_4956, SV2V_UNCONNECTED_4957, SV2V_UNCONNECTED_4958, SV2V_UNCONNECTED_4959, SV2V_UNCONNECTED_4960, SV2V_UNCONNECTED_4961, SV2V_UNCONNECTED_4962, SV2V_UNCONNECTED_4963, SV2V_UNCONNECTED_4964, SV2V_UNCONNECTED_4965, SV2V_UNCONNECTED_4966, SV2V_UNCONNECTED_4967, SV2V_UNCONNECTED_4968, SV2V_UNCONNECTED_4969, SV2V_UNCONNECTED_4970, SV2V_UNCONNECTED_4971, SV2V_UNCONNECTED_4972, SV2V_UNCONNECTED_4973, SV2V_UNCONNECTED_4974, SV2V_UNCONNECTED_4975, SV2V_UNCONNECTED_4976, SV2V_UNCONNECTED_4977, SV2V_UNCONNECTED_4978, SV2V_UNCONNECTED_4979, SV2V_UNCONNECTED_4980, SV2V_UNCONNECTED_4981, SV2V_UNCONNECTED_4982, SV2V_UNCONNECTED_4983, SV2V_UNCONNECTED_4984, SV2V_UNCONNECTED_4985, SV2V_UNCONNECTED_4986, SV2V_UNCONNECTED_4987, SV2V_UNCONNECTED_4988, SV2V_UNCONNECTED_4989, SV2V_UNCONNECTED_4990, SV2V_UNCONNECTED_4991, SV2V_UNCONNECTED_4992, SV2V_UNCONNECTED_4993, SV2V_UNCONNECTED_4994, SV2V_UNCONNECTED_4995, SV2V_UNCONNECTED_4996, SV2V_UNCONNECTED_4997, SV2V_UNCONNECTED_4998, SV2V_UNCONNECTED_4999, SV2V_UNCONNECTED_5000, SV2V_UNCONNECTED_5001, SV2V_UNCONNECTED_5002, SV2V_UNCONNECTED_5003, SV2V_UNCONNECTED_5004, SV2V_UNCONNECTED_5005, SV2V_UNCONNECTED_5006, SV2V_UNCONNECTED_5007, SV2V_UNCONNECTED_5008, SV2V_UNCONNECTED_5009, SV2V_UNCONNECTED_5010, SV2V_UNCONNECTED_5011, SV2V_UNCONNECTED_5012, SV2V_UNCONNECTED_5013, SV2V_UNCONNECTED_5014, SV2V_UNCONNECTED_5015, SV2V_UNCONNECTED_5016, SV2V_UNCONNECTED_5017, SV2V_UNCONNECTED_5018, SV2V_UNCONNECTED_5019, SV2V_UNCONNECTED_5020, SV2V_UNCONNECTED_5021, SV2V_UNCONNECTED_5022, SV2V_UNCONNECTED_5023, SV2V_UNCONNECTED_5024, SV2V_UNCONNECTED_5025, SV2V_UNCONNECTED_5026, SV2V_UNCONNECTED_5027, SV2V_UNCONNECTED_5028, SV2V_UNCONNECTED_5029, SV2V_UNCONNECTED_5030, SV2V_UNCONNECTED_5031, SV2V_UNCONNECTED_5032, SV2V_UNCONNECTED_5033, SV2V_UNCONNECTED_5034, SV2V_UNCONNECTED_5035, SV2V_UNCONNECTED_5036, SV2V_UNCONNECTED_5037, SV2V_UNCONNECTED_5038, SV2V_UNCONNECTED_5039, SV2V_UNCONNECTED_5040, SV2V_UNCONNECTED_5041, SV2V_UNCONNECTED_5042, SV2V_UNCONNECTED_5043, SV2V_UNCONNECTED_5044, SV2V_UNCONNECTED_5045, SV2V_UNCONNECTED_5046, SV2V_UNCONNECTED_5047, SV2V_UNCONNECTED_5048, SV2V_UNCONNECTED_5049, SV2V_UNCONNECTED_5050, SV2V_UNCONNECTED_5051, SV2V_UNCONNECTED_5052, SV2V_UNCONNECTED_5053, SV2V_UNCONNECTED_5054, SV2V_UNCONNECTED_5055, SV2V_UNCONNECTED_5056, SV2V_UNCONNECTED_5057, SV2V_UNCONNECTED_5058, SV2V_UNCONNECTED_5059, SV2V_UNCONNECTED_5060, SV2V_UNCONNECTED_5061, SV2V_UNCONNECTED_5062, SV2V_UNCONNECTED_5063, SV2V_UNCONNECTED_5064, SV2V_UNCONNECTED_5065, SV2V_UNCONNECTED_5066, SV2V_UNCONNECTED_5067, SV2V_UNCONNECTED_5068, SV2V_UNCONNECTED_5069, SV2V_UNCONNECTED_5070, SV2V_UNCONNECTED_5071, SV2V_UNCONNECTED_5072, SV2V_UNCONNECTED_5073, SV2V_UNCONNECTED_5074, SV2V_UNCONNECTED_5075, SV2V_UNCONNECTED_5076, SV2V_UNCONNECTED_5077, SV2V_UNCONNECTED_5078, SV2V_UNCONNECTED_5079, SV2V_UNCONNECTED_5080, SV2V_UNCONNECTED_5081, SV2V_UNCONNECTED_5082, SV2V_UNCONNECTED_5083, SV2V_UNCONNECTED_5084, SV2V_UNCONNECTED_5085, SV2V_UNCONNECTED_5086, SV2V_UNCONNECTED_5087, SV2V_UNCONNECTED_5088, SV2V_UNCONNECTED_5089, SV2V_UNCONNECTED_5090, SV2V_UNCONNECTED_5091, SV2V_UNCONNECTED_5092, SV2V_UNCONNECTED_5093, SV2V_UNCONNECTED_5094, SV2V_UNCONNECTED_5095, SV2V_UNCONNECTED_5096, SV2V_UNCONNECTED_5097, SV2V_UNCONNECTED_5098, SV2V_UNCONNECTED_5099, SV2V_UNCONNECTED_5100, SV2V_UNCONNECTED_5101, SV2V_UNCONNECTED_5102, SV2V_UNCONNECTED_5103, SV2V_UNCONNECTED_5104, SV2V_UNCONNECTED_5105, SV2V_UNCONNECTED_5106, SV2V_UNCONNECTED_5107, SV2V_UNCONNECTED_5108, SV2V_UNCONNECTED_5109, SV2V_UNCONNECTED_5110, SV2V_UNCONNECTED_5111, SV2V_UNCONNECTED_5112, SV2V_UNCONNECTED_5113, SV2V_UNCONNECTED_5114, SV2V_UNCONNECTED_5115, SV2V_UNCONNECTED_5116, SV2V_UNCONNECTED_5117, SV2V_UNCONNECTED_5118, SV2V_UNCONNECTED_5119, SV2V_UNCONNECTED_5120, SV2V_UNCONNECTED_5121, SV2V_UNCONNECTED_5122, SV2V_UNCONNECTED_5123, SV2V_UNCONNECTED_5124, SV2V_UNCONNECTED_5125, SV2V_UNCONNECTED_5126, SV2V_UNCONNECTED_5127, SV2V_UNCONNECTED_5128, SV2V_UNCONNECTED_5129, SV2V_UNCONNECTED_5130, SV2V_UNCONNECTED_5131, SV2V_UNCONNECTED_5132, SV2V_UNCONNECTED_5133, SV2V_UNCONNECTED_5134, SV2V_UNCONNECTED_5135, SV2V_UNCONNECTED_5136, SV2V_UNCONNECTED_5137, SV2V_UNCONNECTED_5138, SV2V_UNCONNECTED_5139, SV2V_UNCONNECTED_5140, SV2V_UNCONNECTED_5141, SV2V_UNCONNECTED_5142, SV2V_UNCONNECTED_5143, SV2V_UNCONNECTED_5144, SV2V_UNCONNECTED_5145, SV2V_UNCONNECTED_5146, SV2V_UNCONNECTED_5147, SV2V_UNCONNECTED_5148, SV2V_UNCONNECTED_5149, SV2V_UNCONNECTED_5150, SV2V_UNCONNECTED_5151, SV2V_UNCONNECTED_5152, SV2V_UNCONNECTED_5153, SV2V_UNCONNECTED_5154, SV2V_UNCONNECTED_5155, SV2V_UNCONNECTED_5156, SV2V_UNCONNECTED_5157, SV2V_UNCONNECTED_5158, SV2V_UNCONNECTED_5159, SV2V_UNCONNECTED_5160, SV2V_UNCONNECTED_5161, SV2V_UNCONNECTED_5162, SV2V_UNCONNECTED_5163, SV2V_UNCONNECTED_5164, SV2V_UNCONNECTED_5165, SV2V_UNCONNECTED_5166, SV2V_UNCONNECTED_5167, SV2V_UNCONNECTED_5168, SV2V_UNCONNECTED_5169, SV2V_UNCONNECTED_5170, SV2V_UNCONNECTED_5171, SV2V_UNCONNECTED_5172, SV2V_UNCONNECTED_5173, SV2V_UNCONNECTED_5174, SV2V_UNCONNECTED_5175, SV2V_UNCONNECTED_5176, SV2V_UNCONNECTED_5177, SV2V_UNCONNECTED_5178, SV2V_UNCONNECTED_5179, SV2V_UNCONNECTED_5180, SV2V_UNCONNECTED_5181, SV2V_UNCONNECTED_5182, SV2V_UNCONNECTED_5183, SV2V_UNCONNECTED_5184, SV2V_UNCONNECTED_5185, SV2V_UNCONNECTED_5186, SV2V_UNCONNECTED_5187, SV2V_UNCONNECTED_5188, SV2V_UNCONNECTED_5189, SV2V_UNCONNECTED_5190, SV2V_UNCONNECTED_5191, SV2V_UNCONNECTED_5192, SV2V_UNCONNECTED_5193, SV2V_UNCONNECTED_5194, SV2V_UNCONNECTED_5195, SV2V_UNCONNECTED_5196, SV2V_UNCONNECTED_5197, SV2V_UNCONNECTED_5198, SV2V_UNCONNECTED_5199, SV2V_UNCONNECTED_5200, SV2V_UNCONNECTED_5201, SV2V_UNCONNECTED_5202, SV2V_UNCONNECTED_5203, SV2V_UNCONNECTED_5204, SV2V_UNCONNECTED_5205, SV2V_UNCONNECTED_5206, SV2V_UNCONNECTED_5207, SV2V_UNCONNECTED_5208, SV2V_UNCONNECTED_5209, SV2V_UNCONNECTED_5210, SV2V_UNCONNECTED_5211, SV2V_UNCONNECTED_5212, SV2V_UNCONNECTED_5213, SV2V_UNCONNECTED_5214, SV2V_UNCONNECTED_5215, SV2V_UNCONNECTED_5216, SV2V_UNCONNECTED_5217, SV2V_UNCONNECTED_5218, SV2V_UNCONNECTED_5219, SV2V_UNCONNECTED_5220, SV2V_UNCONNECTED_5221, SV2V_UNCONNECTED_5222, SV2V_UNCONNECTED_5223, SV2V_UNCONNECTED_5224, SV2V_UNCONNECTED_5225, SV2V_UNCONNECTED_5226, SV2V_UNCONNECTED_5227, SV2V_UNCONNECTED_5228, SV2V_UNCONNECTED_5229, SV2V_UNCONNECTED_5230, SV2V_UNCONNECTED_5231, SV2V_UNCONNECTED_5232, SV2V_UNCONNECTED_5233, SV2V_UNCONNECTED_5234, SV2V_UNCONNECTED_5235, SV2V_UNCONNECTED_5236, SV2V_UNCONNECTED_5237, SV2V_UNCONNECTED_5238, SV2V_UNCONNECTED_5239, SV2V_UNCONNECTED_5240, SV2V_UNCONNECTED_5241, SV2V_UNCONNECTED_5242, SV2V_UNCONNECTED_5243, SV2V_UNCONNECTED_5244, SV2V_UNCONNECTED_5245, SV2V_UNCONNECTED_5246, SV2V_UNCONNECTED_5247, SV2V_UNCONNECTED_5248, SV2V_UNCONNECTED_5249, SV2V_UNCONNECTED_5250, SV2V_UNCONNECTED_5251, SV2V_UNCONNECTED_5252, SV2V_UNCONNECTED_5253, SV2V_UNCONNECTED_5254, SV2V_UNCONNECTED_5255, SV2V_UNCONNECTED_5256, SV2V_UNCONNECTED_5257, SV2V_UNCONNECTED_5258, SV2V_UNCONNECTED_5259, SV2V_UNCONNECTED_5260, SV2V_UNCONNECTED_5261, SV2V_UNCONNECTED_5262, SV2V_UNCONNECTED_5263, SV2V_UNCONNECTED_5264, SV2V_UNCONNECTED_5265, SV2V_UNCONNECTED_5266, SV2V_UNCONNECTED_5267, SV2V_UNCONNECTED_5268, SV2V_UNCONNECTED_5269, SV2V_UNCONNECTED_5270, SV2V_UNCONNECTED_5271, SV2V_UNCONNECTED_5272, SV2V_UNCONNECTED_5273, SV2V_UNCONNECTED_5274, SV2V_UNCONNECTED_5275, SV2V_UNCONNECTED_5276, SV2V_UNCONNECTED_5277, SV2V_UNCONNECTED_5278, SV2V_UNCONNECTED_5279, SV2V_UNCONNECTED_5280, SV2V_UNCONNECTED_5281, SV2V_UNCONNECTED_5282, SV2V_UNCONNECTED_5283, SV2V_UNCONNECTED_5284, SV2V_UNCONNECTED_5285, SV2V_UNCONNECTED_5286, SV2V_UNCONNECTED_5287, SV2V_UNCONNECTED_5288, SV2V_UNCONNECTED_5289, SV2V_UNCONNECTED_5290, SV2V_UNCONNECTED_5291, SV2V_UNCONNECTED_5292, SV2V_UNCONNECTED_5293, SV2V_UNCONNECTED_5294, SV2V_UNCONNECTED_5295, SV2V_UNCONNECTED_5296, SV2V_UNCONNECTED_5297, SV2V_UNCONNECTED_5298, SV2V_UNCONNECTED_5299, SV2V_UNCONNECTED_5300, SV2V_UNCONNECTED_5301, SV2V_UNCONNECTED_5302, SV2V_UNCONNECTED_5303, SV2V_UNCONNECTED_5304, SV2V_UNCONNECTED_5305, SV2V_UNCONNECTED_5306, SV2V_UNCONNECTED_5307, SV2V_UNCONNECTED_5308, SV2V_UNCONNECTED_5309, SV2V_UNCONNECTED_5310, SV2V_UNCONNECTED_5311, SV2V_UNCONNECTED_5312, SV2V_UNCONNECTED_5313, SV2V_UNCONNECTED_5314, SV2V_UNCONNECTED_5315, SV2V_UNCONNECTED_5316, SV2V_UNCONNECTED_5317, SV2V_UNCONNECTED_5318, SV2V_UNCONNECTED_5319, SV2V_UNCONNECTED_5320, SV2V_UNCONNECTED_5321, SV2V_UNCONNECTED_5322, SV2V_UNCONNECTED_5323, SV2V_UNCONNECTED_5324, SV2V_UNCONNECTED_5325, SV2V_UNCONNECTED_5326, SV2V_UNCONNECTED_5327, SV2V_UNCONNECTED_5328, SV2V_UNCONNECTED_5329, SV2V_UNCONNECTED_5330, SV2V_UNCONNECTED_5331, SV2V_UNCONNECTED_5332, SV2V_UNCONNECTED_5333, SV2V_UNCONNECTED_5334, SV2V_UNCONNECTED_5335, SV2V_UNCONNECTED_5336, SV2V_UNCONNECTED_5337, SV2V_UNCONNECTED_5338, SV2V_UNCONNECTED_5339, SV2V_UNCONNECTED_5340, SV2V_UNCONNECTED_5341, SV2V_UNCONNECTED_5342, SV2V_UNCONNECTED_5343, SV2V_UNCONNECTED_5344, SV2V_UNCONNECTED_5345, SV2V_UNCONNECTED_5346, SV2V_UNCONNECTED_5347, SV2V_UNCONNECTED_5348, SV2V_UNCONNECTED_5349, SV2V_UNCONNECTED_5350, SV2V_UNCONNECTED_5351, SV2V_UNCONNECTED_5352, SV2V_UNCONNECTED_5353, SV2V_UNCONNECTED_5354, SV2V_UNCONNECTED_5355, SV2V_UNCONNECTED_5356, SV2V_UNCONNECTED_5357, SV2V_UNCONNECTED_5358, SV2V_UNCONNECTED_5359, SV2V_UNCONNECTED_5360, SV2V_UNCONNECTED_5361, SV2V_UNCONNECTED_5362, SV2V_UNCONNECTED_5363, SV2V_UNCONNECTED_5364, SV2V_UNCONNECTED_5365, SV2V_UNCONNECTED_5366, SV2V_UNCONNECTED_5367, SV2V_UNCONNECTED_5368, SV2V_UNCONNECTED_5369, SV2V_UNCONNECTED_5370, SV2V_UNCONNECTED_5371, SV2V_UNCONNECTED_5372, SV2V_UNCONNECTED_5373, SV2V_UNCONNECTED_5374, SV2V_UNCONNECTED_5375, SV2V_UNCONNECTED_5376, SV2V_UNCONNECTED_5377, SV2V_UNCONNECTED_5378, SV2V_UNCONNECTED_5379, SV2V_UNCONNECTED_5380, SV2V_UNCONNECTED_5381, SV2V_UNCONNECTED_5382, SV2V_UNCONNECTED_5383, SV2V_UNCONNECTED_5384, SV2V_UNCONNECTED_5385, SV2V_UNCONNECTED_5386, SV2V_UNCONNECTED_5387, SV2V_UNCONNECTED_5388, SV2V_UNCONNECTED_5389, SV2V_UNCONNECTED_5390, SV2V_UNCONNECTED_5391, SV2V_UNCONNECTED_5392, SV2V_UNCONNECTED_5393, SV2V_UNCONNECTED_5394, SV2V_UNCONNECTED_5395, SV2V_UNCONNECTED_5396, SV2V_UNCONNECTED_5397, SV2V_UNCONNECTED_5398, SV2V_UNCONNECTED_5399, SV2V_UNCONNECTED_5400, SV2V_UNCONNECTED_5401, SV2V_UNCONNECTED_5402, SV2V_UNCONNECTED_5403, SV2V_UNCONNECTED_5404, SV2V_UNCONNECTED_5405, SV2V_UNCONNECTED_5406, SV2V_UNCONNECTED_5407, SV2V_UNCONNECTED_5408, SV2V_UNCONNECTED_5409, SV2V_UNCONNECTED_5410, SV2V_UNCONNECTED_5411, SV2V_UNCONNECTED_5412, SV2V_UNCONNECTED_5413, SV2V_UNCONNECTED_5414, SV2V_UNCONNECTED_5415, SV2V_UNCONNECTED_5416, SV2V_UNCONNECTED_5417, SV2V_UNCONNECTED_5418, SV2V_UNCONNECTED_5419, SV2V_UNCONNECTED_5420, SV2V_UNCONNECTED_5421, SV2V_UNCONNECTED_5422, SV2V_UNCONNECTED_5423, SV2V_UNCONNECTED_5424, SV2V_UNCONNECTED_5425, SV2V_UNCONNECTED_5426, SV2V_UNCONNECTED_5427, SV2V_UNCONNECTED_5428, SV2V_UNCONNECTED_5429, SV2V_UNCONNECTED_5430, SV2V_UNCONNECTED_5431, SV2V_UNCONNECTED_5432, SV2V_UNCONNECTED_5433, SV2V_UNCONNECTED_5434, SV2V_UNCONNECTED_5435, SV2V_UNCONNECTED_5436, SV2V_UNCONNECTED_5437, SV2V_UNCONNECTED_5438, SV2V_UNCONNECTED_5439, SV2V_UNCONNECTED_5440, SV2V_UNCONNECTED_5441, SV2V_UNCONNECTED_5442, SV2V_UNCONNECTED_5443, SV2V_UNCONNECTED_5444, SV2V_UNCONNECTED_5445, SV2V_UNCONNECTED_5446, SV2V_UNCONNECTED_5447, SV2V_UNCONNECTED_5448, SV2V_UNCONNECTED_5449, SV2V_UNCONNECTED_5450, SV2V_UNCONNECTED_5451, SV2V_UNCONNECTED_5452, SV2V_UNCONNECTED_5453, SV2V_UNCONNECTED_5454, SV2V_UNCONNECTED_5455, SV2V_UNCONNECTED_5456, SV2V_UNCONNECTED_5457, SV2V_UNCONNECTED_5458, SV2V_UNCONNECTED_5459, SV2V_UNCONNECTED_5460, SV2V_UNCONNECTED_5461, SV2V_UNCONNECTED_5462, SV2V_UNCONNECTED_5463, SV2V_UNCONNECTED_5464, SV2V_UNCONNECTED_5465, SV2V_UNCONNECTED_5466, SV2V_UNCONNECTED_5467, SV2V_UNCONNECTED_5468, SV2V_UNCONNECTED_5469, SV2V_UNCONNECTED_5470, SV2V_UNCONNECTED_5471, SV2V_UNCONNECTED_5472, SV2V_UNCONNECTED_5473, SV2V_UNCONNECTED_5474, SV2V_UNCONNECTED_5475, SV2V_UNCONNECTED_5476, SV2V_UNCONNECTED_5477, SV2V_UNCONNECTED_5478, SV2V_UNCONNECTED_5479, SV2V_UNCONNECTED_5480, SV2V_UNCONNECTED_5481, SV2V_UNCONNECTED_5482, SV2V_UNCONNECTED_5483, SV2V_UNCONNECTED_5484, SV2V_UNCONNECTED_5485, SV2V_UNCONNECTED_5486, SV2V_UNCONNECTED_5487, SV2V_UNCONNECTED_5488, SV2V_UNCONNECTED_5489, SV2V_UNCONNECTED_5490, SV2V_UNCONNECTED_5491, SV2V_UNCONNECTED_5492, SV2V_UNCONNECTED_5493, SV2V_UNCONNECTED_5494, SV2V_UNCONNECTED_5495, SV2V_UNCONNECTED_5496, SV2V_UNCONNECTED_5497, SV2V_UNCONNECTED_5498, SV2V_UNCONNECTED_5499, SV2V_UNCONNECTED_5500, SV2V_UNCONNECTED_5501, SV2V_UNCONNECTED_5502, SV2V_UNCONNECTED_5503, SV2V_UNCONNECTED_5504, SV2V_UNCONNECTED_5505, SV2V_UNCONNECTED_5506, SV2V_UNCONNECTED_5507, SV2V_UNCONNECTED_5508, SV2V_UNCONNECTED_5509, SV2V_UNCONNECTED_5510, SV2V_UNCONNECTED_5511, SV2V_UNCONNECTED_5512, SV2V_UNCONNECTED_5513, SV2V_UNCONNECTED_5514, SV2V_UNCONNECTED_5515, SV2V_UNCONNECTED_5516, SV2V_UNCONNECTED_5517, SV2V_UNCONNECTED_5518, SV2V_UNCONNECTED_5519, SV2V_UNCONNECTED_5520, SV2V_UNCONNECTED_5521, SV2V_UNCONNECTED_5522, SV2V_UNCONNECTED_5523, SV2V_UNCONNECTED_5524, SV2V_UNCONNECTED_5525, SV2V_UNCONNECTED_5526, SV2V_UNCONNECTED_5527, SV2V_UNCONNECTED_5528, SV2V_UNCONNECTED_5529, SV2V_UNCONNECTED_5530, SV2V_UNCONNECTED_5531, SV2V_UNCONNECTED_5532, SV2V_UNCONNECTED_5533, SV2V_UNCONNECTED_5534, SV2V_UNCONNECTED_5535, SV2V_UNCONNECTED_5536, SV2V_UNCONNECTED_5537, SV2V_UNCONNECTED_5538, SV2V_UNCONNECTED_5539, SV2V_UNCONNECTED_5540, SV2V_UNCONNECTED_5541, SV2V_UNCONNECTED_5542, SV2V_UNCONNECTED_5543, SV2V_UNCONNECTED_5544, SV2V_UNCONNECTED_5545, SV2V_UNCONNECTED_5546, SV2V_UNCONNECTED_5547, SV2V_UNCONNECTED_5548, SV2V_UNCONNECTED_5549, SV2V_UNCONNECTED_5550, SV2V_UNCONNECTED_5551, SV2V_UNCONNECTED_5552, SV2V_UNCONNECTED_5553, SV2V_UNCONNECTED_5554, SV2V_UNCONNECTED_5555, SV2V_UNCONNECTED_5556, SV2V_UNCONNECTED_5557, SV2V_UNCONNECTED_5558, SV2V_UNCONNECTED_5559, SV2V_UNCONNECTED_5560, SV2V_UNCONNECTED_5561, SV2V_UNCONNECTED_5562, SV2V_UNCONNECTED_5563, SV2V_UNCONNECTED_5564, SV2V_UNCONNECTED_5565, SV2V_UNCONNECTED_5566, SV2V_UNCONNECTED_5567, SV2V_UNCONNECTED_5568, SV2V_UNCONNECTED_5569, SV2V_UNCONNECTED_5570, SV2V_UNCONNECTED_5571, SV2V_UNCONNECTED_5572, SV2V_UNCONNECTED_5573, SV2V_UNCONNECTED_5574, SV2V_UNCONNECTED_5575, SV2V_UNCONNECTED_5576, SV2V_UNCONNECTED_5577, SV2V_UNCONNECTED_5578, SV2V_UNCONNECTED_5579, SV2V_UNCONNECTED_5580, SV2V_UNCONNECTED_5581, SV2V_UNCONNECTED_5582, SV2V_UNCONNECTED_5583, SV2V_UNCONNECTED_5584, SV2V_UNCONNECTED_5585, SV2V_UNCONNECTED_5586, SV2V_UNCONNECTED_5587, SV2V_UNCONNECTED_5588, SV2V_UNCONNECTED_5589, SV2V_UNCONNECTED_5590, SV2V_UNCONNECTED_5591, SV2V_UNCONNECTED_5592, SV2V_UNCONNECTED_5593, SV2V_UNCONNECTED_5594, SV2V_UNCONNECTED_5595, SV2V_UNCONNECTED_5596, SV2V_UNCONNECTED_5597, SV2V_UNCONNECTED_5598, SV2V_UNCONNECTED_5599, SV2V_UNCONNECTED_5600, SV2V_UNCONNECTED_5601, SV2V_UNCONNECTED_5602, SV2V_UNCONNECTED_5603, SV2V_UNCONNECTED_5604, SV2V_UNCONNECTED_5605, SV2V_UNCONNECTED_5606, SV2V_UNCONNECTED_5607, SV2V_UNCONNECTED_5608, SV2V_UNCONNECTED_5609, SV2V_UNCONNECTED_5610, SV2V_UNCONNECTED_5611, SV2V_UNCONNECTED_5612, SV2V_UNCONNECTED_5613, SV2V_UNCONNECTED_5614, SV2V_UNCONNECTED_5615, SV2V_UNCONNECTED_5616, SV2V_UNCONNECTED_5617, SV2V_UNCONNECTED_5618, SV2V_UNCONNECTED_5619, SV2V_UNCONNECTED_5620, SV2V_UNCONNECTED_5621, SV2V_UNCONNECTED_5622, SV2V_UNCONNECTED_5623, SV2V_UNCONNECTED_5624, SV2V_UNCONNECTED_5625, SV2V_UNCONNECTED_5626, SV2V_UNCONNECTED_5627, SV2V_UNCONNECTED_5628, SV2V_UNCONNECTED_5629, SV2V_UNCONNECTED_5630, SV2V_UNCONNECTED_5631, SV2V_UNCONNECTED_5632, SV2V_UNCONNECTED_5633, SV2V_UNCONNECTED_5634, SV2V_UNCONNECTED_5635, SV2V_UNCONNECTED_5636, SV2V_UNCONNECTED_5637, SV2V_UNCONNECTED_5638, SV2V_UNCONNECTED_5639, SV2V_UNCONNECTED_5640, SV2V_UNCONNECTED_5641, SV2V_UNCONNECTED_5642, SV2V_UNCONNECTED_5643, SV2V_UNCONNECTED_5644, SV2V_UNCONNECTED_5645, SV2V_UNCONNECTED_5646, SV2V_UNCONNECTED_5647, SV2V_UNCONNECTED_5648, SV2V_UNCONNECTED_5649, SV2V_UNCONNECTED_5650, SV2V_UNCONNECTED_5651, SV2V_UNCONNECTED_5652, SV2V_UNCONNECTED_5653, SV2V_UNCONNECTED_5654, SV2V_UNCONNECTED_5655, SV2V_UNCONNECTED_5656, SV2V_UNCONNECTED_5657, SV2V_UNCONNECTED_5658, SV2V_UNCONNECTED_5659, SV2V_UNCONNECTED_5660, SV2V_UNCONNECTED_5661, SV2V_UNCONNECTED_5662, SV2V_UNCONNECTED_5663, SV2V_UNCONNECTED_5664, SV2V_UNCONNECTED_5665, SV2V_UNCONNECTED_5666, SV2V_UNCONNECTED_5667, SV2V_UNCONNECTED_5668, SV2V_UNCONNECTED_5669, SV2V_UNCONNECTED_5670, SV2V_UNCONNECTED_5671, SV2V_UNCONNECTED_5672, SV2V_UNCONNECTED_5673, SV2V_UNCONNECTED_5674, SV2V_UNCONNECTED_5675, SV2V_UNCONNECTED_5676, SV2V_UNCONNECTED_5677, SV2V_UNCONNECTED_5678, SV2V_UNCONNECTED_5679, SV2V_UNCONNECTED_5680, SV2V_UNCONNECTED_5681, SV2V_UNCONNECTED_5682, SV2V_UNCONNECTED_5683, SV2V_UNCONNECTED_5684, SV2V_UNCONNECTED_5685, SV2V_UNCONNECTED_5686, SV2V_UNCONNECTED_5687, SV2V_UNCONNECTED_5688, SV2V_UNCONNECTED_5689, SV2V_UNCONNECTED_5690, SV2V_UNCONNECTED_5691, SV2V_UNCONNECTED_5692, SV2V_UNCONNECTED_5693, SV2V_UNCONNECTED_5694, SV2V_UNCONNECTED_5695, SV2V_UNCONNECTED_5696, SV2V_UNCONNECTED_5697, SV2V_UNCONNECTED_5698, SV2V_UNCONNECTED_5699, SV2V_UNCONNECTED_5700, SV2V_UNCONNECTED_5701, SV2V_UNCONNECTED_5702, SV2V_UNCONNECTED_5703, SV2V_UNCONNECTED_5704, SV2V_UNCONNECTED_5705, SV2V_UNCONNECTED_5706, SV2V_UNCONNECTED_5707, SV2V_UNCONNECTED_5708, SV2V_UNCONNECTED_5709, SV2V_UNCONNECTED_5710, SV2V_UNCONNECTED_5711, SV2V_UNCONNECTED_5712, SV2V_UNCONNECTED_5713, SV2V_UNCONNECTED_5714, SV2V_UNCONNECTED_5715, SV2V_UNCONNECTED_5716, SV2V_UNCONNECTED_5717, SV2V_UNCONNECTED_5718, SV2V_UNCONNECTED_5719, SV2V_UNCONNECTED_5720, SV2V_UNCONNECTED_5721, SV2V_UNCONNECTED_5722, SV2V_UNCONNECTED_5723, SV2V_UNCONNECTED_5724, SV2V_UNCONNECTED_5725, SV2V_UNCONNECTED_5726, SV2V_UNCONNECTED_5727, SV2V_UNCONNECTED_5728, SV2V_UNCONNECTED_5729, SV2V_UNCONNECTED_5730, SV2V_UNCONNECTED_5731, SV2V_UNCONNECTED_5732, SV2V_UNCONNECTED_5733, SV2V_UNCONNECTED_5734, SV2V_UNCONNECTED_5735, SV2V_UNCONNECTED_5736, SV2V_UNCONNECTED_5737, SV2V_UNCONNECTED_5738, SV2V_UNCONNECTED_5739, SV2V_UNCONNECTED_5740, SV2V_UNCONNECTED_5741, SV2V_UNCONNECTED_5742, SV2V_UNCONNECTED_5743, SV2V_UNCONNECTED_5744, SV2V_UNCONNECTED_5745, SV2V_UNCONNECTED_5746, SV2V_UNCONNECTED_5747, SV2V_UNCONNECTED_5748, SV2V_UNCONNECTED_5749, SV2V_UNCONNECTED_5750, SV2V_UNCONNECTED_5751, SV2V_UNCONNECTED_5752, SV2V_UNCONNECTED_5753, SV2V_UNCONNECTED_5754, SV2V_UNCONNECTED_5755, SV2V_UNCONNECTED_5756, SV2V_UNCONNECTED_5757, SV2V_UNCONNECTED_5758, SV2V_UNCONNECTED_5759, SV2V_UNCONNECTED_5760, SV2V_UNCONNECTED_5761, SV2V_UNCONNECTED_5762, SV2V_UNCONNECTED_5763, SV2V_UNCONNECTED_5764, SV2V_UNCONNECTED_5765, SV2V_UNCONNECTED_5766, SV2V_UNCONNECTED_5767, SV2V_UNCONNECTED_5768, SV2V_UNCONNECTED_5769, SV2V_UNCONNECTED_5770, SV2V_UNCONNECTED_5771, SV2V_UNCONNECTED_5772, SV2V_UNCONNECTED_5773, SV2V_UNCONNECTED_5774, SV2V_UNCONNECTED_5775, SV2V_UNCONNECTED_5776, SV2V_UNCONNECTED_5777, SV2V_UNCONNECTED_5778, SV2V_UNCONNECTED_5779, SV2V_UNCONNECTED_5780, SV2V_UNCONNECTED_5781, SV2V_UNCONNECTED_5782, SV2V_UNCONNECTED_5783, SV2V_UNCONNECTED_5784, SV2V_UNCONNECTED_5785, SV2V_UNCONNECTED_5786, SV2V_UNCONNECTED_5787, SV2V_UNCONNECTED_5788, SV2V_UNCONNECTED_5789, SV2V_UNCONNECTED_5790, SV2V_UNCONNECTED_5791, SV2V_UNCONNECTED_5792, SV2V_UNCONNECTED_5793, SV2V_UNCONNECTED_5794, SV2V_UNCONNECTED_5795, SV2V_UNCONNECTED_5796, SV2V_UNCONNECTED_5797, SV2V_UNCONNECTED_5798, SV2V_UNCONNECTED_5799, SV2V_UNCONNECTED_5800, SV2V_UNCONNECTED_5801, SV2V_UNCONNECTED_5802, SV2V_UNCONNECTED_5803, SV2V_UNCONNECTED_5804, SV2V_UNCONNECTED_5805, SV2V_UNCONNECTED_5806, SV2V_UNCONNECTED_5807, SV2V_UNCONNECTED_5808, SV2V_UNCONNECTED_5809, SV2V_UNCONNECTED_5810, SV2V_UNCONNECTED_5811, SV2V_UNCONNECTED_5812, SV2V_UNCONNECTED_5813, SV2V_UNCONNECTED_5814, SV2V_UNCONNECTED_5815, SV2V_UNCONNECTED_5816, SV2V_UNCONNECTED_5817, SV2V_UNCONNECTED_5818, SV2V_UNCONNECTED_5819, SV2V_UNCONNECTED_5820, SV2V_UNCONNECTED_5821, SV2V_UNCONNECTED_5822, SV2V_UNCONNECTED_5823, SV2V_UNCONNECTED_5824, SV2V_UNCONNECTED_5825, SV2V_UNCONNECTED_5826, SV2V_UNCONNECTED_5827, SV2V_UNCONNECTED_5828, SV2V_UNCONNECTED_5829, SV2V_UNCONNECTED_5830, SV2V_UNCONNECTED_5831, SV2V_UNCONNECTED_5832, SV2V_UNCONNECTED_5833, SV2V_UNCONNECTED_5834, SV2V_UNCONNECTED_5835, SV2V_UNCONNECTED_5836, SV2V_UNCONNECTED_5837, SV2V_UNCONNECTED_5838, SV2V_UNCONNECTED_5839, SV2V_UNCONNECTED_5840, SV2V_UNCONNECTED_5841, SV2V_UNCONNECTED_5842, SV2V_UNCONNECTED_5843, SV2V_UNCONNECTED_5844, SV2V_UNCONNECTED_5845, SV2V_UNCONNECTED_5846, SV2V_UNCONNECTED_5847, SV2V_UNCONNECTED_5848, SV2V_UNCONNECTED_5849, SV2V_UNCONNECTED_5850, SV2V_UNCONNECTED_5851, SV2V_UNCONNECTED_5852, SV2V_UNCONNECTED_5853, SV2V_UNCONNECTED_5854, SV2V_UNCONNECTED_5855, SV2V_UNCONNECTED_5856, SV2V_UNCONNECTED_5857, SV2V_UNCONNECTED_5858, SV2V_UNCONNECTED_5859, SV2V_UNCONNECTED_5860, SV2V_UNCONNECTED_5861, SV2V_UNCONNECTED_5862, SV2V_UNCONNECTED_5863, SV2V_UNCONNECTED_5864, SV2V_UNCONNECTED_5865, SV2V_UNCONNECTED_5866, SV2V_UNCONNECTED_5867, SV2V_UNCONNECTED_5868, SV2V_UNCONNECTED_5869, SV2V_UNCONNECTED_5870, SV2V_UNCONNECTED_5871, SV2V_UNCONNECTED_5872, SV2V_UNCONNECTED_5873, SV2V_UNCONNECTED_5874, SV2V_UNCONNECTED_5875, SV2V_UNCONNECTED_5876, SV2V_UNCONNECTED_5877, SV2V_UNCONNECTED_5878, SV2V_UNCONNECTED_5879, SV2V_UNCONNECTED_5880, SV2V_UNCONNECTED_5881, SV2V_UNCONNECTED_5882, SV2V_UNCONNECTED_5883, SV2V_UNCONNECTED_5884, SV2V_UNCONNECTED_5885, SV2V_UNCONNECTED_5886, SV2V_UNCONNECTED_5887, SV2V_UNCONNECTED_5888, SV2V_UNCONNECTED_5889, SV2V_UNCONNECTED_5890, SV2V_UNCONNECTED_5891, SV2V_UNCONNECTED_5892, SV2V_UNCONNECTED_5893, SV2V_UNCONNECTED_5894, SV2V_UNCONNECTED_5895, SV2V_UNCONNECTED_5896, SV2V_UNCONNECTED_5897, SV2V_UNCONNECTED_5898, SV2V_UNCONNECTED_5899, SV2V_UNCONNECTED_5900, SV2V_UNCONNECTED_5901, SV2V_UNCONNECTED_5902, SV2V_UNCONNECTED_5903, SV2V_UNCONNECTED_5904, SV2V_UNCONNECTED_5905, SV2V_UNCONNECTED_5906, SV2V_UNCONNECTED_5907, SV2V_UNCONNECTED_5908, SV2V_UNCONNECTED_5909, SV2V_UNCONNECTED_5910, SV2V_UNCONNECTED_5911, SV2V_UNCONNECTED_5912, SV2V_UNCONNECTED_5913, SV2V_UNCONNECTED_5914, SV2V_UNCONNECTED_5915, SV2V_UNCONNECTED_5916, SV2V_UNCONNECTED_5917, SV2V_UNCONNECTED_5918, SV2V_UNCONNECTED_5919, SV2V_UNCONNECTED_5920, SV2V_UNCONNECTED_5921, SV2V_UNCONNECTED_5922, SV2V_UNCONNECTED_5923, SV2V_UNCONNECTED_5924, SV2V_UNCONNECTED_5925, SV2V_UNCONNECTED_5926, SV2V_UNCONNECTED_5927, SV2V_UNCONNECTED_5928, SV2V_UNCONNECTED_5929, SV2V_UNCONNECTED_5930, SV2V_UNCONNECTED_5931, SV2V_UNCONNECTED_5932, SV2V_UNCONNECTED_5933, SV2V_UNCONNECTED_5934, SV2V_UNCONNECTED_5935, SV2V_UNCONNECTED_5936, SV2V_UNCONNECTED_5937, SV2V_UNCONNECTED_5938, SV2V_UNCONNECTED_5939, SV2V_UNCONNECTED_5940, SV2V_UNCONNECTED_5941, SV2V_UNCONNECTED_5942, SV2V_UNCONNECTED_5943, SV2V_UNCONNECTED_5944, SV2V_UNCONNECTED_5945, SV2V_UNCONNECTED_5946, SV2V_UNCONNECTED_5947, SV2V_UNCONNECTED_5948, SV2V_UNCONNECTED_5949, SV2V_UNCONNECTED_5950, SV2V_UNCONNECTED_5951, SV2V_UNCONNECTED_5952, SV2V_UNCONNECTED_5953, SV2V_UNCONNECTED_5954, SV2V_UNCONNECTED_5955, SV2V_UNCONNECTED_5956, SV2V_UNCONNECTED_5957, SV2V_UNCONNECTED_5958, SV2V_UNCONNECTED_5959, SV2V_UNCONNECTED_5960, SV2V_UNCONNECTED_5961, SV2V_UNCONNECTED_5962, SV2V_UNCONNECTED_5963, SV2V_UNCONNECTED_5964, SV2V_UNCONNECTED_5965, SV2V_UNCONNECTED_5966, SV2V_UNCONNECTED_5967, SV2V_UNCONNECTED_5968, SV2V_UNCONNECTED_5969, SV2V_UNCONNECTED_5970, SV2V_UNCONNECTED_5971, SV2V_UNCONNECTED_5972, SV2V_UNCONNECTED_5973, SV2V_UNCONNECTED_5974, SV2V_UNCONNECTED_5975, SV2V_UNCONNECTED_5976, SV2V_UNCONNECTED_5977, SV2V_UNCONNECTED_5978, SV2V_UNCONNECTED_5979, SV2V_UNCONNECTED_5980, SV2V_UNCONNECTED_5981, SV2V_UNCONNECTED_5982, SV2V_UNCONNECTED_5983, SV2V_UNCONNECTED_5984, SV2V_UNCONNECTED_5985, SV2V_UNCONNECTED_5986, SV2V_UNCONNECTED_5987, SV2V_UNCONNECTED_5988, SV2V_UNCONNECTED_5989, SV2V_UNCONNECTED_5990, SV2V_UNCONNECTED_5991, SV2V_UNCONNECTED_5992, SV2V_UNCONNECTED_5993, SV2V_UNCONNECTED_5994, SV2V_UNCONNECTED_5995, SV2V_UNCONNECTED_5996, SV2V_UNCONNECTED_5997, SV2V_UNCONNECTED_5998, SV2V_UNCONNECTED_5999, SV2V_UNCONNECTED_6000, SV2V_UNCONNECTED_6001, SV2V_UNCONNECTED_6002, SV2V_UNCONNECTED_6003, SV2V_UNCONNECTED_6004, SV2V_UNCONNECTED_6005, SV2V_UNCONNECTED_6006, SV2V_UNCONNECTED_6007, SV2V_UNCONNECTED_6008, SV2V_UNCONNECTED_6009, SV2V_UNCONNECTED_6010, SV2V_UNCONNECTED_6011, SV2V_UNCONNECTED_6012, SV2V_UNCONNECTED_6013, SV2V_UNCONNECTED_6014, SV2V_UNCONNECTED_6015, SV2V_UNCONNECTED_6016, SV2V_UNCONNECTED_6017, SV2V_UNCONNECTED_6018, SV2V_UNCONNECTED_6019, SV2V_UNCONNECTED_6020, SV2V_UNCONNECTED_6021, SV2V_UNCONNECTED_6022, SV2V_UNCONNECTED_6023, SV2V_UNCONNECTED_6024, SV2V_UNCONNECTED_6025, SV2V_UNCONNECTED_6026, SV2V_UNCONNECTED_6027, SV2V_UNCONNECTED_6028, SV2V_UNCONNECTED_6029, SV2V_UNCONNECTED_6030, SV2V_UNCONNECTED_6031, SV2V_UNCONNECTED_6032, SV2V_UNCONNECTED_6033, SV2V_UNCONNECTED_6034, SV2V_UNCONNECTED_6035, SV2V_UNCONNECTED_6036, SV2V_UNCONNECTED_6037, SV2V_UNCONNECTED_6038, SV2V_UNCONNECTED_6039, SV2V_UNCONNECTED_6040, SV2V_UNCONNECTED_6041, SV2V_UNCONNECTED_6042, SV2V_UNCONNECTED_6043, SV2V_UNCONNECTED_6044, SV2V_UNCONNECTED_6045, SV2V_UNCONNECTED_6046, SV2V_UNCONNECTED_6047, SV2V_UNCONNECTED_6048, SV2V_UNCONNECTED_6049, SV2V_UNCONNECTED_6050, SV2V_UNCONNECTED_6051, SV2V_UNCONNECTED_6052, SV2V_UNCONNECTED_6053, SV2V_UNCONNECTED_6054, SV2V_UNCONNECTED_6055, SV2V_UNCONNECTED_6056, SV2V_UNCONNECTED_6057, SV2V_UNCONNECTED_6058, SV2V_UNCONNECTED_6059, SV2V_UNCONNECTED_6060, SV2V_UNCONNECTED_6061, SV2V_UNCONNECTED_6062, SV2V_UNCONNECTED_6063, SV2V_UNCONNECTED_6064, SV2V_UNCONNECTED_6065, SV2V_UNCONNECTED_6066, SV2V_UNCONNECTED_6067, SV2V_UNCONNECTED_6068, SV2V_UNCONNECTED_6069, SV2V_UNCONNECTED_6070, SV2V_UNCONNECTED_6071, SV2V_UNCONNECTED_6072, SV2V_UNCONNECTED_6073, SV2V_UNCONNECTED_6074, SV2V_UNCONNECTED_6075, SV2V_UNCONNECTED_6076, SV2V_UNCONNECTED_6077, SV2V_UNCONNECTED_6078, SV2V_UNCONNECTED_6079, SV2V_UNCONNECTED_6080, SV2V_UNCONNECTED_6081, SV2V_UNCONNECTED_6082, SV2V_UNCONNECTED_6083, SV2V_UNCONNECTED_6084, SV2V_UNCONNECTED_6085, SV2V_UNCONNECTED_6086, SV2V_UNCONNECTED_6087, SV2V_UNCONNECTED_6088, SV2V_UNCONNECTED_6089, SV2V_UNCONNECTED_6090, SV2V_UNCONNECTED_6091, SV2V_UNCONNECTED_6092, SV2V_UNCONNECTED_6093, SV2V_UNCONNECTED_6094, SV2V_UNCONNECTED_6095, SV2V_UNCONNECTED_6096, SV2V_UNCONNECTED_6097, SV2V_UNCONNECTED_6098, SV2V_UNCONNECTED_6099, SV2V_UNCONNECTED_6100, SV2V_UNCONNECTED_6101, SV2V_UNCONNECTED_6102, SV2V_UNCONNECTED_6103, SV2V_UNCONNECTED_6104, SV2V_UNCONNECTED_6105, SV2V_UNCONNECTED_6106, SV2V_UNCONNECTED_6107, SV2V_UNCONNECTED_6108, SV2V_UNCONNECTED_6109, SV2V_UNCONNECTED_6110, SV2V_UNCONNECTED_6111, SV2V_UNCONNECTED_6112, SV2V_UNCONNECTED_6113, SV2V_UNCONNECTED_6114, SV2V_UNCONNECTED_6115, SV2V_UNCONNECTED_6116, SV2V_UNCONNECTED_6117, SV2V_UNCONNECTED_6118, SV2V_UNCONNECTED_6119, SV2V_UNCONNECTED_6120, SV2V_UNCONNECTED_6121, SV2V_UNCONNECTED_6122, SV2V_UNCONNECTED_6123, SV2V_UNCONNECTED_6124, SV2V_UNCONNECTED_6125, SV2V_UNCONNECTED_6126, SV2V_UNCONNECTED_6127, SV2V_UNCONNECTED_6128, SV2V_UNCONNECTED_6129, SV2V_UNCONNECTED_6130, SV2V_UNCONNECTED_6131, SV2V_UNCONNECTED_6132, SV2V_UNCONNECTED_6133, SV2V_UNCONNECTED_6134, SV2V_UNCONNECTED_6135, SV2V_UNCONNECTED_6136, SV2V_UNCONNECTED_6137, SV2V_UNCONNECTED_6138, SV2V_UNCONNECTED_6139, SV2V_UNCONNECTED_6140, SV2V_UNCONNECTED_6141, SV2V_UNCONNECTED_6142, SV2V_UNCONNECTED_6143, SV2V_UNCONNECTED_6144, SV2V_UNCONNECTED_6145, SV2V_UNCONNECTED_6146, SV2V_UNCONNECTED_6147, SV2V_UNCONNECTED_6148, SV2V_UNCONNECTED_6149, SV2V_UNCONNECTED_6150, SV2V_UNCONNECTED_6151, SV2V_UNCONNECTED_6152, SV2V_UNCONNECTED_6153, SV2V_UNCONNECTED_6154, SV2V_UNCONNECTED_6155, SV2V_UNCONNECTED_6156, SV2V_UNCONNECTED_6157, SV2V_UNCONNECTED_6158, SV2V_UNCONNECTED_6159, SV2V_UNCONNECTED_6160, SV2V_UNCONNECTED_6161, SV2V_UNCONNECTED_6162, SV2V_UNCONNECTED_6163, SV2V_UNCONNECTED_6164, SV2V_UNCONNECTED_6165, SV2V_UNCONNECTED_6166, SV2V_UNCONNECTED_6167, SV2V_UNCONNECTED_6168, SV2V_UNCONNECTED_6169, SV2V_UNCONNECTED_6170, SV2V_UNCONNECTED_6171, SV2V_UNCONNECTED_6172, SV2V_UNCONNECTED_6173, SV2V_UNCONNECTED_6174, SV2V_UNCONNECTED_6175, SV2V_UNCONNECTED_6176, SV2V_UNCONNECTED_6177, SV2V_UNCONNECTED_6178, SV2V_UNCONNECTED_6179, SV2V_UNCONNECTED_6180, SV2V_UNCONNECTED_6181, SV2V_UNCONNECTED_6182, SV2V_UNCONNECTED_6183, SV2V_UNCONNECTED_6184, SV2V_UNCONNECTED_6185, SV2V_UNCONNECTED_6186, SV2V_UNCONNECTED_6187, SV2V_UNCONNECTED_6188, SV2V_UNCONNECTED_6189, SV2V_UNCONNECTED_6190, SV2V_UNCONNECTED_6191, SV2V_UNCONNECTED_6192, SV2V_UNCONNECTED_6193, SV2V_UNCONNECTED_6194, SV2V_UNCONNECTED_6195, SV2V_UNCONNECTED_6196, SV2V_UNCONNECTED_6197, SV2V_UNCONNECTED_6198, SV2V_UNCONNECTED_6199, SV2V_UNCONNECTED_6200, SV2V_UNCONNECTED_6201, SV2V_UNCONNECTED_6202, SV2V_UNCONNECTED_6203, SV2V_UNCONNECTED_6204, SV2V_UNCONNECTED_6205, SV2V_UNCONNECTED_6206, SV2V_UNCONNECTED_6207, SV2V_UNCONNECTED_6208, SV2V_UNCONNECTED_6209, SV2V_UNCONNECTED_6210, SV2V_UNCONNECTED_6211, SV2V_UNCONNECTED_6212, SV2V_UNCONNECTED_6213, SV2V_UNCONNECTED_6214, SV2V_UNCONNECTED_6215, SV2V_UNCONNECTED_6216, SV2V_UNCONNECTED_6217, SV2V_UNCONNECTED_6218, SV2V_UNCONNECTED_6219, SV2V_UNCONNECTED_6220, SV2V_UNCONNECTED_6221, SV2V_UNCONNECTED_6222, SV2V_UNCONNECTED_6223, SV2V_UNCONNECTED_6224, SV2V_UNCONNECTED_6225, SV2V_UNCONNECTED_6226, SV2V_UNCONNECTED_6227, SV2V_UNCONNECTED_6228, SV2V_UNCONNECTED_6229, SV2V_UNCONNECTED_6230, SV2V_UNCONNECTED_6231, SV2V_UNCONNECTED_6232, SV2V_UNCONNECTED_6233, SV2V_UNCONNECTED_6234, SV2V_UNCONNECTED_6235, SV2V_UNCONNECTED_6236, SV2V_UNCONNECTED_6237, SV2V_UNCONNECTED_6238, SV2V_UNCONNECTED_6239, SV2V_UNCONNECTED_6240, SV2V_UNCONNECTED_6241, SV2V_UNCONNECTED_6242, SV2V_UNCONNECTED_6243, SV2V_UNCONNECTED_6244, SV2V_UNCONNECTED_6245, SV2V_UNCONNECTED_6246, SV2V_UNCONNECTED_6247, SV2V_UNCONNECTED_6248, SV2V_UNCONNECTED_6249, SV2V_UNCONNECTED_6250, SV2V_UNCONNECTED_6251, SV2V_UNCONNECTED_6252, SV2V_UNCONNECTED_6253, SV2V_UNCONNECTED_6254, SV2V_UNCONNECTED_6255, SV2V_UNCONNECTED_6256, SV2V_UNCONNECTED_6257, SV2V_UNCONNECTED_6258, SV2V_UNCONNECTED_6259, SV2V_UNCONNECTED_6260, SV2V_UNCONNECTED_6261, SV2V_UNCONNECTED_6262, SV2V_UNCONNECTED_6263, SV2V_UNCONNECTED_6264, SV2V_UNCONNECTED_6265, SV2V_UNCONNECTED_6266, SV2V_UNCONNECTED_6267, SV2V_UNCONNECTED_6268, SV2V_UNCONNECTED_6269, SV2V_UNCONNECTED_6270, SV2V_UNCONNECTED_6271, SV2V_UNCONNECTED_6272, SV2V_UNCONNECTED_6273, SV2V_UNCONNECTED_6274, SV2V_UNCONNECTED_6275, SV2V_UNCONNECTED_6276, SV2V_UNCONNECTED_6277, SV2V_UNCONNECTED_6278, SV2V_UNCONNECTED_6279, SV2V_UNCONNECTED_6280, SV2V_UNCONNECTED_6281, SV2V_UNCONNECTED_6282, SV2V_UNCONNECTED_6283, SV2V_UNCONNECTED_6284, SV2V_UNCONNECTED_6285, SV2V_UNCONNECTED_6286, SV2V_UNCONNECTED_6287, SV2V_UNCONNECTED_6288, SV2V_UNCONNECTED_6289, SV2V_UNCONNECTED_6290, SV2V_UNCONNECTED_6291, SV2V_UNCONNECTED_6292, SV2V_UNCONNECTED_6293, SV2V_UNCONNECTED_6294, SV2V_UNCONNECTED_6295, SV2V_UNCONNECTED_6296, SV2V_UNCONNECTED_6297, SV2V_UNCONNECTED_6298, SV2V_UNCONNECTED_6299, SV2V_UNCONNECTED_6300, SV2V_UNCONNECTED_6301, SV2V_UNCONNECTED_6302, SV2V_UNCONNECTED_6303, SV2V_UNCONNECTED_6304, SV2V_UNCONNECTED_6305, SV2V_UNCONNECTED_6306, SV2V_UNCONNECTED_6307, SV2V_UNCONNECTED_6308, SV2V_UNCONNECTED_6309, SV2V_UNCONNECTED_6310, SV2V_UNCONNECTED_6311, SV2V_UNCONNECTED_6312, SV2V_UNCONNECTED_6313, SV2V_UNCONNECTED_6314, SV2V_UNCONNECTED_6315, SV2V_UNCONNECTED_6316, SV2V_UNCONNECTED_6317, SV2V_UNCONNECTED_6318, SV2V_UNCONNECTED_6319, SV2V_UNCONNECTED_6320, SV2V_UNCONNECTED_6321, SV2V_UNCONNECTED_6322, SV2V_UNCONNECTED_6323, SV2V_UNCONNECTED_6324, SV2V_UNCONNECTED_6325, SV2V_UNCONNECTED_6326, SV2V_UNCONNECTED_6327, SV2V_UNCONNECTED_6328, SV2V_UNCONNECTED_6329, SV2V_UNCONNECTED_6330, SV2V_UNCONNECTED_6331, SV2V_UNCONNECTED_6332, SV2V_UNCONNECTED_6333, SV2V_UNCONNECTED_6334, SV2V_UNCONNECTED_6335, SV2V_UNCONNECTED_6336, SV2V_UNCONNECTED_6337, SV2V_UNCONNECTED_6338, SV2V_UNCONNECTED_6339, SV2V_UNCONNECTED_6340, SV2V_UNCONNECTED_6341, SV2V_UNCONNECTED_6342, SV2V_UNCONNECTED_6343, SV2V_UNCONNECTED_6344, SV2V_UNCONNECTED_6345, SV2V_UNCONNECTED_6346, SV2V_UNCONNECTED_6347, SV2V_UNCONNECTED_6348, SV2V_UNCONNECTED_6349, SV2V_UNCONNECTED_6350, SV2V_UNCONNECTED_6351, SV2V_UNCONNECTED_6352, SV2V_UNCONNECTED_6353, SV2V_UNCONNECTED_6354, SV2V_UNCONNECTED_6355, SV2V_UNCONNECTED_6356, SV2V_UNCONNECTED_6357, SV2V_UNCONNECTED_6358, SV2V_UNCONNECTED_6359, SV2V_UNCONNECTED_6360, SV2V_UNCONNECTED_6361, SV2V_UNCONNECTED_6362, SV2V_UNCONNECTED_6363, SV2V_UNCONNECTED_6364, SV2V_UNCONNECTED_6365, SV2V_UNCONNECTED_6366, SV2V_UNCONNECTED_6367, SV2V_UNCONNECTED_6368, SV2V_UNCONNECTED_6369, SV2V_UNCONNECTED_6370, SV2V_UNCONNECTED_6371, SV2V_UNCONNECTED_6372, SV2V_UNCONNECTED_6373, SV2V_UNCONNECTED_6374, SV2V_UNCONNECTED_6375, SV2V_UNCONNECTED_6376, SV2V_UNCONNECTED_6377, SV2V_UNCONNECTED_6378, SV2V_UNCONNECTED_6379, SV2V_UNCONNECTED_6380, SV2V_UNCONNECTED_6381, SV2V_UNCONNECTED_6382, SV2V_UNCONNECTED_6383, SV2V_UNCONNECTED_6384, SV2V_UNCONNECTED_6385, SV2V_UNCONNECTED_6386, SV2V_UNCONNECTED_6387, SV2V_UNCONNECTED_6388, SV2V_UNCONNECTED_6389, SV2V_UNCONNECTED_6390, SV2V_UNCONNECTED_6391, SV2V_UNCONNECTED_6392, SV2V_UNCONNECTED_6393, SV2V_UNCONNECTED_6394, SV2V_UNCONNECTED_6395, SV2V_UNCONNECTED_6396, SV2V_UNCONNECTED_6397, SV2V_UNCONNECTED_6398, SV2V_UNCONNECTED_6399, SV2V_UNCONNECTED_6400, SV2V_UNCONNECTED_6401, SV2V_UNCONNECTED_6402, SV2V_UNCONNECTED_6403, SV2V_UNCONNECTED_6404, SV2V_UNCONNECTED_6405, SV2V_UNCONNECTED_6406, SV2V_UNCONNECTED_6407, SV2V_UNCONNECTED_6408, SV2V_UNCONNECTED_6409, SV2V_UNCONNECTED_6410, SV2V_UNCONNECTED_6411, SV2V_UNCONNECTED_6412, SV2V_UNCONNECTED_6413, SV2V_UNCONNECTED_6414, SV2V_UNCONNECTED_6415, SV2V_UNCONNECTED_6416, SV2V_UNCONNECTED_6417, SV2V_UNCONNECTED_6418, SV2V_UNCONNECTED_6419, SV2V_UNCONNECTED_6420, SV2V_UNCONNECTED_6421, SV2V_UNCONNECTED_6422, SV2V_UNCONNECTED_6423, SV2V_UNCONNECTED_6424, SV2V_UNCONNECTED_6425, SV2V_UNCONNECTED_6426, SV2V_UNCONNECTED_6427, SV2V_UNCONNECTED_6428, SV2V_UNCONNECTED_6429, SV2V_UNCONNECTED_6430, SV2V_UNCONNECTED_6431, SV2V_UNCONNECTED_6432, SV2V_UNCONNECTED_6433, SV2V_UNCONNECTED_6434, SV2V_UNCONNECTED_6435, SV2V_UNCONNECTED_6436, SV2V_UNCONNECTED_6437, SV2V_UNCONNECTED_6438, SV2V_UNCONNECTED_6439, SV2V_UNCONNECTED_6440, SV2V_UNCONNECTED_6441, SV2V_UNCONNECTED_6442, SV2V_UNCONNECTED_6443, SV2V_UNCONNECTED_6444, SV2V_UNCONNECTED_6445, SV2V_UNCONNECTED_6446, SV2V_UNCONNECTED_6447, SV2V_UNCONNECTED_6448, SV2V_UNCONNECTED_6449, SV2V_UNCONNECTED_6450, SV2V_UNCONNECTED_6451, SV2V_UNCONNECTED_6452, SV2V_UNCONNECTED_6453, SV2V_UNCONNECTED_6454, SV2V_UNCONNECTED_6455, SV2V_UNCONNECTED_6456, SV2V_UNCONNECTED_6457, SV2V_UNCONNECTED_6458, SV2V_UNCONNECTED_6459, SV2V_UNCONNECTED_6460, SV2V_UNCONNECTED_6461, SV2V_UNCONNECTED_6462, SV2V_UNCONNECTED_6463, SV2V_UNCONNECTED_6464, SV2V_UNCONNECTED_6465, SV2V_UNCONNECTED_6466, SV2V_UNCONNECTED_6467, SV2V_UNCONNECTED_6468, SV2V_UNCONNECTED_6469, SV2V_UNCONNECTED_6470, SV2V_UNCONNECTED_6471, SV2V_UNCONNECTED_6472, SV2V_UNCONNECTED_6473, SV2V_UNCONNECTED_6474, SV2V_UNCONNECTED_6475, SV2V_UNCONNECTED_6476, SV2V_UNCONNECTED_6477, SV2V_UNCONNECTED_6478, SV2V_UNCONNECTED_6479, SV2V_UNCONNECTED_6480, SV2V_UNCONNECTED_6481, SV2V_UNCONNECTED_6482, SV2V_UNCONNECTED_6483, SV2V_UNCONNECTED_6484, SV2V_UNCONNECTED_6485, SV2V_UNCONNECTED_6486, SV2V_UNCONNECTED_6487, SV2V_UNCONNECTED_6488, SV2V_UNCONNECTED_6489, SV2V_UNCONNECTED_6490, SV2V_UNCONNECTED_6491, SV2V_UNCONNECTED_6492, SV2V_UNCONNECTED_6493, SV2V_UNCONNECTED_6494, SV2V_UNCONNECTED_6495, SV2V_UNCONNECTED_6496, SV2V_UNCONNECTED_6497, SV2V_UNCONNECTED_6498, SV2V_UNCONNECTED_6499, SV2V_UNCONNECTED_6500, SV2V_UNCONNECTED_6501, SV2V_UNCONNECTED_6502, SV2V_UNCONNECTED_6503, SV2V_UNCONNECTED_6504, SV2V_UNCONNECTED_6505, SV2V_UNCONNECTED_6506, SV2V_UNCONNECTED_6507, SV2V_UNCONNECTED_6508, SV2V_UNCONNECTED_6509, SV2V_UNCONNECTED_6510, SV2V_UNCONNECTED_6511, SV2V_UNCONNECTED_6512, SV2V_UNCONNECTED_6513, SV2V_UNCONNECTED_6514, SV2V_UNCONNECTED_6515, SV2V_UNCONNECTED_6516, SV2V_UNCONNECTED_6517, SV2V_UNCONNECTED_6518, SV2V_UNCONNECTED_6519, SV2V_UNCONNECTED_6520, SV2V_UNCONNECTED_6521, SV2V_UNCONNECTED_6522, SV2V_UNCONNECTED_6523, SV2V_UNCONNECTED_6524, SV2V_UNCONNECTED_6525, SV2V_UNCONNECTED_6526, SV2V_UNCONNECTED_6527, SV2V_UNCONNECTED_6528, SV2V_UNCONNECTED_6529, SV2V_UNCONNECTED_6530, SV2V_UNCONNECTED_6531, SV2V_UNCONNECTED_6532, SV2V_UNCONNECTED_6533, SV2V_UNCONNECTED_6534, SV2V_UNCONNECTED_6535, SV2V_UNCONNECTED_6536, SV2V_UNCONNECTED_6537, SV2V_UNCONNECTED_6538, SV2V_UNCONNECTED_6539, SV2V_UNCONNECTED_6540, SV2V_UNCONNECTED_6541, SV2V_UNCONNECTED_6542, SV2V_UNCONNECTED_6543, SV2V_UNCONNECTED_6544, SV2V_UNCONNECTED_6545, SV2V_UNCONNECTED_6546, SV2V_UNCONNECTED_6547, SV2V_UNCONNECTED_6548, SV2V_UNCONNECTED_6549, SV2V_UNCONNECTED_6550, SV2V_UNCONNECTED_6551, SV2V_UNCONNECTED_6552, SV2V_UNCONNECTED_6553, SV2V_UNCONNECTED_6554, SV2V_UNCONNECTED_6555, SV2V_UNCONNECTED_6556, SV2V_UNCONNECTED_6557, SV2V_UNCONNECTED_6558, SV2V_UNCONNECTED_6559, SV2V_UNCONNECTED_6560, SV2V_UNCONNECTED_6561, SV2V_UNCONNECTED_6562, SV2V_UNCONNECTED_6563, SV2V_UNCONNECTED_6564, SV2V_UNCONNECTED_6565, SV2V_UNCONNECTED_6566, SV2V_UNCONNECTED_6567, SV2V_UNCONNECTED_6568, SV2V_UNCONNECTED_6569, SV2V_UNCONNECTED_6570, SV2V_UNCONNECTED_6571, SV2V_UNCONNECTED_6572, SV2V_UNCONNECTED_6573, SV2V_UNCONNECTED_6574, SV2V_UNCONNECTED_6575, SV2V_UNCONNECTED_6576, SV2V_UNCONNECTED_6577, SV2V_UNCONNECTED_6578, SV2V_UNCONNECTED_6579, SV2V_UNCONNECTED_6580, SV2V_UNCONNECTED_6581, SV2V_UNCONNECTED_6582, SV2V_UNCONNECTED_6583, SV2V_UNCONNECTED_6584, SV2V_UNCONNECTED_6585, SV2V_UNCONNECTED_6586, SV2V_UNCONNECTED_6587, SV2V_UNCONNECTED_6588, SV2V_UNCONNECTED_6589, SV2V_UNCONNECTED_6590, SV2V_UNCONNECTED_6591, SV2V_UNCONNECTED_6592, SV2V_UNCONNECTED_6593, SV2V_UNCONNECTED_6594, SV2V_UNCONNECTED_6595, SV2V_UNCONNECTED_6596, SV2V_UNCONNECTED_6597, SV2V_UNCONNECTED_6598, SV2V_UNCONNECTED_6599, SV2V_UNCONNECTED_6600, SV2V_UNCONNECTED_6601, SV2V_UNCONNECTED_6602, SV2V_UNCONNECTED_6603, SV2V_UNCONNECTED_6604, SV2V_UNCONNECTED_6605, SV2V_UNCONNECTED_6606, SV2V_UNCONNECTED_6607, SV2V_UNCONNECTED_6608, SV2V_UNCONNECTED_6609, SV2V_UNCONNECTED_6610, SV2V_UNCONNECTED_6611, SV2V_UNCONNECTED_6612, SV2V_UNCONNECTED_6613, SV2V_UNCONNECTED_6614, SV2V_UNCONNECTED_6615, SV2V_UNCONNECTED_6616, SV2V_UNCONNECTED_6617, SV2V_UNCONNECTED_6618, SV2V_UNCONNECTED_6619, SV2V_UNCONNECTED_6620, SV2V_UNCONNECTED_6621, SV2V_UNCONNECTED_6622, SV2V_UNCONNECTED_6623, SV2V_UNCONNECTED_6624, SV2V_UNCONNECTED_6625, SV2V_UNCONNECTED_6626, SV2V_UNCONNECTED_6627, SV2V_UNCONNECTED_6628, SV2V_UNCONNECTED_6629, SV2V_UNCONNECTED_6630, SV2V_UNCONNECTED_6631, SV2V_UNCONNECTED_6632, SV2V_UNCONNECTED_6633, SV2V_UNCONNECTED_6634, SV2V_UNCONNECTED_6635, SV2V_UNCONNECTED_6636, SV2V_UNCONNECTED_6637, SV2V_UNCONNECTED_6638, SV2V_UNCONNECTED_6639, SV2V_UNCONNECTED_6640, SV2V_UNCONNECTED_6641, SV2V_UNCONNECTED_6642, SV2V_UNCONNECTED_6643, SV2V_UNCONNECTED_6644, SV2V_UNCONNECTED_6645, SV2V_UNCONNECTED_6646, SV2V_UNCONNECTED_6647, SV2V_UNCONNECTED_6648, SV2V_UNCONNECTED_6649, SV2V_UNCONNECTED_6650, SV2V_UNCONNECTED_6651, SV2V_UNCONNECTED_6652, SV2V_UNCONNECTED_6653, SV2V_UNCONNECTED_6654, SV2V_UNCONNECTED_6655, SV2V_UNCONNECTED_6656, SV2V_UNCONNECTED_6657, SV2V_UNCONNECTED_6658, SV2V_UNCONNECTED_6659, SV2V_UNCONNECTED_6660, SV2V_UNCONNECTED_6661, SV2V_UNCONNECTED_6662, SV2V_UNCONNECTED_6663, SV2V_UNCONNECTED_6664, SV2V_UNCONNECTED_6665, SV2V_UNCONNECTED_6666, SV2V_UNCONNECTED_6667, SV2V_UNCONNECTED_6668, SV2V_UNCONNECTED_6669, SV2V_UNCONNECTED_6670, SV2V_UNCONNECTED_6671, SV2V_UNCONNECTED_6672, SV2V_UNCONNECTED_6673, SV2V_UNCONNECTED_6674, SV2V_UNCONNECTED_6675, SV2V_UNCONNECTED_6676, SV2V_UNCONNECTED_6677, SV2V_UNCONNECTED_6678, SV2V_UNCONNECTED_6679, SV2V_UNCONNECTED_6680, SV2V_UNCONNECTED_6681, SV2V_UNCONNECTED_6682, SV2V_UNCONNECTED_6683, SV2V_UNCONNECTED_6684, SV2V_UNCONNECTED_6685, SV2V_UNCONNECTED_6686, SV2V_UNCONNECTED_6687, SV2V_UNCONNECTED_6688, SV2V_UNCONNECTED_6689, SV2V_UNCONNECTED_6690, SV2V_UNCONNECTED_6691, SV2V_UNCONNECTED_6692, SV2V_UNCONNECTED_6693, SV2V_UNCONNECTED_6694, SV2V_UNCONNECTED_6695, SV2V_UNCONNECTED_6696, SV2V_UNCONNECTED_6697, SV2V_UNCONNECTED_6698, SV2V_UNCONNECTED_6699, SV2V_UNCONNECTED_6700, SV2V_UNCONNECTED_6701, SV2V_UNCONNECTED_6702, SV2V_UNCONNECTED_6703, SV2V_UNCONNECTED_6704, SV2V_UNCONNECTED_6705, SV2V_UNCONNECTED_6706, SV2V_UNCONNECTED_6707, SV2V_UNCONNECTED_6708, SV2V_UNCONNECTED_6709, SV2V_UNCONNECTED_6710, SV2V_UNCONNECTED_6711, SV2V_UNCONNECTED_6712, SV2V_UNCONNECTED_6713, SV2V_UNCONNECTED_6714, SV2V_UNCONNECTED_6715, SV2V_UNCONNECTED_6716, SV2V_UNCONNECTED_6717, SV2V_UNCONNECTED_6718, SV2V_UNCONNECTED_6719, SV2V_UNCONNECTED_6720, SV2V_UNCONNECTED_6721, SV2V_UNCONNECTED_6722, SV2V_UNCONNECTED_6723, SV2V_UNCONNECTED_6724, SV2V_UNCONNECTED_6725, SV2V_UNCONNECTED_6726, SV2V_UNCONNECTED_6727, SV2V_UNCONNECTED_6728, SV2V_UNCONNECTED_6729, SV2V_UNCONNECTED_6730, SV2V_UNCONNECTED_6731, SV2V_UNCONNECTED_6732, SV2V_UNCONNECTED_6733, SV2V_UNCONNECTED_6734, SV2V_UNCONNECTED_6735, SV2V_UNCONNECTED_6736, SV2V_UNCONNECTED_6737, SV2V_UNCONNECTED_6738, SV2V_UNCONNECTED_6739, SV2V_UNCONNECTED_6740, SV2V_UNCONNECTED_6741, SV2V_UNCONNECTED_6742, SV2V_UNCONNECTED_6743, SV2V_UNCONNECTED_6744, SV2V_UNCONNECTED_6745, SV2V_UNCONNECTED_6746, SV2V_UNCONNECTED_6747, SV2V_UNCONNECTED_6748, SV2V_UNCONNECTED_6749, SV2V_UNCONNECTED_6750, SV2V_UNCONNECTED_6751, SV2V_UNCONNECTED_6752, SV2V_UNCONNECTED_6753, SV2V_UNCONNECTED_6754, SV2V_UNCONNECTED_6755, SV2V_UNCONNECTED_6756, SV2V_UNCONNECTED_6757, SV2V_UNCONNECTED_6758, SV2V_UNCONNECTED_6759, SV2V_UNCONNECTED_6760, SV2V_UNCONNECTED_6761, SV2V_UNCONNECTED_6762, SV2V_UNCONNECTED_6763, SV2V_UNCONNECTED_6764, SV2V_UNCONNECTED_6765, SV2V_UNCONNECTED_6766, SV2V_UNCONNECTED_6767, SV2V_UNCONNECTED_6768, SV2V_UNCONNECTED_6769, SV2V_UNCONNECTED_6770, SV2V_UNCONNECTED_6771, SV2V_UNCONNECTED_6772, SV2V_UNCONNECTED_6773, SV2V_UNCONNECTED_6774, SV2V_UNCONNECTED_6775, SV2V_UNCONNECTED_6776, SV2V_UNCONNECTED_6777, SV2V_UNCONNECTED_6778, SV2V_UNCONNECTED_6779, SV2V_UNCONNECTED_6780, SV2V_UNCONNECTED_6781, SV2V_UNCONNECTED_6782, SV2V_UNCONNECTED_6783, SV2V_UNCONNECTED_6784, SV2V_UNCONNECTED_6785, SV2V_UNCONNECTED_6786, SV2V_UNCONNECTED_6787, SV2V_UNCONNECTED_6788, SV2V_UNCONNECTED_6789, SV2V_UNCONNECTED_6790, SV2V_UNCONNECTED_6791, SV2V_UNCONNECTED_6792, SV2V_UNCONNECTED_6793, SV2V_UNCONNECTED_6794, SV2V_UNCONNECTED_6795, SV2V_UNCONNECTED_6796, SV2V_UNCONNECTED_6797, SV2V_UNCONNECTED_6798, SV2V_UNCONNECTED_6799, SV2V_UNCONNECTED_6800, SV2V_UNCONNECTED_6801, SV2V_UNCONNECTED_6802, SV2V_UNCONNECTED_6803, SV2V_UNCONNECTED_6804, SV2V_UNCONNECTED_6805, SV2V_UNCONNECTED_6806, SV2V_UNCONNECTED_6807, SV2V_UNCONNECTED_6808, SV2V_UNCONNECTED_6809, SV2V_UNCONNECTED_6810, SV2V_UNCONNECTED_6811, SV2V_UNCONNECTED_6812, SV2V_UNCONNECTED_6813, SV2V_UNCONNECTED_6814, SV2V_UNCONNECTED_6815, SV2V_UNCONNECTED_6816, SV2V_UNCONNECTED_6817, SV2V_UNCONNECTED_6818, SV2V_UNCONNECTED_6819, SV2V_UNCONNECTED_6820, SV2V_UNCONNECTED_6821, SV2V_UNCONNECTED_6822, SV2V_UNCONNECTED_6823, SV2V_UNCONNECTED_6824, SV2V_UNCONNECTED_6825, SV2V_UNCONNECTED_6826, SV2V_UNCONNECTED_6827, SV2V_UNCONNECTED_6828, SV2V_UNCONNECTED_6829, SV2V_UNCONNECTED_6830, SV2V_UNCONNECTED_6831, SV2V_UNCONNECTED_6832, SV2V_UNCONNECTED_6833, SV2V_UNCONNECTED_6834, SV2V_UNCONNECTED_6835, SV2V_UNCONNECTED_6836, SV2V_UNCONNECTED_6837, SV2V_UNCONNECTED_6838, SV2V_UNCONNECTED_6839, SV2V_UNCONNECTED_6840, SV2V_UNCONNECTED_6841, SV2V_UNCONNECTED_6842, SV2V_UNCONNECTED_6843, SV2V_UNCONNECTED_6844, SV2V_UNCONNECTED_6845, SV2V_UNCONNECTED_6846, SV2V_UNCONNECTED_6847, SV2V_UNCONNECTED_6848, SV2V_UNCONNECTED_6849, SV2V_UNCONNECTED_6850, SV2V_UNCONNECTED_6851, SV2V_UNCONNECTED_6852, SV2V_UNCONNECTED_6853, SV2V_UNCONNECTED_6854, SV2V_UNCONNECTED_6855, SV2V_UNCONNECTED_6856, SV2V_UNCONNECTED_6857, SV2V_UNCONNECTED_6858, SV2V_UNCONNECTED_6859, SV2V_UNCONNECTED_6860, SV2V_UNCONNECTED_6861, SV2V_UNCONNECTED_6862, SV2V_UNCONNECTED_6863, SV2V_UNCONNECTED_6864, SV2V_UNCONNECTED_6865, SV2V_UNCONNECTED_6866, SV2V_UNCONNECTED_6867, SV2V_UNCONNECTED_6868, SV2V_UNCONNECTED_6869, SV2V_UNCONNECTED_6870, SV2V_UNCONNECTED_6871, SV2V_UNCONNECTED_6872, SV2V_UNCONNECTED_6873, SV2V_UNCONNECTED_6874, SV2V_UNCONNECTED_6875, SV2V_UNCONNECTED_6876, SV2V_UNCONNECTED_6877, SV2V_UNCONNECTED_6878, SV2V_UNCONNECTED_6879, SV2V_UNCONNECTED_6880, SV2V_UNCONNECTED_6881, SV2V_UNCONNECTED_6882, SV2V_UNCONNECTED_6883, SV2V_UNCONNECTED_6884, SV2V_UNCONNECTED_6885, SV2V_UNCONNECTED_6886, SV2V_UNCONNECTED_6887, SV2V_UNCONNECTED_6888, SV2V_UNCONNECTED_6889, SV2V_UNCONNECTED_6890, SV2V_UNCONNECTED_6891, SV2V_UNCONNECTED_6892, SV2V_UNCONNECTED_6893, SV2V_UNCONNECTED_6894, SV2V_UNCONNECTED_6895, SV2V_UNCONNECTED_6896, SV2V_UNCONNECTED_6897, SV2V_UNCONNECTED_6898, SV2V_UNCONNECTED_6899, SV2V_UNCONNECTED_6900, SV2V_UNCONNECTED_6901, SV2V_UNCONNECTED_6902, SV2V_UNCONNECTED_6903, SV2V_UNCONNECTED_6904, SV2V_UNCONNECTED_6905, SV2V_UNCONNECTED_6906, SV2V_UNCONNECTED_6907, SV2V_UNCONNECTED_6908, SV2V_UNCONNECTED_6909, SV2V_UNCONNECTED_6910, SV2V_UNCONNECTED_6911, SV2V_UNCONNECTED_6912, SV2V_UNCONNECTED_6913, SV2V_UNCONNECTED_6914, SV2V_UNCONNECTED_6915, SV2V_UNCONNECTED_6916, SV2V_UNCONNECTED_6917, SV2V_UNCONNECTED_6918, SV2V_UNCONNECTED_6919, SV2V_UNCONNECTED_6920, SV2V_UNCONNECTED_6921, SV2V_UNCONNECTED_6922, SV2V_UNCONNECTED_6923, SV2V_UNCONNECTED_6924, SV2V_UNCONNECTED_6925, SV2V_UNCONNECTED_6926, SV2V_UNCONNECTED_6927, SV2V_UNCONNECTED_6928, SV2V_UNCONNECTED_6929, SV2V_UNCONNECTED_6930, SV2V_UNCONNECTED_6931, SV2V_UNCONNECTED_6932, SV2V_UNCONNECTED_6933, SV2V_UNCONNECTED_6934, SV2V_UNCONNECTED_6935, SV2V_UNCONNECTED_6936, SV2V_UNCONNECTED_6937, SV2V_UNCONNECTED_6938, SV2V_UNCONNECTED_6939, SV2V_UNCONNECTED_6940, SV2V_UNCONNECTED_6941, SV2V_UNCONNECTED_6942, SV2V_UNCONNECTED_6943, SV2V_UNCONNECTED_6944, SV2V_UNCONNECTED_6945, SV2V_UNCONNECTED_6946, SV2V_UNCONNECTED_6947, SV2V_UNCONNECTED_6948, SV2V_UNCONNECTED_6949, SV2V_UNCONNECTED_6950, SV2V_UNCONNECTED_6951, SV2V_UNCONNECTED_6952, SV2V_UNCONNECTED_6953, SV2V_UNCONNECTED_6954, SV2V_UNCONNECTED_6955, SV2V_UNCONNECTED_6956, SV2V_UNCONNECTED_6957, SV2V_UNCONNECTED_6958, SV2V_UNCONNECTED_6959, SV2V_UNCONNECTED_6960, SV2V_UNCONNECTED_6961, SV2V_UNCONNECTED_6962, SV2V_UNCONNECTED_6963, SV2V_UNCONNECTED_6964, SV2V_UNCONNECTED_6965, SV2V_UNCONNECTED_6966, SV2V_UNCONNECTED_6967, SV2V_UNCONNECTED_6968, SV2V_UNCONNECTED_6969, SV2V_UNCONNECTED_6970, SV2V_UNCONNECTED_6971, SV2V_UNCONNECTED_6972, SV2V_UNCONNECTED_6973, SV2V_UNCONNECTED_6974, SV2V_UNCONNECTED_6975, SV2V_UNCONNECTED_6976, SV2V_UNCONNECTED_6977, SV2V_UNCONNECTED_6978, SV2V_UNCONNECTED_6979, SV2V_UNCONNECTED_6980, SV2V_UNCONNECTED_6981, SV2V_UNCONNECTED_6982, SV2V_UNCONNECTED_6983, SV2V_UNCONNECTED_6984, SV2V_UNCONNECTED_6985, SV2V_UNCONNECTED_6986, SV2V_UNCONNECTED_6987, SV2V_UNCONNECTED_6988, SV2V_UNCONNECTED_6989, SV2V_UNCONNECTED_6990, SV2V_UNCONNECTED_6991, SV2V_UNCONNECTED_6992, SV2V_UNCONNECTED_6993, SV2V_UNCONNECTED_6994, SV2V_UNCONNECTED_6995, SV2V_UNCONNECTED_6996, SV2V_UNCONNECTED_6997, SV2V_UNCONNECTED_6998, SV2V_UNCONNECTED_6999, SV2V_UNCONNECTED_7000, SV2V_UNCONNECTED_7001, SV2V_UNCONNECTED_7002, SV2V_UNCONNECTED_7003, SV2V_UNCONNECTED_7004, SV2V_UNCONNECTED_7005, SV2V_UNCONNECTED_7006, SV2V_UNCONNECTED_7007, SV2V_UNCONNECTED_7008, SV2V_UNCONNECTED_7009, SV2V_UNCONNECTED_7010, SV2V_UNCONNECTED_7011, SV2V_UNCONNECTED_7012, SV2V_UNCONNECTED_7013, SV2V_UNCONNECTED_7014, SV2V_UNCONNECTED_7015, SV2V_UNCONNECTED_7016, SV2V_UNCONNECTED_7017, SV2V_UNCONNECTED_7018, SV2V_UNCONNECTED_7019, SV2V_UNCONNECTED_7020, SV2V_UNCONNECTED_7021, SV2V_UNCONNECTED_7022, SV2V_UNCONNECTED_7023, SV2V_UNCONNECTED_7024, SV2V_UNCONNECTED_7025, SV2V_UNCONNECTED_7026, SV2V_UNCONNECTED_7027, SV2V_UNCONNECTED_7028, SV2V_UNCONNECTED_7029, SV2V_UNCONNECTED_7030, SV2V_UNCONNECTED_7031, SV2V_UNCONNECTED_7032, SV2V_UNCONNECTED_7033, SV2V_UNCONNECTED_7034, SV2V_UNCONNECTED_7035, SV2V_UNCONNECTED_7036, SV2V_UNCONNECTED_7037, SV2V_UNCONNECTED_7038, SV2V_UNCONNECTED_7039, SV2V_UNCONNECTED_7040, SV2V_UNCONNECTED_7041, SV2V_UNCONNECTED_7042, SV2V_UNCONNECTED_7043, SV2V_UNCONNECTED_7044, SV2V_UNCONNECTED_7045, SV2V_UNCONNECTED_7046, SV2V_UNCONNECTED_7047, SV2V_UNCONNECTED_7048, SV2V_UNCONNECTED_7049, SV2V_UNCONNECTED_7050, SV2V_UNCONNECTED_7051, SV2V_UNCONNECTED_7052, SV2V_UNCONNECTED_7053, SV2V_UNCONNECTED_7054, SV2V_UNCONNECTED_7055, SV2V_UNCONNECTED_7056, SV2V_UNCONNECTED_7057, SV2V_UNCONNECTED_7058, SV2V_UNCONNECTED_7059, SV2V_UNCONNECTED_7060, SV2V_UNCONNECTED_7061, SV2V_UNCONNECTED_7062, SV2V_UNCONNECTED_7063, SV2V_UNCONNECTED_7064, SV2V_UNCONNECTED_7065, SV2V_UNCONNECTED_7066, SV2V_UNCONNECTED_7067, SV2V_UNCONNECTED_7068, SV2V_UNCONNECTED_7069, SV2V_UNCONNECTED_7070, SV2V_UNCONNECTED_7071, SV2V_UNCONNECTED_7072, SV2V_UNCONNECTED_7073, SV2V_UNCONNECTED_7074, SV2V_UNCONNECTED_7075, SV2V_UNCONNECTED_7076, SV2V_UNCONNECTED_7077, SV2V_UNCONNECTED_7078, SV2V_UNCONNECTED_7079, SV2V_UNCONNECTED_7080, SV2V_UNCONNECTED_7081, SV2V_UNCONNECTED_7082, SV2V_UNCONNECTED_7083, SV2V_UNCONNECTED_7084, SV2V_UNCONNECTED_7085, SV2V_UNCONNECTED_7086, SV2V_UNCONNECTED_7087, SV2V_UNCONNECTED_7088, SV2V_UNCONNECTED_7089, SV2V_UNCONNECTED_7090, SV2V_UNCONNECTED_7091, SV2V_UNCONNECTED_7092, SV2V_UNCONNECTED_7093, SV2V_UNCONNECTED_7094, SV2V_UNCONNECTED_7095, SV2V_UNCONNECTED_7096, SV2V_UNCONNECTED_7097, SV2V_UNCONNECTED_7098, SV2V_UNCONNECTED_7099, SV2V_UNCONNECTED_7100, SV2V_UNCONNECTED_7101, SV2V_UNCONNECTED_7102, SV2V_UNCONNECTED_7103, SV2V_UNCONNECTED_7104, SV2V_UNCONNECTED_7105, SV2V_UNCONNECTED_7106, SV2V_UNCONNECTED_7107, SV2V_UNCONNECTED_7108, SV2V_UNCONNECTED_7109, SV2V_UNCONNECTED_7110, SV2V_UNCONNECTED_7111, SV2V_UNCONNECTED_7112, SV2V_UNCONNECTED_7113, SV2V_UNCONNECTED_7114, SV2V_UNCONNECTED_7115, SV2V_UNCONNECTED_7116, SV2V_UNCONNECTED_7117, SV2V_UNCONNECTED_7118, SV2V_UNCONNECTED_7119, SV2V_UNCONNECTED_7120, SV2V_UNCONNECTED_7121, SV2V_UNCONNECTED_7122, SV2V_UNCONNECTED_7123, SV2V_UNCONNECTED_7124, SV2V_UNCONNECTED_7125, SV2V_UNCONNECTED_7126, SV2V_UNCONNECTED_7127, SV2V_UNCONNECTED_7128, SV2V_UNCONNECTED_7129, SV2V_UNCONNECTED_7130, SV2V_UNCONNECTED_7131, SV2V_UNCONNECTED_7132, SV2V_UNCONNECTED_7133, SV2V_UNCONNECTED_7134, SV2V_UNCONNECTED_7135, SV2V_UNCONNECTED_7136, SV2V_UNCONNECTED_7137, SV2V_UNCONNECTED_7138, SV2V_UNCONNECTED_7139, SV2V_UNCONNECTED_7140, SV2V_UNCONNECTED_7141, SV2V_UNCONNECTED_7142, SV2V_UNCONNECTED_7143, SV2V_UNCONNECTED_7144, SV2V_UNCONNECTED_7145, SV2V_UNCONNECTED_7146, SV2V_UNCONNECTED_7147, SV2V_UNCONNECTED_7148, SV2V_UNCONNECTED_7149, SV2V_UNCONNECTED_7150, SV2V_UNCONNECTED_7151, SV2V_UNCONNECTED_7152, SV2V_UNCONNECTED_7153, SV2V_UNCONNECTED_7154, SV2V_UNCONNECTED_7155, SV2V_UNCONNECTED_7156, SV2V_UNCONNECTED_7157, SV2V_UNCONNECTED_7158, SV2V_UNCONNECTED_7159, SV2V_UNCONNECTED_7160, SV2V_UNCONNECTED_7161, SV2V_UNCONNECTED_7162, SV2V_UNCONNECTED_7163, SV2V_UNCONNECTED_7164, SV2V_UNCONNECTED_7165, SV2V_UNCONNECTED_7166, SV2V_UNCONNECTED_7167, SV2V_UNCONNECTED_7168, SV2V_UNCONNECTED_7169, SV2V_UNCONNECTED_7170, SV2V_UNCONNECTED_7171, SV2V_UNCONNECTED_7172, SV2V_UNCONNECTED_7173, SV2V_UNCONNECTED_7174, SV2V_UNCONNECTED_7175, SV2V_UNCONNECTED_7176, SV2V_UNCONNECTED_7177, SV2V_UNCONNECTED_7178, SV2V_UNCONNECTED_7179, SV2V_UNCONNECTED_7180, SV2V_UNCONNECTED_7181, SV2V_UNCONNECTED_7182, SV2V_UNCONNECTED_7183, SV2V_UNCONNECTED_7184, SV2V_UNCONNECTED_7185, SV2V_UNCONNECTED_7186, SV2V_UNCONNECTED_7187, SV2V_UNCONNECTED_7188, SV2V_UNCONNECTED_7189, SV2V_UNCONNECTED_7190, SV2V_UNCONNECTED_7191, SV2V_UNCONNECTED_7192, SV2V_UNCONNECTED_7193, SV2V_UNCONNECTED_7194, SV2V_UNCONNECTED_7195, SV2V_UNCONNECTED_7196, SV2V_UNCONNECTED_7197, T9_0, T14[0:0], T15, T16, T17 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> T19;
  assign N641 = N811 | N694;
  assign N642 = T199[10] | T199[11];
  assign N643 = T199[9] | N642;
  assign N644 = T199[8] | N643;
  assign N645 = T199[7] | N644;
  assign N646 = T199[6] | N645;
  assign N647 = T199[5] | N646;
  assign N648 = T199[4] | N647;
  assign N649 = T199[3] | N648;
  assign N650 = T199[2] | N649;
  assign N651 = T199[1] | N650;
  assign N652 = ~N651;
  assign N653 = io_mulAddResult[9] | io_mulAddResult[10];
  assign N654 = io_mulAddResult[8] | N653;
  assign N655 = io_mulAddResult[7] | N654;
  assign N656 = io_mulAddResult[6] | N655;
  assign N657 = io_mulAddResult[5] | N656;
  assign N658 = io_mulAddResult[4] | N657;
  assign N659 = io_mulAddResult[3] | N658;
  assign N660 = io_mulAddResult[2] | N659;
  assign N661 = io_mulAddResult[1] | N660;
  assign N662 = io_mulAddResult[0] | N661;
  assign N663 = N737 | N768;
  assign N664 = notSigSum[74] | notSigSum[75];
  assign N665 = notSigSum[73] | N664;
  assign N666 = notSigSum[72] | N665;
  assign N667 = notSigSum[71] | N666;
  assign N668 = notSigSum[70] | N667;
  assign N669 = notSigSum[69] | N668;
  assign N670 = notSigSum[68] | N669;
  assign N671 = notSigSum[67] | N670;
  assign N672 = notSigSum[66] | N671;
  assign N673 = notSigSum[65] | N672;
  assign N674 = notSigSum[64] | N673;
  assign N675 = notSigSum[63] | N674;
  assign N676 = notSigSum[62] | N675;
  assign N677 = notSigSum[61] | N676;
  assign N678 = notSigSum[60] | N677;
  assign N679 = notSigSum[59] | N678;
  assign N680 = notSigSum[58] | N679;
  assign N681 = notSigSum[57] | N680;
  assign N682 = notSigSum[56] | N681;
  assign N683 = notSigSum[55] | N682;
  assign N684 = notSigSum[54] | N683;
  assign N685 = notSigSum[53] | N684;
  assign N686 = notSigSum[52] | N685;
  assign N687 = notSigSum[51] | N686;
  assign N688 = notSigSum[50] | N687;
  assign N689 = notSigSum[49] | N688;
  assign N690 = notSigSum[48] | N689;
  assign N691 = notSigSum[47] | N690;
  assign N692 = notSigSum[46] | N691;
  assign N693 = notSigSum[45] | N692;
  assign N694 = notSigSum[44] | N693;
  assign N695 = io_mulAddResult[41] | io_mulAddResult[42];
  assign N696 = io_mulAddResult[40] | N695;
  assign N697 = io_mulAddResult[39] | N696;
  assign N698 = io_mulAddResult[38] | N697;
  assign N699 = io_mulAddResult[37] | N698;
  assign N700 = io_mulAddResult[36] | N699;
  assign N701 = io_mulAddResult[35] | N700;
  assign N702 = io_mulAddResult[34] | N701;
  assign N703 = io_mulAddResult[33] | N702;
  assign N704 = io_mulAddResult[32] | N703;
  assign N705 = io_mulAddResult[31] | N704;
  assign N706 = io_mulAddResult[30] | N705;
  assign N707 = io_mulAddResult[29] | N706;
  assign N708 = io_mulAddResult[28] | N707;
  assign N709 = io_mulAddResult[27] | N708;
  assign N710 = io_mulAddResult[26] | N709;
  assign N711 = io_mulAddResult[25] | N710;
  assign N712 = io_mulAddResult[24] | N711;
  assign N713 = io_mulAddResult[23] | N712;
  assign N714 = io_mulAddResult[22] | N713;
  assign N715 = io_mulAddResult[21] | N714;
  assign N716 = io_mulAddResult[20] | N715;
  assign N717 = io_mulAddResult[19] | N716;
  assign N718 = io_mulAddResult[18] | N717;
  assign N719 = io_mulAddResult[17] | N718;
  assign N720 = io_mulAddResult[16] | N719;
  assign N721 = io_mulAddResult[15] | N720;
  assign N722 = io_mulAddResult[14] | N721;
  assign N723 = io_mulAddResult[13] | N722;
  assign N724 = io_mulAddResult[12] | N723;
  assign N725 = io_mulAddResult[11] | N724;
  assign N726 = io_mulAddResult[10] | N725;
  assign N727 = io_mulAddResult[9] | N726;
  assign N728 = io_mulAddResult[8] | N727;
  assign N729 = io_mulAddResult[7] | N728;
  assign N730 = io_mulAddResult[6] | N729;
  assign N731 = io_mulAddResult[5] | N730;
  assign N732 = io_mulAddResult[4] | N731;
  assign N733 = io_mulAddResult[3] | N732;
  assign N734 = io_mulAddResult[2] | N733;
  assign N735 = io_mulAddResult[1] | N734;
  assign N736 = io_mulAddResult[0] | N735;
  assign N737 = io_fromPreMul_bit0AlignedNegSigC | N736;
  assign N738 = io_mulAddResult[73] | io_mulAddResult[74];
  assign N739 = io_mulAddResult[72] | N738;
  assign N740 = io_mulAddResult[71] | N739;
  assign N741 = io_mulAddResult[70] | N740;
  assign N742 = io_mulAddResult[69] | N741;
  assign N743 = io_mulAddResult[68] | N742;
  assign N744 = io_mulAddResult[67] | N743;
  assign N745 = io_mulAddResult[66] | N744;
  assign N746 = io_mulAddResult[65] | N745;
  assign N747 = io_mulAddResult[64] | N746;
  assign N748 = io_mulAddResult[63] | N747;
  assign N749 = io_mulAddResult[62] | N748;
  assign N750 = io_mulAddResult[61] | N749;
  assign N751 = io_mulAddResult[60] | N750;
  assign N752 = io_mulAddResult[59] | N751;
  assign N753 = io_mulAddResult[58] | N752;
  assign N754 = io_mulAddResult[57] | N753;
  assign N755 = io_mulAddResult[56] | N754;
  assign N756 = io_mulAddResult[55] | N755;
  assign N757 = io_mulAddResult[54] | N756;
  assign N758 = io_mulAddResult[53] | N757;
  assign N759 = io_mulAddResult[52] | N758;
  assign N760 = io_mulAddResult[51] | N759;
  assign N761 = io_mulAddResult[50] | N760;
  assign N762 = io_mulAddResult[49] | N761;
  assign N763 = io_mulAddResult[48] | N762;
  assign N764 = io_mulAddResult[47] | N763;
  assign N765 = io_mulAddResult[46] | N764;
  assign N766 = io_mulAddResult[45] | N765;
  assign N767 = io_mulAddResult[44] | N766;
  assign N768 = io_mulAddResult[43] | N767;
  assign N769 = T199[42] | T199[43];
  assign N770 = T199[41] | N769;
  assign N771 = T199[40] | N770;
  assign N772 = T199[39] | N771;
  assign N773 = T199[38] | N772;
  assign N774 = T199[37] | N773;
  assign N775 = T199[36] | N774;
  assign N776 = T199[35] | N775;
  assign N777 = T199[34] | N776;
  assign N778 = T199[33] | N777;
  assign N779 = T199[32] | N778;
  assign N780 = T199[31] | N779;
  assign N781 = T199[30] | N780;
  assign N782 = T199[29] | N781;
  assign N783 = T199[28] | N782;
  assign N784 = T199[27] | N783;
  assign N785 = T199[26] | N784;
  assign N786 = T199[25] | N785;
  assign N787 = T199[24] | N786;
  assign N788 = T199[23] | N787;
  assign N789 = T199[22] | N788;
  assign N790 = T199[21] | N789;
  assign N791 = T199[20] | N790;
  assign N792 = T199[19] | N791;
  assign N793 = T199[18] | N792;
  assign N794 = T199[17] | N793;
  assign N795 = T199[16] | N794;
  assign N796 = T199[15] | N795;
  assign N797 = T199[14] | N796;
  assign N798 = T199[13] | N797;
  assign N799 = T199[12] | N798;
  assign N800 = T199[11] | N799;
  assign N801 = T199[10] | N800;
  assign N802 = T199[9] | N801;
  assign N803 = T199[8] | N802;
  assign N804 = T199[7] | N803;
  assign N805 = T199[6] | N804;
  assign N806 = T199[5] | N805;
  assign N807 = T199[4] | N806;
  assign N808 = T199[3] | N807;
  assign N809 = T199[2] | N808;
  assign N810 = T199[1] | N809;
  assign N811 = T199[0] | N810;
  assign T31 = io_fromPreMul_highAlignedNegSigC + 1'b1;
  assign T663 = io_fromPreMul_CAlignDist[5:0] - 1'b1;
  assign { T182[53:53], T182_0 } = 1'b0 - T682[0];
  assign { T186[85:85], T186_0 } = 1'b0 - T682[0];
  assign { T213[21:21], T213_0 } = 1'b0 - T682[0];
  assign T20 = { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } - T448;
  assign { sExpX3[13:13], sExpX3_13 } = io_fromPreMul_sExpSum - T447;
  assign T306 = sExpX3_13 - 1'b1;
  assign T356 = sExpX3_13 + 1'b1;
  assign { T104[55:55], T104_0 } = 1'b0 - sExpX3[13];
  assign roundUp_sigY3 = T314 + 1'b1;
  assign { T385[51:51], T385_0 } = 1'b0 - T698[0];
  assign inexactY = (N0)? T287 : 
                    (N1)? anyRound : 1'b0;
  assign N0 = doIncrSig;
  assign N1 = N250;
  assign T447 = (N2)? CDom_estNormDist : 
                (N3)? T20 : 1'b0;
  assign N2 = io_fromPreMul_isCDominant;
  assign N3 = N369;
  assign T448 = (N4)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N5)? T450 : 1'b0;
  assign N4 = T22[107];
  assign N5 = N251;
  assign T450 = (N6)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N7)? T451 : 1'b0;
  assign N6 = T22[106];
  assign N7 = N252;
  assign T451 = (N8)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N9)? T452 : 1'b0;
  assign N8 = T22[105];
  assign N9 = N253;
  assign T452 = (N10)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N11)? T453 : 1'b0;
  assign N10 = T22[104];
  assign N11 = N254;
  assign T453 = (N12)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N13)? T454 : 1'b0;
  assign N12 = T22[103];
  assign N13 = N255;
  assign T454 = (N14)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N15)? T455 : 1'b0;
  assign N14 = T22[102];
  assign N15 = N256;
  assign T455 = (N16)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N17)? T456 : 1'b0;
  assign N16 = T22[101];
  assign N17 = N257;
  assign T456 = (N18)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N19)? T457 : 1'b0;
  assign N18 = T22[100];
  assign N19 = N258;
  assign T457 = (N20)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N21)? T458 : 1'b0;
  assign N20 = T22[99];
  assign N21 = N259;
  assign T458 = (N22)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N23)? T459 : 1'b0;
  assign N22 = T22[98];
  assign N23 = N260;
  assign T459 = (N24)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N25)? T460 : 1'b0;
  assign N24 = T22[97];
  assign N25 = N261;
  assign T460 = (N26)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N27)? T461 : 1'b0;
  assign N26 = T22[96];
  assign N27 = N262;
  assign T461 = (N28)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N29)? T462 : 1'b0;
  assign N28 = T22[95];
  assign N29 = N263;
  assign T462 = (N30)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N31)? T463 : 1'b0;
  assign N30 = T22[94];
  assign N31 = N264;
  assign T463 = (N32)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N33)? T464 : 1'b0;
  assign N32 = T22[93];
  assign N33 = N265;
  assign T464 = (N34)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N35)? T465 : 1'b0;
  assign N34 = T22[92];
  assign N35 = N266;
  assign T465 = (N36)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N37)? T466 : 1'b0;
  assign N36 = T22[91];
  assign N37 = N267;
  assign T466 = (N38)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N39)? T467 : 1'b0;
  assign N38 = T22[90];
  assign N39 = N268;
  assign T467 = (N40)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N41)? T468 : 1'b0;
  assign N40 = T22[89];
  assign N41 = N269;
  assign T468 = (N42)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N43)? T469 : 1'b0;
  assign N42 = T22[88];
  assign N43 = N270;
  assign T469 = (N44)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N45)? T470 : 1'b0;
  assign N44 = T22[87];
  assign N45 = N271;
  assign T470 = (N46)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N47)? T471 : 1'b0;
  assign N46 = T22[86];
  assign N47 = N272;
  assign T471 = (N48)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N49)? T472 : 1'b0;
  assign N48 = T22[85];
  assign N49 = N273;
  assign T472 = (N50)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N51)? T473 : 1'b0;
  assign N50 = T22[84];
  assign N51 = N274;
  assign T473 = (N52)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N53)? T474 : 1'b0;
  assign N52 = T22[83];
  assign N53 = N275;
  assign T474 = (N54)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N55)? T475 : 1'b0;
  assign N54 = T22[82];
  assign N55 = N276;
  assign T475 = (N56)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N57)? T476 : 1'b0;
  assign N56 = T22[81];
  assign N57 = N277;
  assign T476 = (N58)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N59)? T477 : 1'b0;
  assign N58 = T22[80];
  assign N59 = N278;
  assign T477 = (N60)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N61)? T478 : 1'b0;
  assign N60 = T22[79];
  assign N61 = N279;
  assign T478 = (N62)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N63)? T479 : 1'b0;
  assign N62 = T22[78];
  assign N63 = N280;
  assign T479 = (N64)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N65)? T480 : 1'b0;
  assign N64 = T22[77];
  assign N65 = N281;
  assign T480 = (N66)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N67)? T481 : 1'b0;
  assign N66 = T22[76];
  assign N67 = N282;
  assign T481 = (N68)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N69)? T482 : 1'b0;
  assign N68 = T22[75];
  assign N69 = N283;
  assign T482 = (N70)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N71)? T483 : 1'b0;
  assign N70 = T22[74];
  assign N71 = N284;
  assign T483 = (N72)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N73)? T484 : 1'b0;
  assign N72 = T22[73];
  assign N73 = N285;
  assign T484 = (N74)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N75)? T485 : 1'b0;
  assign N74 = T22[72];
  assign N75 = N286;
  assign T485 = (N76)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N77)? T486 : 1'b0;
  assign N76 = T22[71];
  assign N77 = N287;
  assign T486 = (N78)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N79)? T487 : 1'b0;
  assign N78 = T22[70];
  assign N79 = N288;
  assign T487 = (N80)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N81)? T488 : 1'b0;
  assign N80 = T22[69];
  assign N81 = N289;
  assign T488 = (N82)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N83)? T489 : 1'b0;
  assign N82 = T22[68];
  assign N83 = N290;
  assign T489 = (N84)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N85)? T490 : 1'b0;
  assign N84 = T22[67];
  assign N85 = N291;
  assign T490 = (N86)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N87)? T491 : 1'b0;
  assign N86 = T22[66];
  assign N87 = N292;
  assign T491 = (N88)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N89)? T492 : 1'b0;
  assign N88 = T22[65];
  assign N89 = N293;
  assign T492[5:0] = (N90)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N91)? T493 : 1'b0;
  assign N90 = T492[6];
  assign N91 = N294;
  assign T493 = (N92)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N93)? T494 : 1'b0;
  assign N92 = T22[63];
  assign N93 = N295;
  assign T494 = (N94)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N95)? T495 : 1'b0;
  assign N94 = T22[62];
  assign N95 = N296;
  assign T495 = (N96)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N97)? T496 : 1'b0;
  assign N96 = T22[61];
  assign N97 = N297;
  assign T496 = (N98)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N99)? T497 : 1'b0;
  assign N98 = T22[60];
  assign N99 = N298;
  assign T497 = (N100)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N101)? T498 : 1'b0;
  assign N100 = T22[59];
  assign N101 = N299;
  assign T498 = (N102)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N103)? T499 : 1'b0;
  assign N102 = T22[58];
  assign N103 = N300;
  assign T499 = (N104)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N105)? T500 : 1'b0;
  assign N104 = T22[57];
  assign N105 = N301;
  assign T500 = (N106)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N107)? T501 : 1'b0;
  assign N106 = T22[56];
  assign N107 = N302;
  assign T501 = (N108)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N109)? T502 : 1'b0;
  assign N108 = T22[55];
  assign N109 = N303;
  assign T502 = (N110)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N111)? T503 : 1'b0;
  assign N110 = T22[54];
  assign N111 = N304;
  assign T503 = (N112)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N113)? T504 : 1'b0;
  assign N112 = T22[53];
  assign N113 = N305;
  assign T504 = (N114)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N115)? T505 : 1'b0;
  assign N114 = T22[52];
  assign N115 = N306;
  assign T505 = (N116)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N117)? T506 : 1'b0;
  assign N116 = T22[51];
  assign N117 = N307;
  assign T506 = (N118)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N119)? T507 : 1'b0;
  assign N118 = T22[50];
  assign N119 = N308;
  assign T507 = (N120)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N121)? T508 : 1'b0;
  assign N120 = T22[49];
  assign N121 = N309;
  assign T508 = (N122)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N123)? T509 : 1'b0;
  assign N122 = T22[48];
  assign N123 = N310;
  assign T509 = (N124)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N125)? T510 : 1'b0;
  assign N124 = T22[47];
  assign N125 = N311;
  assign T510 = (N126)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N127)? T511 : 1'b0;
  assign N126 = T22[46];
  assign N127 = N312;
  assign T511 = (N128)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N129)? T512 : 1'b0;
  assign N128 = T22[45];
  assign N129 = N313;
  assign T512 = (N130)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N131)? T513 : 1'b0;
  assign N130 = T22[44];
  assign N131 = N314;
  assign T513 = (N132)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N133)? T514 : 1'b0;
  assign N132 = T22[43];
  assign N133 = N315;
  assign T514 = (N134)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N135)? T515 : 1'b0;
  assign N134 = T22[42];
  assign N135 = N316;
  assign T515 = (N136)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N137)? T516 : 1'b0;
  assign N136 = T22[41];
  assign N137 = N317;
  assign T516 = (N138)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N139)? T517 : 1'b0;
  assign N138 = T22[40];
  assign N139 = N318;
  assign T517 = (N140)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N141)? T518 : 1'b0;
  assign N140 = T22[39];
  assign N141 = N319;
  assign T518 = (N142)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N143)? T519 : 1'b0;
  assign N142 = T22[38];
  assign N143 = N320;
  assign T519 = (N144)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N145)? T520 : 1'b0;
  assign N144 = T22[37];
  assign N145 = N321;
  assign T520 = (N146)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N147)? T521 : 1'b0;
  assign N146 = T22[36];
  assign N147 = N322;
  assign T521 = (N148)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N149)? T522 : 1'b0;
  assign N148 = T22[35];
  assign N149 = N323;
  assign T522 = (N150)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N151)? T523 : 1'b0;
  assign N150 = T22[34];
  assign N151 = N324;
  assign T523 = (N152)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N153)? T524 : 1'b0;
  assign N152 = T22[33];
  assign N153 = N325;
  assign T524[4:0] = (N154)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N155)? T525 : 1'b0;
  assign N154 = T524[5];
  assign N155 = N326;
  assign T525 = (N156)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N157)? T526 : 1'b0;
  assign N156 = T22[31];
  assign N157 = N327;
  assign T526 = (N158)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N159)? T527 : 1'b0;
  assign N158 = T22[30];
  assign N159 = N328;
  assign T527 = (N160)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N161)? T528 : 1'b0;
  assign N160 = T22[29];
  assign N161 = N329;
  assign T528 = (N162)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N163)? T529 : 1'b0;
  assign N162 = T22[28];
  assign N163 = N330;
  assign T529 = (N164)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N165)? T530 : 1'b0;
  assign N164 = T22[27];
  assign N165 = N331;
  assign T530 = (N166)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N167)? T531 : 1'b0;
  assign N166 = T22[26];
  assign N167 = N332;
  assign T531 = (N168)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N169)? T532 : 1'b0;
  assign N168 = T22[25];
  assign N169 = N333;
  assign T532 = (N170)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N171)? T533 : 1'b0;
  assign N170 = T22[24];
  assign N171 = N334;
  assign T533 = (N172)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N173)? T534 : 1'b0;
  assign N172 = T22[23];
  assign N173 = N335;
  assign T534 = (N174)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N175)? T535 : 1'b0;
  assign N174 = T22[22];
  assign N175 = N336;
  assign T535 = (N176)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N177)? T536 : 1'b0;
  assign N176 = T22[21];
  assign N177 = N337;
  assign T536 = (N178)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N179)? T537 : 1'b0;
  assign N178 = T22[20];
  assign N179 = N338;
  assign T537 = (N180)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N181)? T538 : 1'b0;
  assign N180 = T22[19];
  assign N181 = N339;
  assign T538 = (N182)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N183)? T539 : 1'b0;
  assign N182 = T22[18];
  assign N183 = N340;
  assign T539 = (N184)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N185)? T540 : 1'b0;
  assign N184 = T22[17];
  assign N185 = N341;
  assign T540[3:0] = (N186)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N187)? T541 : 1'b0;
  assign N186 = T540[4];
  assign N187 = N342;
  assign T541 = (N188)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N189)? T542 : 1'b0;
  assign N188 = T22[15];
  assign N189 = N343;
  assign T542 = (N190)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N191)? T543 : 1'b0;
  assign N190 = T22[14];
  assign N191 = N344;
  assign T543 = (N192)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N193)? T544 : 1'b0;
  assign N192 = T22[13];
  assign N193 = N345;
  assign T544 = (N194)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N195)? T545 : 1'b0;
  assign N194 = T22[12];
  assign N195 = N346;
  assign T545 = (N196)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N197)? T546 : 1'b0;
  assign N196 = T22[11];
  assign N197 = N347;
  assign T546 = (N198)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N199)? T547 : 1'b0;
  assign N198 = T22[10];
  assign N199 = N348;
  assign T547 = (N200)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N201)? T548 : 1'b0;
  assign N200 = T22[9];
  assign N201 = N349;
  assign T548[2:0] = (N202)? { 1'b0, 1'b0, 1'b0 } : 
                     (N203)? T549 : 1'b0;
  assign N202 = T548[3];
  assign N203 = N350;
  assign T549 = (N204)? { 1'b1, 1'b1, 1'b1 } : 
                (N205)? T550 : 1'b0;
  assign N204 = T22[7];
  assign N205 = N351;
  assign T550 = (N206)? { 1'b1, 1'b1, 1'b0 } : 
                (N207)? T551 : 1'b0;
  assign N206 = T22[6];
  assign N207 = N352;
  assign T551 = (N208)? { 1'b1, 1'b0, 1'b1 } : 
                (N209)? T552 : 1'b0;
  assign N208 = T22[5];
  assign N209 = N353;
  assign T552[1:0] = (N210)? { 1'b0, 1'b0 } : 
                     (N211)? T553 : 1'b0;
  assign N210 = T552[2];
  assign N211 = N354;
  assign T553 = (N212)? { 1'b1, 1'b1 } : 
                (N213)? T554 : 1'b0;
  assign N212 = T22[3];
  assign N213 = N355;
  assign T554[0] = (N214)? 1'b0 : 
                   (N215)? T22[1] : 1'b0;
  assign N214 = T554[1];
  assign N215 = N356;
  assign { sigSum, T25 } = (N216)? T31 : 
                           (N217)? io_fromPreMul_highAlignedNegSigC : 1'b0;
  assign N216 = io_mulAddResult[106];
  assign N217 = N357;
  assign CDom_estNormDist = (N218)? io_fromPreMul_CAlignDist : 
                            (N219)? { 1'b0, 1'b0, T663 } : 1'b0;
  assign N218 = T36;
  assign N219 = N358;
  assign sigX3[0] = (N0)? N593 : 
                    (N1)? N624 : 1'b0;
  assign { cFirstNormAbsSigSum, T179 } = (N220)? T257 : 
                                         (N221)? { 1'b0, T681 } : 1'b0;
  assign N220 = sigSum[109];
  assign N221 = N359;
  assign T681 = (N2)? CDom_firstNormAbsSigSum : 
                (N3)? notCDom_pos_firstNormAbsSigSum : 1'b0;
  assign notCDom_pos_firstNormAbsSigSum = (N222)? T205 : 
                                          (N223)? T181 : 1'b0;
  assign N222 = T20[6];
  assign N223 = N360;
  assign T181 = (N224)? T185 : 
                (N225)? { io_mulAddResult[32:0], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182[53:53], T182_0 } : 1'b0;
  assign N224 = T20[5];
  assign N225 = N361;
  assign T185 = (N226)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T25, io_mulAddResult[105:43], T684[0:0] } : 
                (N227)? { io_mulAddResult[0:0], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186[85:85], T186_0 } : 1'b0;
  assign N226 = T20[4];
  assign N227 = N362;
  assign T684[0] = (N228)? T196 : 
                   (N229)? N737 : 1'b0;
  assign N228 = T682[0];
  assign N229 = N363;
  assign T205 = (N224)? { io_mulAddResult[64:0], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213[21:21], T213_0 } : 
                (N225)? { io_mulAddResult[96:11], T206[0:0] } : 1'b0;
  assign T206[0] = (N228)? N652 : 
                   (N229)? N662 : 1'b0;
  assign T257 = (N2)? { 1'b0, CDom_firstNormAbsSigSum } : 
                (N3)? notCDom_neg_cFirstNormAbsSigSum : 1'b0;
  assign notCDom_neg_cFirstNormAbsSigSum = (N222)? T269 : 
                                           (N223)? T258 : 1'b0;
  assign T258 = (N224)? { T261_87, T261_86, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T261 } : 
                (N225)? { T199[34:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { T261_87, T261_86, T261 } = (N226)? { 1'b0, 1'b0, notSigSum[107:44], N811 } : 
                                      (N227)? { T199[2:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T269 = (N224)? { notSigSum[66:44], T199[43:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N225)? { notSigSum[98:44], T199[43:12], N640 } : 1'b0;
  assign T305 = (N230)? T306 : 
                (N231)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N230 = N389;
  assign N231 = N388;
  assign T309 = (N232)? T310 : 
                (N233)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N232 = roundEven;
  assign N233 = N365;
  assign roundEven = (N0)? T319 : 
                     (N1)? T316 : 1'b0;
  assign T323 = (N234)? roundUp_sigY3 : 
                (N235)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N234 = T324;
  assign N235 = N366;
  assign roundDirectUp = (N236)? N627 : 
                         (N237)? N561 : 1'b0;
  assign N236 = signY;
  assign N237 = N367;
  assign signY = (N238)? N627 : 
                 (N239)? T327 : 1'b0;
  assign N238 = isZeroY;
  assign N239 = N368;
  assign doNegSignSum = (N2)? T328 : 
                        (N3)? sigSum[109] : 1'b0;
  assign T344 = (N240)? T345 : 
                (N241)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N240 = T348;
  assign N241 = N370;
  assign T353 = (N242)? sExpX3_13 : 
                (N243)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N242 = T308[0];
  assign N243 = N371;
  assign T355 = (N244)? T356 : 
                (N245)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N244 = T308[1];
  assign N245 = N372;
  assign T394 = (N246)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N247)? fractY : 1'b0;
  assign N246 = T397;
  assign N247 = N373;
  assign fractY = (N248)? sigY3[51:0] : 
                  (N249)? sigY3[52:1] : 1'b0;
  assign N248 = sigX3Shift1;
  assign N249 = N364;
  assign io_exceptionFlags[0] = io_exceptionFlags[2] | T3;
  assign T3 = commonCase & inexactY;
  assign N250 = ~doIncrSig;
  assign anyRound = N502 | N558;
  assign T4[56] = sigX3_56 & 1'b0;
  assign T4[55] = T446[0] & 1'b0;
  assign T4[54] = sigX3[54] & T445[54];
  assign T4[53] = sigX3[53] & T445[53];
  assign T4[52] = sigX3[52] & T445[52];
  assign T4[51] = sigX3[51] & T445[51];
  assign T4[50] = sigX3[50] & T445[50];
  assign T4[49] = sigX3[49] & T445[49];
  assign T4[48] = sigX3[48] & T445[48];
  assign T4[47] = sigX3[47] & T445[47];
  assign T4[46] = sigX3[46] & T445[46];
  assign T4[45] = sigX3[45] & T445[45];
  assign T4[44] = sigX3[44] & T445[44];
  assign T4[43] = sigX3[43] & T445[43];
  assign T4[42] = sigX3[42] & T445[42];
  assign T4[41] = sigX3[41] & T445[41];
  assign T4[40] = sigX3[40] & T445[40];
  assign T4[39] = sigX3[39] & T445[39];
  assign T4[38] = sigX3[38] & T445[38];
  assign T4[37] = sigX3[37] & T445[37];
  assign T4[36] = sigX3[36] & T445[36];
  assign T4[35] = sigX3[35] & T445[35];
  assign T4[34] = sigX3[34] & T445[34];
  assign T4[33] = sigX3[33] & T445[33];
  assign T4[32] = sigX3[32] & T445[32];
  assign T4[31] = sigX3[31] & T445[31];
  assign T4[30] = sigX3[30] & T445[30];
  assign T4[29] = sigX3[29] & T445[29];
  assign T4[28] = sigX3[28] & T445[28];
  assign T4[27] = sigX3[27] & T445[27];
  assign T4[26] = sigX3[26] & T445[26];
  assign T4[25] = sigX3[25] & T445[25];
  assign T4[24] = sigX3[24] & T445[24];
  assign T4[23] = sigX3[23] & T445[23];
  assign T4[22] = sigX3[22] & T445[22];
  assign T4[21] = sigX3[21] & T445[21];
  assign T4[20] = sigX3[20] & T445[20];
  assign T4[19] = sigX3[19] & T445[19];
  assign T4[18] = sigX3[18] & T445[18];
  assign T4[17] = sigX3[17] & T445[17];
  assign T4[16] = sigX3[16] & T445[16];
  assign T4[15] = sigX3[15] & T445[15];
  assign T4[14] = sigX3[14] & T445[14];
  assign T4[13] = sigX3[13] & T445[13];
  assign T4[12] = sigX3[12] & T445[12];
  assign T4[11] = sigX3[11] & T445[11];
  assign T4[10] = sigX3[10] & T445[10];
  assign T4[9] = sigX3[9] & T445[9];
  assign T4[8] = sigX3[8] & T445[8];
  assign T4[7] = sigX3[7] & T445[7];
  assign T4[6] = sigX3[6] & T445[6];
  assign T4[5] = sigX3[5] & T445[5];
  assign T4[4] = sigX3[4] & T445[4];
  assign T4[3] = sigX3[3] & T445[3];
  assign T4[2] = sigX3[2] & T445[2];
  assign T4[1] = sigX3[1] & T445[1];
  assign T4[0] = sigX3[0] & T445[0];
  assign T445[54] = T104[55] | T6[55];
  assign T445[53] = T104[55] | T6[54];
  assign T445[52] = T104[55] | T6[53];
  assign T445[51] = T104[55] | T6[52];
  assign T445[50] = T104[55] | T6[51];
  assign T445[49] = T104[55] | T6[50];
  assign T445[48] = T104[55] | T6[49];
  assign T445[47] = T104[55] | T6[48];
  assign T445[46] = T104[55] | T6[47];
  assign T445[45] = T104[55] | T6[46];
  assign T445[44] = T104[55] | T6[45];
  assign T445[43] = T104[55] | T6[44];
  assign T445[42] = T104[55] | T6[43];
  assign T445[41] = T104[55] | T6[42];
  assign T445[40] = T104[55] | T6[41];
  assign T445[39] = T104[55] | T6[40];
  assign T445[38] = T104[55] | T6[39];
  assign T445[37] = T104[55] | T6[38];
  assign T445[36] = T104[55] | T6[37];
  assign T445[35] = T104[55] | T6[36];
  assign T445[34] = T104[55] | T6[35];
  assign T445[33] = T104[55] | T6[34];
  assign T445[32] = T104[55] | T6[33];
  assign T445[31] = T104[55] | T6[32];
  assign T445[30] = T104[55] | T6[31];
  assign T445[29] = T104[55] | T6[30];
  assign T445[28] = T104[55] | T6[29];
  assign T445[27] = T104[55] | T6[28];
  assign T445[26] = T104[55] | T6[27];
  assign T445[25] = T104[55] | T6[26];
  assign T445[24] = T104[55] | T6[25];
  assign T445[23] = T104[55] | T6[24];
  assign T445[22] = T104[55] | T6[23];
  assign T445[21] = T104[55] | T6[22];
  assign T445[20] = T104[55] | T6[21];
  assign T445[19] = T104[55] | T6[20];
  assign T445[18] = T104[55] | T6[19];
  assign T445[17] = T104[55] | T6[18];
  assign T445[16] = T104[55] | T6[17];
  assign T445[15] = T104[55] | T6[16];
  assign T445[14] = T104[55] | T6[15];
  assign T445[13] = T104[55] | T6[14];
  assign T445[12] = T104[55] | T6[13];
  assign T445[11] = T104[55] | T6[12];
  assign T445[10] = T104[55] | T6[11];
  assign T445[9] = T104[55] | T6[10];
  assign T445[8] = T104[55] | T6[9];
  assign T445[7] = T104[55] | T6[8];
  assign T445[6] = T104[55] | T6[7];
  assign T445[5] = T104[55] | T6[6];
  assign T445[4] = T104[55] | T6[5];
  assign T445[3] = T104[55] | T6[4];
  assign T445[2] = T104[55] | T6[3];
  assign T445[1] = T104[55] | T6[2];
  assign T445[0] = T104[55] | 1'b1;
  assign roundMask[0] = T104_0 | 1'b1;
  assign T6[55] = T9[53] | 1'b0;
  assign T6[54] = T9[52] | 1'b0;
  assign T6[53] = T9[51] | 1'b0;
  assign T6[52] = T9[50] | 1'b0;
  assign T6[51] = T9[49] | 1'b0;
  assign T6[50] = T9[48] | 1'b0;
  assign T6[49] = T9[47] | 1'b0;
  assign T6[48] = T9[46] | 1'b0;
  assign T6[47] = T9[45] | 1'b0;
  assign T6[46] = T9[44] | 1'b0;
  assign T6[45] = T9[43] | 1'b0;
  assign T6[44] = T9[42] | 1'b0;
  assign T6[43] = T9[41] | 1'b0;
  assign T6[42] = T9[40] | 1'b0;
  assign T6[41] = T9[39] | 1'b0;
  assign T6[40] = T9[38] | 1'b0;
  assign T6[39] = T9[37] | 1'b0;
  assign T6[38] = T9[36] | 1'b0;
  assign T6[37] = T9[35] | 1'b0;
  assign T6[36] = T9[34] | 1'b0;
  assign T6[35] = T9[33] | 1'b0;
  assign T6[34] = T9[32] | 1'b0;
  assign T6[33] = T9[31] | 1'b0;
  assign T6[32] = T9[30] | 1'b0;
  assign T6[31] = T9[29] | 1'b0;
  assign T6[30] = T9[28] | 1'b0;
  assign T6[29] = T9[27] | 1'b0;
  assign T6[28] = T9[26] | 1'b0;
  assign T6[27] = T9[25] | 1'b0;
  assign T6[26] = T9[24] | 1'b0;
  assign T6[25] = T9[23] | 1'b0;
  assign T6[24] = T9[22] | 1'b0;
  assign T6[23] = T9[21] | 1'b0;
  assign T6[22] = T9[20] | 1'b0;
  assign T6[21] = T9[19] | 1'b0;
  assign T6[20] = T9[18] | 1'b0;
  assign T6[19] = T9[17] | 1'b0;
  assign T6[18] = T9[16] | 1'b0;
  assign T6[17] = T9[15] | 1'b0;
  assign T6[16] = T9[14] | 1'b0;
  assign T6[15] = T9[13] | 1'b0;
  assign T6[14] = T9[12] | 1'b0;
  assign T6[13] = T9[11] | 1'b0;
  assign T6[12] = T9[10] | 1'b0;
  assign T6[11] = T9[9] | 1'b0;
  assign T6[10] = T9[8] | 1'b0;
  assign T6[9] = T9[7] | 1'b0;
  assign T6[8] = T9[6] | 1'b0;
  assign T6[7] = T15[0] | 1'b0;
  assign T6[6] = T15[1] | 1'b0;
  assign T6[5] = T15[2] | 1'b0;
  assign T6[4] = T15[3] | 1'b0;
  assign T6[3] = T14[0] | 1'b0;
  assign T6[2] = T9_0 | T446[0];
  assign T19[12] = ~sExpX3_13[12];
  assign T19[11] = ~sExpX3_13[11];
  assign T19[10] = ~sExpX3_13[10];
  assign T19[9] = ~sExpX3_13[9];
  assign T19[8] = ~sExpX3_13[8];
  assign T19[7] = ~sExpX3_13[7];
  assign T19[6] = ~sExpX3_13[6];
  assign T19[5] = ~sExpX3_13[5];
  assign T19[4] = ~sExpX3_13[4];
  assign T19[3] = ~sExpX3_13[3];
  assign T19[2] = ~sExpX3_13[2];
  assign T19[1] = ~sExpX3_13[1];
  assign T19[0] = ~sExpX3_13[0];
  assign N251 = ~T22[107];
  assign N252 = ~T22[106];
  assign N253 = ~T22[105];
  assign N254 = ~T22[104];
  assign N255 = ~T22[103];
  assign N256 = ~T22[102];
  assign N257 = ~T22[101];
  assign N258 = ~T22[100];
  assign N259 = ~T22[99];
  assign N260 = ~T22[98];
  assign N261 = ~T22[97];
  assign N262 = ~T22[96];
  assign N263 = ~T22[95];
  assign N264 = ~T22[94];
  assign N265 = ~T22[93];
  assign N266 = ~T22[92];
  assign N267 = ~T22[91];
  assign N268 = ~T22[90];
  assign N269 = ~T22[89];
  assign N270 = ~T22[88];
  assign N271 = ~T22[87];
  assign N272 = ~T22[86];
  assign N273 = ~T22[85];
  assign N274 = ~T22[84];
  assign N275 = ~T22[83];
  assign N276 = ~T22[82];
  assign N277 = ~T22[81];
  assign N278 = ~T22[80];
  assign N279 = ~T22[79];
  assign N280 = ~T22[78];
  assign N281 = ~T22[77];
  assign N282 = ~T22[76];
  assign N283 = ~T22[75];
  assign N284 = ~T22[74];
  assign N285 = ~T22[73];
  assign N286 = ~T22[72];
  assign N287 = ~T22[71];
  assign N288 = ~T22[70];
  assign N289 = ~T22[69];
  assign N290 = ~T22[68];
  assign N291 = ~T22[67];
  assign N292 = ~T22[66];
  assign N293 = ~T22[65];
  assign N294 = ~T22[64];
  assign T492[6] = T22[64];
  assign N295 = ~T22[63];
  assign N296 = ~T22[62];
  assign N297 = ~T22[61];
  assign N298 = ~T22[60];
  assign N299 = ~T22[59];
  assign N300 = ~T22[58];
  assign N301 = ~T22[57];
  assign N302 = ~T22[56];
  assign N303 = ~T22[55];
  assign N304 = ~T22[54];
  assign N305 = ~T22[53];
  assign N306 = ~T22[52];
  assign N307 = ~T22[51];
  assign N308 = ~T22[50];
  assign N309 = ~T22[49];
  assign N310 = ~T22[48];
  assign N311 = ~T22[47];
  assign N312 = ~T22[46];
  assign N313 = ~T22[45];
  assign N314 = ~T22[44];
  assign N315 = ~T22[43];
  assign N316 = ~T22[42];
  assign N317 = ~T22[41];
  assign N318 = ~T22[40];
  assign N319 = ~T22[39];
  assign N320 = ~T22[38];
  assign N321 = ~T22[37];
  assign N322 = ~T22[36];
  assign N323 = ~T22[35];
  assign N324 = ~T22[34];
  assign N325 = ~T22[33];
  assign N326 = ~T22[32];
  assign T524[5] = T22[32];
  assign N327 = ~T22[31];
  assign N328 = ~T22[30];
  assign N329 = ~T22[29];
  assign N330 = ~T22[28];
  assign N331 = ~T22[27];
  assign N332 = ~T22[26];
  assign N333 = ~T22[25];
  assign N334 = ~T22[24];
  assign N335 = ~T22[23];
  assign N336 = ~T22[22];
  assign N337 = ~T22[21];
  assign N338 = ~T22[20];
  assign N339 = ~T22[19];
  assign N340 = ~T22[18];
  assign N341 = ~T22[17];
  assign N342 = ~T22[16];
  assign T540[4] = T22[16];
  assign N343 = ~T22[15];
  assign N344 = ~T22[14];
  assign N345 = ~T22[13];
  assign N346 = ~T22[12];
  assign N347 = ~T22[11];
  assign N348 = ~T22[10];
  assign N349 = ~T22[9];
  assign N350 = ~T22[8];
  assign T548[3] = T22[8];
  assign N351 = ~T22[7];
  assign N352 = ~T22[6];
  assign N353 = ~T22[5];
  assign N354 = ~T22[4];
  assign T552[2] = T22[4];
  assign N355 = ~T22[3];
  assign N356 = ~T22[2];
  assign T554[1] = T22[2];
  assign T22[107] = T25[108] ^ T25[107];
  assign T22[106] = T25[107] ^ io_mulAddResult[105];
  assign T22[105] = io_mulAddResult[105] ^ io_mulAddResult[104];
  assign T22[104] = io_mulAddResult[104] ^ io_mulAddResult[103];
  assign T22[103] = io_mulAddResult[103] ^ io_mulAddResult[102];
  assign T22[102] = io_mulAddResult[102] ^ io_mulAddResult[101];
  assign T22[101] = io_mulAddResult[101] ^ io_mulAddResult[100];
  assign T22[100] = io_mulAddResult[100] ^ io_mulAddResult[99];
  assign T22[99] = io_mulAddResult[99] ^ io_mulAddResult[98];
  assign T22[98] = io_mulAddResult[98] ^ io_mulAddResult[97];
  assign T22[97] = io_mulAddResult[97] ^ io_mulAddResult[96];
  assign T22[96] = io_mulAddResult[96] ^ io_mulAddResult[95];
  assign T22[95] = io_mulAddResult[95] ^ io_mulAddResult[94];
  assign T22[94] = io_mulAddResult[94] ^ io_mulAddResult[93];
  assign T22[93] = io_mulAddResult[93] ^ io_mulAddResult[92];
  assign T22[92] = io_mulAddResult[92] ^ io_mulAddResult[91];
  assign T22[91] = io_mulAddResult[91] ^ io_mulAddResult[90];
  assign T22[90] = io_mulAddResult[90] ^ io_mulAddResult[89];
  assign T22[89] = io_mulAddResult[89] ^ io_mulAddResult[88];
  assign T22[88] = io_mulAddResult[88] ^ io_mulAddResult[87];
  assign T22[87] = io_mulAddResult[87] ^ io_mulAddResult[86];
  assign T22[86] = io_mulAddResult[86] ^ io_mulAddResult[85];
  assign T22[85] = io_mulAddResult[85] ^ io_mulAddResult[84];
  assign T22[84] = io_mulAddResult[84] ^ io_mulAddResult[83];
  assign T22[83] = io_mulAddResult[83] ^ io_mulAddResult[82];
  assign T22[82] = io_mulAddResult[82] ^ io_mulAddResult[81];
  assign T22[81] = io_mulAddResult[81] ^ io_mulAddResult[80];
  assign T22[80] = io_mulAddResult[80] ^ io_mulAddResult[79];
  assign T22[79] = io_mulAddResult[79] ^ io_mulAddResult[78];
  assign T22[78] = io_mulAddResult[78] ^ io_mulAddResult[77];
  assign T22[77] = io_mulAddResult[77] ^ io_mulAddResult[76];
  assign T22[76] = io_mulAddResult[76] ^ io_mulAddResult[75];
  assign T22[75] = io_mulAddResult[75] ^ io_mulAddResult[74];
  assign T22[74] = io_mulAddResult[74] ^ io_mulAddResult[73];
  assign T22[73] = io_mulAddResult[73] ^ io_mulAddResult[72];
  assign T22[72] = io_mulAddResult[72] ^ io_mulAddResult[71];
  assign T22[71] = io_mulAddResult[71] ^ io_mulAddResult[70];
  assign T22[70] = io_mulAddResult[70] ^ io_mulAddResult[69];
  assign T22[69] = io_mulAddResult[69] ^ io_mulAddResult[68];
  assign T22[68] = io_mulAddResult[68] ^ io_mulAddResult[67];
  assign T22[67] = io_mulAddResult[67] ^ io_mulAddResult[66];
  assign T22[66] = io_mulAddResult[66] ^ io_mulAddResult[65];
  assign T22[65] = io_mulAddResult[65] ^ io_mulAddResult[64];
  assign T22[64] = io_mulAddResult[64] ^ io_mulAddResult[63];
  assign T22[63] = io_mulAddResult[63] ^ io_mulAddResult[62];
  assign T22[62] = io_mulAddResult[62] ^ io_mulAddResult[61];
  assign T22[61] = io_mulAddResult[61] ^ io_mulAddResult[60];
  assign T22[60] = io_mulAddResult[60] ^ io_mulAddResult[59];
  assign T22[59] = io_mulAddResult[59] ^ io_mulAddResult[58];
  assign T22[58] = io_mulAddResult[58] ^ io_mulAddResult[57];
  assign T22[57] = io_mulAddResult[57] ^ io_mulAddResult[56];
  assign T22[56] = io_mulAddResult[56] ^ io_mulAddResult[55];
  assign T22[55] = io_mulAddResult[55] ^ io_mulAddResult[54];
  assign T22[54] = io_mulAddResult[54] ^ io_mulAddResult[53];
  assign T22[53] = io_mulAddResult[53] ^ io_mulAddResult[52];
  assign T22[52] = io_mulAddResult[52] ^ io_mulAddResult[51];
  assign T22[51] = io_mulAddResult[51] ^ io_mulAddResult[50];
  assign T22[50] = io_mulAddResult[50] ^ io_mulAddResult[49];
  assign T22[49] = io_mulAddResult[49] ^ io_mulAddResult[48];
  assign T22[48] = io_mulAddResult[48] ^ io_mulAddResult[47];
  assign T22[47] = io_mulAddResult[47] ^ io_mulAddResult[46];
  assign T22[46] = io_mulAddResult[46] ^ io_mulAddResult[45];
  assign T22[45] = io_mulAddResult[45] ^ io_mulAddResult[44];
  assign T22[44] = io_mulAddResult[44] ^ io_mulAddResult[43];
  assign T22[43] = io_mulAddResult[43] ^ io_mulAddResult[42];
  assign T22[42] = io_mulAddResult[42] ^ io_mulAddResult[41];
  assign T22[41] = io_mulAddResult[41] ^ io_mulAddResult[40];
  assign T22[40] = io_mulAddResult[40] ^ io_mulAddResult[39];
  assign T22[39] = io_mulAddResult[39] ^ io_mulAddResult[38];
  assign T22[38] = io_mulAddResult[38] ^ io_mulAddResult[37];
  assign T22[37] = io_mulAddResult[37] ^ io_mulAddResult[36];
  assign T22[36] = io_mulAddResult[36] ^ io_mulAddResult[35];
  assign T22[35] = io_mulAddResult[35] ^ io_mulAddResult[34];
  assign T22[34] = io_mulAddResult[34] ^ io_mulAddResult[33];
  assign T22[33] = io_mulAddResult[33] ^ io_mulAddResult[32];
  assign T22[32] = io_mulAddResult[32] ^ io_mulAddResult[31];
  assign T22[31] = io_mulAddResult[31] ^ io_mulAddResult[30];
  assign T22[30] = io_mulAddResult[30] ^ io_mulAddResult[29];
  assign T22[29] = io_mulAddResult[29] ^ io_mulAddResult[28];
  assign T22[28] = io_mulAddResult[28] ^ io_mulAddResult[27];
  assign T22[27] = io_mulAddResult[27] ^ io_mulAddResult[26];
  assign T22[26] = io_mulAddResult[26] ^ io_mulAddResult[25];
  assign T22[25] = io_mulAddResult[25] ^ io_mulAddResult[24];
  assign T22[24] = io_mulAddResult[24] ^ io_mulAddResult[23];
  assign T22[23] = io_mulAddResult[23] ^ io_mulAddResult[22];
  assign T22[22] = io_mulAddResult[22] ^ io_mulAddResult[21];
  assign T22[21] = io_mulAddResult[21] ^ io_mulAddResult[20];
  assign T22[20] = io_mulAddResult[20] ^ io_mulAddResult[19];
  assign T22[19] = io_mulAddResult[19] ^ io_mulAddResult[18];
  assign T22[18] = io_mulAddResult[18] ^ io_mulAddResult[17];
  assign T22[17] = io_mulAddResult[17] ^ io_mulAddResult[16];
  assign T22[16] = io_mulAddResult[16] ^ io_mulAddResult[15];
  assign T22[15] = io_mulAddResult[15] ^ io_mulAddResult[14];
  assign T22[14] = io_mulAddResult[14] ^ io_mulAddResult[13];
  assign T22[13] = io_mulAddResult[13] ^ io_mulAddResult[12];
  assign T22[12] = io_mulAddResult[12] ^ io_mulAddResult[11];
  assign T22[11] = io_mulAddResult[11] ^ io_mulAddResult[10];
  assign T22[10] = io_mulAddResult[10] ^ io_mulAddResult[9];
  assign T22[9] = io_mulAddResult[9] ^ io_mulAddResult[8];
  assign T22[8] = io_mulAddResult[8] ^ io_mulAddResult[7];
  assign T22[7] = io_mulAddResult[7] ^ io_mulAddResult[6];
  assign T22[6] = io_mulAddResult[6] ^ io_mulAddResult[5];
  assign T22[5] = io_mulAddResult[5] ^ io_mulAddResult[4];
  assign T22[4] = io_mulAddResult[4] ^ io_mulAddResult[3];
  assign T22[3] = io_mulAddResult[3] ^ io_mulAddResult[2];
  assign T22[2] = io_mulAddResult[2] ^ io_mulAddResult[1];
  assign T22[1] = io_mulAddResult[1] ^ io_mulAddResult[0];
  assign N357 = ~io_mulAddResult[106];
  assign N358 = ~T36;
  assign T36 = io_fromPreMul_CAlignDist_0 | T682[0];
  assign T682[0] = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T9[21] = 1'b0 | T49[15];
  assign T9[20] = T52[15] | 1'b0;
  assign T9[19] = 1'b0 | T49_13;
  assign T9[18] = T50[14] | 1'b0;
  assign T9[17] = 1'b0 | T49_11;
  assign T9[16] = T50_12 | 1'b0;
  assign T9[15] = 1'b0 | T49_9;
  assign T9[14] = T50_10 | 1'b0;
  assign T9[13] = 1'b0 | T49_7;
  assign T9[12] = T50_8 | 1'b0;
  assign T9[11] = 1'b0 | T49_5;
  assign T9[10] = T50_6 | 1'b0;
  assign T9[9] = 1'b0 | T49_3;
  assign T9[8] = T50_4 | 1'b0;
  assign T9[7] = 1'b0 | T49_1;
  assign T9[6] = T50_2 | 1'b0;
  assign T52[15] = 1'b0 | T53[15];
  assign T49[15] = 1'b0 | T53[14];
  assign T50[14] = T56[15] | 1'b0;
  assign T49_13 = T56[14] | 1'b0;
  assign T50_12 = 1'b0 | T53_11;
  assign T49_11 = 1'b0 | T53_10;
  assign T50_10 = T54[13] | 1'b0;
  assign T49_9 = T54[12] | 1'b0;
  assign T50_8 = 1'b0 | T53_7;
  assign T49_7 = 1'b0 | T53_6;
  assign T50_6 = T54_9 | 1'b0;
  assign T49_5 = T54_8 | 1'b0;
  assign T50_4 = 1'b0 | T53_3;
  assign T49_3 = 1'b0 | T53_2;
  assign T50_2 = T54_5 | 1'b0;
  assign T49_1 = T54_4 | 1'b0;
  assign T56[15] = 1'b0 | T57[15];
  assign T56[14] = 1'b0 | T57[14];
  assign T53[15] = 1'b0 | T57[13];
  assign T53[14] = 1'b0 | T57[12];
  assign T54[13] = T60[15] | 1'b0;
  assign T54[12] = T60[14] | 1'b0;
  assign T53_11 = T60[13] | 1'b0;
  assign T53_10 = T60[12] | 1'b0;
  assign T54_9 = 1'b0 | T57_7;
  assign T54_8 = 1'b0 | T57_6;
  assign T53_7 = 1'b0 | T57_5;
  assign T53_6 = 1'b0 | T57_4;
  assign T54_5 = T58[11] | 1'b0;
  assign T54_4 = T58[10] | 1'b0;
  assign T53_3 = T58[9] | 1'b0;
  assign T53_2 = T58[8] | 1'b0;
  assign T60[15] = 1'b0 | T16[7];
  assign T60[14] = 1'b0 | T16[6];
  assign T60[13] = 1'b0 | T16[5];
  assign T60[12] = 1'b0 | T16[4];
  assign T57[15] = 1'b0 | T16[3];
  assign T57[14] = 1'b0 | T16[2];
  assign T57[13] = 1'b0 | T16[1];
  assign T57[12] = 1'b0 | T16[0];
  assign T58[11] = T16[15] | 1'b0;
  assign T58[10] = T16[14] | 1'b0;
  assign T58[9] = T16[13] | 1'b0;
  assign T58[8] = T16[12] | 1'b0;
  assign T57_7 = T16[11] | 1'b0;
  assign T57_6 = T16[10] | 1'b0;
  assign T57_5 = T16[9] | 1'b0;
  assign T57_4 = T16[8] | 1'b0;
  assign T9[53] = 1'b0 | T74[31];
  assign T9[52] = T77[31] | 1'b0;
  assign T9[51] = 1'b0 | T74_29;
  assign T9[50] = T75[30] | 1'b0;
  assign T9[49] = 1'b0 | T74_27;
  assign T9[48] = T75_28 | 1'b0;
  assign T9[47] = 1'b0 | T74_25;
  assign T9[46] = T75_26 | 1'b0;
  assign T9[45] = 1'b0 | T74_23;
  assign T9[44] = T75_24 | 1'b0;
  assign T9[43] = 1'b0 | T74_21;
  assign T9[42] = T75_22 | 1'b0;
  assign T9[41] = 1'b0 | T74_19;
  assign T9[40] = T75_20 | 1'b0;
  assign T9[39] = 1'b0 | T74_17;
  assign T9[38] = T75_18 | 1'b0;
  assign T9[37] = 1'b0 | T74_15;
  assign T9[36] = T75_16 | 1'b0;
  assign T9[35] = 1'b0 | T74_13;
  assign T9[34] = T75_14 | 1'b0;
  assign T9[33] = 1'b0 | T74_11;
  assign T9[32] = T75_12 | 1'b0;
  assign T9[31] = 1'b0 | T74_9;
  assign T9[30] = T75_10 | 1'b0;
  assign T9[29] = 1'b0 | T74_7;
  assign T9[28] = T75_8 | 1'b0;
  assign T9[27] = 1'b0 | T74_5;
  assign T9[26] = T75_6 | 1'b0;
  assign T9[25] = 1'b0 | T74_3;
  assign T9[24] = T75_4 | 1'b0;
  assign T9[23] = 1'b0 | T74_1;
  assign T9[22] = T75_2 | 1'b0;
  assign T77[31] = 1'b0 | T78[31];
  assign T74[31] = 1'b0 | T78[30];
  assign T75[30] = T81[31] | 1'b0;
  assign T74_29 = T81[30] | 1'b0;
  assign T75_28 = 1'b0 | T78_27;
  assign T74_27 = 1'b0 | T78_26;
  assign T75_26 = T79[29] | 1'b0;
  assign T74_25 = T79[28] | 1'b0;
  assign T75_24 = 1'b0 | T78_23;
  assign T74_23 = 1'b0 | T78_22;
  assign T75_22 = T79_25 | 1'b0;
  assign T74_21 = T79_24 | 1'b0;
  assign T75_20 = 1'b0 | T78_19;
  assign T74_19 = 1'b0 | T78_18;
  assign T75_18 = T79_21 | 1'b0;
  assign T74_17 = T79_20 | 1'b0;
  assign T75_16 = 1'b0 | T78_15;
  assign T74_15 = 1'b0 | T78_14;
  assign T75_14 = T79_17 | 1'b0;
  assign T74_13 = T79_16 | 1'b0;
  assign T75_12 = 1'b0 | T78_11;
  assign T74_11 = 1'b0 | T78_10;
  assign T75_10 = T79_13 | 1'b0;
  assign T74_9 = T79_12 | 1'b0;
  assign T75_8 = 1'b0 | T78_7;
  assign T74_7 = 1'b0 | T78_6;
  assign T75_6 = T79_9 | 1'b0;
  assign T74_5 = T79_8 | 1'b0;
  assign T75_4 = 1'b0 | T78_3;
  assign T74_3 = 1'b0 | T78_2;
  assign T75_2 = T79_5 | 1'b0;
  assign T74_1 = T79_4 | 1'b0;
  assign T81[31] = 1'b0 | T82[31];
  assign T81[30] = 1'b0 | T82[30];
  assign T78[31] = 1'b0 | T82[29];
  assign T78[30] = 1'b0 | T82[28];
  assign T79[29] = T85[31] | 1'b0;
  assign T79[28] = T85[30] | 1'b0;
  assign T78_27 = T85[29] | 1'b0;
  assign T78_26 = T85[28] | 1'b0;
  assign T79_25 = 1'b0 | T82_23;
  assign T79_24 = 1'b0 | T82_22;
  assign T78_23 = 1'b0 | T82_21;
  assign T78_22 = 1'b0 | T82_20;
  assign T79_21 = T83[27] | 1'b0;
  assign T79_20 = T83[26] | 1'b0;
  assign T78_19 = T83[25] | 1'b0;
  assign T78_18 = T83[24] | 1'b0;
  assign T79_17 = 1'b0 | T82_15;
  assign T79_16 = 1'b0 | T82_14;
  assign T78_15 = 1'b0 | T82_13;
  assign T78_14 = 1'b0 | T82_12;
  assign T79_13 = T83_19 | 1'b0;
  assign T79_12 = T83_18 | 1'b0;
  assign T78_11 = T83_17 | 1'b0;
  assign T78_10 = T83_16 | 1'b0;
  assign T79_9 = 1'b0 | T82_7;
  assign T79_8 = 1'b0 | T82_6;
  assign T78_7 = 1'b0 | T82_5;
  assign T78_6 = 1'b0 | T82_4;
  assign T79_5 = T83_11 | 1'b0;
  assign T79_4 = T83_10 | 1'b0;
  assign T78_3 = T83_9 | 1'b0;
  assign T78_2 = T83_8 | 1'b0;
  assign T85[31] = 1'b0 | T86[31];
  assign T85[30] = 1'b0 | T86[30];
  assign T85[29] = 1'b0 | T86[29];
  assign T85[28] = 1'b0 | T86[28];
  assign T82[31] = 1'b0 | T86[27];
  assign T82[30] = 1'b0 | T86[26];
  assign T82[29] = 1'b0 | T86[25];
  assign T82[28] = 1'b0 | T86[24];
  assign T83[27] = T89[31] | 1'b0;
  assign T83[26] = T89[30] | 1'b0;
  assign T83[25] = T89[29] | 1'b0;
  assign T83[24] = T89[28] | 1'b0;
  assign T82_23 = T89[27] | 1'b0;
  assign T82_22 = T89[26] | 1'b0;
  assign T82_21 = T89[25] | 1'b0;
  assign T82_20 = T89[24] | 1'b0;
  assign T83_19 = 1'b0 | T86_15;
  assign T83_18 = 1'b0 | T86_14;
  assign T83_17 = 1'b0 | T86_13;
  assign T83_16 = 1'b0 | T86_12;
  assign T82_15 = 1'b0 | T86_11;
  assign T82_14 = 1'b0 | T86_10;
  assign T82_13 = 1'b0 | T86_9;
  assign T82_12 = 1'b0 | T86_8;
  assign T83_11 = T87[23] | 1'b0;
  assign T83_10 = T87[22] | 1'b0;
  assign T83_9 = T87[21] | 1'b0;
  assign T83_8 = T87[20] | 1'b0;
  assign T82_7 = T87[19] | 1'b0;
  assign T82_6 = T87[18] | 1'b0;
  assign T82_5 = T87[17] | 1'b0;
  assign T82_4 = T87[16] | 1'b0;
  assign T89[31] = 1'b0 | T17[15];
  assign T89[30] = 1'b0 | T17[14];
  assign T89[29] = 1'b0 | T17[13];
  assign T89[28] = 1'b0 | T17[12];
  assign T89[27] = 1'b0 | T17[11];
  assign T89[26] = 1'b0 | T17[10];
  assign T89[25] = 1'b0 | T17[9];
  assign T89[24] = 1'b0 | T17[8];
  assign T86[31] = 1'b0 | T17[7];
  assign T86[30] = 1'b0 | T17[6];
  assign T86[29] = 1'b0 | T17[5];
  assign T86[28] = 1'b0 | T17[4];
  assign T86[27] = 1'b0 | T17[3];
  assign T86[26] = 1'b0 | T17[2];
  assign T86[25] = 1'b0 | T17[1];
  assign T86[24] = 1'b0 | T17[0];
  assign T87[23] = T17[31] | 1'b0;
  assign T87[22] = T17[30] | 1'b0;
  assign T87[21] = T17[29] | 1'b0;
  assign T87[20] = T17[28] | 1'b0;
  assign T87[19] = T17[27] | 1'b0;
  assign T87[18] = T17[26] | 1'b0;
  assign T87[17] = T17[25] | 1'b0;
  assign T87[16] = T17[24] | 1'b0;
  assign T86_15 = T17[23] | 1'b0;
  assign T86_14 = T17[22] | 1'b0;
  assign T86_13 = T17[21] | 1'b0;
  assign T86_12 = T17[20] | 1'b0;
  assign T86_11 = T17[19] | 1'b0;
  assign T86_10 = T17[18] | 1'b0;
  assign T86_9 = T17[17] | 1'b0;
  assign T86_8 = T17[16] | 1'b0;
  assign T109[31] = T179[31] & absSigSumExtraMask[31];
  assign T109[30] = T179[30] & absSigSumExtraMask[30];
  assign T109[29] = T179[29] & absSigSumExtraMask[29];
  assign T109[28] = T179[28] & absSigSumExtraMask[28];
  assign T109[27] = T179[27] & absSigSumExtraMask[27];
  assign T109[26] = T179[26] & absSigSumExtraMask[26];
  assign T109[25] = T179[25] & absSigSumExtraMask[25];
  assign T109[24] = T179[24] & absSigSumExtraMask[24];
  assign T109[23] = T179[23] & absSigSumExtraMask[23];
  assign T109[22] = T179[22] & absSigSumExtraMask[22];
  assign T109[21] = T179[21] & absSigSumExtraMask[21];
  assign T109[20] = T179[20] & absSigSumExtraMask[20];
  assign T109[19] = T179[19] & absSigSumExtraMask[19];
  assign T109[18] = T179[18] & absSigSumExtraMask[18];
  assign T109[17] = T179[17] & absSigSumExtraMask[17];
  assign T109[16] = T179[16] & absSigSumExtraMask[16];
  assign T109[15] = T179[15] & absSigSumExtraMask[15];
  assign T109[14] = T179[14] & absSigSumExtraMask[14];
  assign T109[13] = T179[13] & absSigSumExtraMask[13];
  assign T109[12] = T179[12] & absSigSumExtraMask[12];
  assign T109[11] = T179[11] & absSigSumExtraMask[11];
  assign T109[10] = T179[10] & absSigSumExtraMask[10];
  assign T109[9] = T179[9] & absSigSumExtraMask[9];
  assign T109[8] = T179[8] & absSigSumExtraMask[8];
  assign T109[7] = T179[7] & T116[0];
  assign T109[6] = T179[6] & T116[1];
  assign T109[5] = T179[5] & T116[2];
  assign T109[4] = T179[4] & T116[3];
  assign T109[3] = T179[3] & T115[0];
  assign T109[2] = T179[2] & T115[1];
  assign T109[1] = T179[1] & absSigSumExtraMask_1;
  assign T109[0] = T179[0] & 1'b1;
  assign normTo2ShiftDist[4] = ~T447[4];
  assign normTo2ShiftDist[3] = ~T447[3];
  assign normTo2ShiftDist[2] = ~T447[2];
  assign normTo2ShiftDist[1] = ~T447[1];
  assign normTo2ShiftDist[0] = ~T447[0];
  assign absSigSumExtraMask[15] = 1'b0 | T136[7];
  assign absSigSumExtraMask[14] = T139[7] | 1'b0;
  assign absSigSumExtraMask[13] = 1'b0 | T136_5;
  assign absSigSumExtraMask[12] = T137[6] | 1'b0;
  assign absSigSumExtraMask[11] = 1'b0 | T136_3;
  assign absSigSumExtraMask[10] = T137_4 | 1'b0;
  assign absSigSumExtraMask[9] = 1'b0 | T136_1;
  assign absSigSumExtraMask[8] = T137_2 | 1'b0;
  assign T139[7] = 1'b0 | T140[7];
  assign T136[7] = 1'b0 | T140[6];
  assign T137[6] = T143[7] | 1'b0;
  assign T136_5 = T143[6] | 1'b0;
  assign T137_4 = 1'b0 | T140_3;
  assign T136_3 = 1'b0 | T140_2;
  assign T137_2 = T141[5] | 1'b0;
  assign T136_1 = T141[4] | 1'b0;
  assign T143[7] = 1'b0 | T117[3];
  assign T143[6] = 1'b0 | T117[2];
  assign T140[7] = 1'b0 | T117[1];
  assign T140[6] = 1'b0 | T117[0];
  assign T141[5] = T117[7] | 1'b0;
  assign T141[4] = T117[6] | 1'b0;
  assign T140_3 = T117[5] | 1'b0;
  assign T140_2 = T117[4] | 1'b0;
  assign absSigSumExtraMask[31] = 1'b0 | T155[15];
  assign absSigSumExtraMask[30] = T158[15] | 1'b0;
  assign absSigSumExtraMask[29] = 1'b0 | T155_13;
  assign absSigSumExtraMask[28] = T156[14] | 1'b0;
  assign absSigSumExtraMask[27] = 1'b0 | T155_11;
  assign absSigSumExtraMask[26] = T156_12 | 1'b0;
  assign absSigSumExtraMask[25] = 1'b0 | T155_9;
  assign absSigSumExtraMask[24] = T156_10 | 1'b0;
  assign absSigSumExtraMask[23] = 1'b0 | T155_7;
  assign absSigSumExtraMask[22] = T156_8 | 1'b0;
  assign absSigSumExtraMask[21] = 1'b0 | T155_5;
  assign absSigSumExtraMask[20] = T156_6 | 1'b0;
  assign absSigSumExtraMask[19] = 1'b0 | T155_3;
  assign absSigSumExtraMask[18] = T156_4 | 1'b0;
  assign absSigSumExtraMask[17] = 1'b0 | T155_1;
  assign absSigSumExtraMask[16] = T156_2 | 1'b0;
  assign T158[15] = 1'b0 | T159[15];
  assign T155[15] = 1'b0 | T159[14];
  assign T156[14] = T162[15] | 1'b0;
  assign T155_13 = T162[14] | 1'b0;
  assign T156_12 = 1'b0 | T159_11;
  assign T155_11 = 1'b0 | T159_10;
  assign T156_10 = T160[13] | 1'b0;
  assign T155_9 = T160[12] | 1'b0;
  assign T156_8 = 1'b0 | T159_7;
  assign T155_7 = 1'b0 | T159_6;
  assign T156_6 = T160_9 | 1'b0;
  assign T155_5 = T160_8 | 1'b0;
  assign T156_4 = 1'b0 | T159_3;
  assign T155_3 = 1'b0 | T159_2;
  assign T156_2 = T160_5 | 1'b0;
  assign T155_1 = T160_4 | 1'b0;
  assign T162[15] = 1'b0 | T163[15];
  assign T162[14] = 1'b0 | T163[14];
  assign T159[15] = 1'b0 | T163[13];
  assign T159[14] = 1'b0 | T163[12];
  assign T160[13] = T166[15] | 1'b0;
  assign T160[12] = T166[14] | 1'b0;
  assign T159_11 = T166[13] | 1'b0;
  assign T159_10 = T166[12] | 1'b0;
  assign T160_9 = 1'b0 | T163_7;
  assign T160_8 = 1'b0 | T163_6;
  assign T159_7 = 1'b0 | T163_5;
  assign T159_6 = 1'b0 | T163_4;
  assign T160_5 = T164[11] | 1'b0;
  assign T160_4 = T164[10] | 1'b0;
  assign T159_3 = T164[9] | 1'b0;
  assign T159_2 = T164[8] | 1'b0;
  assign T166[15] = 1'b0 | T118[7];
  assign T166[14] = 1'b0 | T118[6];
  assign T166[13] = 1'b0 | T118[5];
  assign T166[12] = 1'b0 | T118[4];
  assign T163[15] = 1'b0 | T118[3];
  assign T163[14] = 1'b0 | T118[2];
  assign T163[13] = 1'b0 | T118[1];
  assign T163[12] = 1'b0 | T118[0];
  assign T164[11] = T118[15] | 1'b0;
  assign T164[10] = T118[14] | 1'b0;
  assign T164[9] = T118[13] | 1'b0;
  assign T164[8] = T118[12] | 1'b0;
  assign T163_7 = T118[11] | 1'b0;
  assign T163_6 = T118[10] | 1'b0;
  assign T163_5 = T118[9] | 1'b0;
  assign T163_4 = T118[8] | 1'b0;
  assign N359 = ~sigSum[109];
  assign N360 = ~T20[6];
  assign N361 = ~T20[5];
  assign N362 = ~T20[4];
  assign N363 = ~T682[0];
  assign T196 = ~N811;
  assign notSigSum[161] = ~sigSum[161];
  assign notSigSum[160] = ~sigSum[160];
  assign notSigSum[159] = ~sigSum[159];
  assign notSigSum[158] = ~sigSum[158];
  assign notSigSum[157] = ~sigSum[157];
  assign notSigSum[156] = ~sigSum[156];
  assign notSigSum[155] = ~sigSum[155];
  assign notSigSum[154] = ~sigSum[154];
  assign notSigSum[153] = ~sigSum[153];
  assign notSigSum[152] = ~sigSum[152];
  assign notSigSum[151] = ~sigSum[151];
  assign notSigSum[150] = ~sigSum[150];
  assign notSigSum[149] = ~sigSum[149];
  assign notSigSum[148] = ~sigSum[148];
  assign notSigSum[147] = ~sigSum[147];
  assign notSigSum[146] = ~sigSum[146];
  assign notSigSum[145] = ~sigSum[145];
  assign notSigSum[144] = ~sigSum[144];
  assign notSigSum[143] = ~sigSum[143];
  assign notSigSum[142] = ~sigSum[142];
  assign notSigSum[141] = ~sigSum[141];
  assign notSigSum[140] = ~sigSum[140];
  assign notSigSum[139] = ~sigSum[139];
  assign notSigSum[138] = ~sigSum[138];
  assign notSigSum[137] = ~sigSum[137];
  assign notSigSum[136] = ~sigSum[136];
  assign notSigSum[135] = ~sigSum[135];
  assign notSigSum[134] = ~sigSum[134];
  assign notSigSum[133] = ~sigSum[133];
  assign notSigSum[132] = ~sigSum[132];
  assign notSigSum[131] = ~sigSum[131];
  assign notSigSum[130] = ~sigSum[130];
  assign notSigSum[129] = ~sigSum[129];
  assign notSigSum[128] = ~sigSum[128];
  assign notSigSum[127] = ~sigSum[127];
  assign notSigSum[126] = ~sigSum[126];
  assign notSigSum[125] = ~sigSum[125];
  assign notSigSum[124] = ~sigSum[124];
  assign notSigSum[123] = ~sigSum[123];
  assign notSigSum[122] = ~sigSum[122];
  assign notSigSum[121] = ~sigSum[121];
  assign notSigSum[120] = ~sigSum[120];
  assign notSigSum[119] = ~sigSum[119];
  assign notSigSum[118] = ~sigSum[118];
  assign notSigSum[117] = ~sigSum[117];
  assign notSigSum[116] = ~sigSum[116];
  assign notSigSum[115] = ~sigSum[115];
  assign notSigSum[114] = ~sigSum[114];
  assign notSigSum[113] = ~sigSum[113];
  assign notSigSum[112] = ~sigSum[112];
  assign notSigSum[111] = ~sigSum[111];
  assign notSigSum[110] = ~sigSum[110];
  assign notSigSum[109] = ~sigSum[109];
  assign notSigSum[108] = ~T25[108];
  assign notSigSum[107] = ~T25[107];
  assign notSigSum[106] = ~io_mulAddResult[105];
  assign notSigSum[105] = ~io_mulAddResult[104];
  assign notSigSum[104] = ~io_mulAddResult[103];
  assign notSigSum[103] = ~io_mulAddResult[102];
  assign notSigSum[102] = ~io_mulAddResult[101];
  assign notSigSum[101] = ~io_mulAddResult[100];
  assign notSigSum[100] = ~io_mulAddResult[99];
  assign notSigSum[99] = ~io_mulAddResult[98];
  assign notSigSum[98] = ~io_mulAddResult[97];
  assign notSigSum[97] = ~io_mulAddResult[96];
  assign notSigSum[96] = ~io_mulAddResult[95];
  assign notSigSum[95] = ~io_mulAddResult[94];
  assign notSigSum[94] = ~io_mulAddResult[93];
  assign notSigSum[93] = ~io_mulAddResult[92];
  assign notSigSum[92] = ~io_mulAddResult[91];
  assign notSigSum[91] = ~io_mulAddResult[90];
  assign notSigSum[90] = ~io_mulAddResult[89];
  assign notSigSum[89] = ~io_mulAddResult[88];
  assign notSigSum[88] = ~io_mulAddResult[87];
  assign notSigSum[87] = ~io_mulAddResult[86];
  assign notSigSum[86] = ~io_mulAddResult[85];
  assign notSigSum[85] = ~io_mulAddResult[84];
  assign notSigSum[84] = ~io_mulAddResult[83];
  assign notSigSum[83] = ~io_mulAddResult[82];
  assign notSigSum[82] = ~io_mulAddResult[81];
  assign notSigSum[81] = ~io_mulAddResult[80];
  assign notSigSum[80] = ~io_mulAddResult[79];
  assign notSigSum[79] = ~io_mulAddResult[78];
  assign notSigSum[78] = ~io_mulAddResult[77];
  assign notSigSum[77] = ~io_mulAddResult[76];
  assign notSigSum[76] = ~io_mulAddResult[75];
  assign notSigSum[75] = ~io_mulAddResult[74];
  assign notSigSum[74] = ~io_mulAddResult[73];
  assign notSigSum[73] = ~io_mulAddResult[72];
  assign notSigSum[72] = ~io_mulAddResult[71];
  assign notSigSum[71] = ~io_mulAddResult[70];
  assign notSigSum[70] = ~io_mulAddResult[69];
  assign notSigSum[69] = ~io_mulAddResult[68];
  assign notSigSum[68] = ~io_mulAddResult[67];
  assign notSigSum[67] = ~io_mulAddResult[66];
  assign notSigSum[66] = ~io_mulAddResult[65];
  assign notSigSum[65] = ~io_mulAddResult[64];
  assign notSigSum[64] = ~io_mulAddResult[63];
  assign notSigSum[63] = ~io_mulAddResult[62];
  assign notSigSum[62] = ~io_mulAddResult[61];
  assign notSigSum[61] = ~io_mulAddResult[60];
  assign notSigSum[60] = ~io_mulAddResult[59];
  assign notSigSum[59] = ~io_mulAddResult[58];
  assign notSigSum[58] = ~io_mulAddResult[57];
  assign notSigSum[57] = ~io_mulAddResult[56];
  assign notSigSum[56] = ~io_mulAddResult[55];
  assign notSigSum[55] = ~io_mulAddResult[54];
  assign notSigSum[54] = ~io_mulAddResult[53];
  assign notSigSum[53] = ~io_mulAddResult[52];
  assign notSigSum[52] = ~io_mulAddResult[51];
  assign notSigSum[51] = ~io_mulAddResult[50];
  assign notSigSum[50] = ~io_mulAddResult[49];
  assign notSigSum[49] = ~io_mulAddResult[48];
  assign notSigSum[48] = ~io_mulAddResult[47];
  assign notSigSum[47] = ~io_mulAddResult[46];
  assign notSigSum[46] = ~io_mulAddResult[45];
  assign notSigSum[45] = ~io_mulAddResult[44];
  assign notSigSum[44] = ~io_mulAddResult[43];
  assign T199[43] = ~io_mulAddResult[42];
  assign T199[42] = ~io_mulAddResult[41];
  assign T199[41] = ~io_mulAddResult[40];
  assign T199[40] = ~io_mulAddResult[39];
  assign T199[39] = ~io_mulAddResult[38];
  assign T199[38] = ~io_mulAddResult[37];
  assign T199[37] = ~io_mulAddResult[36];
  assign T199[36] = ~io_mulAddResult[35];
  assign T199[35] = ~io_mulAddResult[34];
  assign T199[34] = ~io_mulAddResult[33];
  assign T199[33] = ~io_mulAddResult[32];
  assign T199[32] = ~io_mulAddResult[31];
  assign T199[31] = ~io_mulAddResult[30];
  assign T199[30] = ~io_mulAddResult[29];
  assign T199[29] = ~io_mulAddResult[28];
  assign T199[28] = ~io_mulAddResult[27];
  assign T199[27] = ~io_mulAddResult[26];
  assign T199[26] = ~io_mulAddResult[25];
  assign T199[25] = ~io_mulAddResult[24];
  assign T199[24] = ~io_mulAddResult[23];
  assign T199[23] = ~io_mulAddResult[22];
  assign T199[22] = ~io_mulAddResult[21];
  assign T199[21] = ~io_mulAddResult[20];
  assign T199[20] = ~io_mulAddResult[19];
  assign T199[19] = ~io_mulAddResult[18];
  assign T199[18] = ~io_mulAddResult[17];
  assign T199[17] = ~io_mulAddResult[16];
  assign T199[16] = ~io_mulAddResult[15];
  assign T199[15] = ~io_mulAddResult[14];
  assign T199[14] = ~io_mulAddResult[13];
  assign T199[13] = ~io_mulAddResult[12];
  assign T199[12] = ~io_mulAddResult[11];
  assign T199[11] = ~io_mulAddResult[10];
  assign T199[10] = ~io_mulAddResult[9];
  assign T199[9] = ~io_mulAddResult[8];
  assign T199[8] = ~io_mulAddResult[7];
  assign T199[7] = ~io_mulAddResult[6];
  assign T199[6] = ~io_mulAddResult[5];
  assign T199[5] = ~io_mulAddResult[4];
  assign T199[4] = ~io_mulAddResult[3];
  assign T199[3] = ~io_mulAddResult[2];
  assign T199[2] = ~io_mulAddResult[1];
  assign T199[1] = ~io_mulAddResult[0];
  assign T199[0] = ~io_fromPreMul_bit0AlignedNegSigC;
  assign CDom_firstNormAbsSigSum[86] = T227[86] | T219[86];
  assign CDom_firstNormAbsSigSum[85] = T227[85] | T219[85];
  assign CDom_firstNormAbsSigSum[84] = T227[84] | T219[84];
  assign CDom_firstNormAbsSigSum[83] = T227[83] | T219[83];
  assign CDom_firstNormAbsSigSum[82] = T227[82] | T219[82];
  assign CDom_firstNormAbsSigSum[81] = T227[81] | T219[81];
  assign CDom_firstNormAbsSigSum[80] = T227[80] | T219[80];
  assign CDom_firstNormAbsSigSum[79] = T227[79] | T219[79];
  assign CDom_firstNormAbsSigSum[78] = T227[78] | T219[78];
  assign CDom_firstNormAbsSigSum[77] = T227[77] | T219[77];
  assign CDom_firstNormAbsSigSum[76] = T227[76] | T219[76];
  assign CDom_firstNormAbsSigSum[75] = T227[75] | T219[75];
  assign CDom_firstNormAbsSigSum[74] = T227[74] | T219[74];
  assign CDom_firstNormAbsSigSum[73] = T227[73] | T219[73];
  assign CDom_firstNormAbsSigSum[72] = T227[72] | T219[72];
  assign CDom_firstNormAbsSigSum[71] = T227[71] | T219[71];
  assign CDom_firstNormAbsSigSum[70] = T227[70] | T219[70];
  assign CDom_firstNormAbsSigSum[69] = T227[69] | T219[69];
  assign CDom_firstNormAbsSigSum[68] = T227[68] | T219[68];
  assign CDom_firstNormAbsSigSum[67] = T227[67] | T219[67];
  assign CDom_firstNormAbsSigSum[66] = T227[66] | T219[66];
  assign CDom_firstNormAbsSigSum[65] = T227[65] | T219[65];
  assign CDom_firstNormAbsSigSum[64] = T227[64] | T219[64];
  assign CDom_firstNormAbsSigSum[63] = T227[63] | T219[63];
  assign CDom_firstNormAbsSigSum[62] = T227[62] | T219[62];
  assign CDom_firstNormAbsSigSum[61] = T227[61] | T219[61];
  assign CDom_firstNormAbsSigSum[60] = T227[60] | T219[60];
  assign CDom_firstNormAbsSigSum[59] = T227[59] | T219[59];
  assign CDom_firstNormAbsSigSum[58] = T227[58] | T219[58];
  assign CDom_firstNormAbsSigSum[57] = T227[57] | T219[57];
  assign CDom_firstNormAbsSigSum[56] = T227[56] | T219[56];
  assign CDom_firstNormAbsSigSum[55] = T227[55] | T219[55];
  assign CDom_firstNormAbsSigSum[54] = T227[54] | T219[54];
  assign CDom_firstNormAbsSigSum[53] = T227[53] | T219[53];
  assign CDom_firstNormAbsSigSum[52] = T227[52] | T219[52];
  assign CDom_firstNormAbsSigSum[51] = T227[51] | T219[51];
  assign CDom_firstNormAbsSigSum[50] = T227[50] | T219[50];
  assign CDom_firstNormAbsSigSum[49] = T227[49] | T219[49];
  assign CDom_firstNormAbsSigSum[48] = T227[48] | T219[48];
  assign CDom_firstNormAbsSigSum[47] = T227[47] | T219[47];
  assign CDom_firstNormAbsSigSum[46] = T227[46] | T219[46];
  assign CDom_firstNormAbsSigSum[45] = T227[45] | T219[45];
  assign CDom_firstNormAbsSigSum[44] = T227[44] | T219[44];
  assign CDom_firstNormAbsSigSum[43] = T227[43] | T219[43];
  assign CDom_firstNormAbsSigSum[42] = T227[42] | T219[42];
  assign CDom_firstNormAbsSigSum[41] = T227[41] | T219[41];
  assign CDom_firstNormAbsSigSum[40] = T227[40] | T219[40];
  assign CDom_firstNormAbsSigSum[39] = T227[39] | T219[39];
  assign CDom_firstNormAbsSigSum[38] = T227[38] | T219[38];
  assign CDom_firstNormAbsSigSum[37] = T227[37] | T219[37];
  assign CDom_firstNormAbsSigSum[36] = T227[36] | T219[36];
  assign CDom_firstNormAbsSigSum[35] = T227[35] | T219[35];
  assign CDom_firstNormAbsSigSum[34] = T227[34] | T219[34];
  assign CDom_firstNormAbsSigSum[33] = T227[33] | T219[33];
  assign CDom_firstNormAbsSigSum[32] = T227[32] | T219[32];
  assign CDom_firstNormAbsSigSum[31] = T227[31] | T219[31];
  assign CDom_firstNormAbsSigSum[30] = T227[30] | T219[30];
  assign CDom_firstNormAbsSigSum[29] = T227[29] | T219[29];
  assign CDom_firstNormAbsSigSum[28] = T227[28] | T219[28];
  assign CDom_firstNormAbsSigSum[27] = T227[27] | T219[27];
  assign CDom_firstNormAbsSigSum[26] = T227[26] | T219[26];
  assign CDom_firstNormAbsSigSum[25] = T227[25] | T219[25];
  assign CDom_firstNormAbsSigSum[24] = T227[24] | T219[24];
  assign CDom_firstNormAbsSigSum[23] = T227[23] | T219[23];
  assign CDom_firstNormAbsSigSum[22] = T227[22] | T219[22];
  assign CDom_firstNormAbsSigSum[21] = T227[21] | T219[21];
  assign CDom_firstNormAbsSigSum[20] = T227[20] | T219[20];
  assign CDom_firstNormAbsSigSum[19] = T227[19] | T219[19];
  assign CDom_firstNormAbsSigSum[18] = T227[18] | T219[18];
  assign CDom_firstNormAbsSigSum[17] = T227[17] | T219[17];
  assign CDom_firstNormAbsSigSum[16] = T227[16] | T219[16];
  assign CDom_firstNormAbsSigSum[15] = T227[15] | T219[15];
  assign CDom_firstNormAbsSigSum[14] = T227[14] | T219[14];
  assign CDom_firstNormAbsSigSum[13] = T227[13] | T219[13];
  assign CDom_firstNormAbsSigSum[12] = T227[12] | T219[12];
  assign CDom_firstNormAbsSigSum[11] = T227[11] | T219[11];
  assign CDom_firstNormAbsSigSum[10] = T227[10] | T219[10];
  assign CDom_firstNormAbsSigSum[9] = T227[9] | T219[9];
  assign CDom_firstNormAbsSigSum[8] = T227[8] | T219[8];
  assign CDom_firstNormAbsSigSum[7] = T227[7] | T219[7];
  assign CDom_firstNormAbsSigSum[6] = T227[6] | T219[6];
  assign CDom_firstNormAbsSigSum[5] = T227[5] | T219[5];
  assign CDom_firstNormAbsSigSum[4] = T227[4] | T219[4];
  assign CDom_firstNormAbsSigSum[3] = T227[3] | T219[3];
  assign CDom_firstNormAbsSigSum[2] = T227[2] | T219[2];
  assign CDom_firstNormAbsSigSum[1] = T227[1] | T219[1];
  assign CDom_firstNormAbsSigSum[0] = T227[0] | T219[0];
  assign T219[86] = T686[86] & notSigSum[129];
  assign T219[85] = T686[86] & notSigSum[128];
  assign T219[84] = T686[86] & notSigSum[127];
  assign T219[83] = T686[86] & notSigSum[126];
  assign T219[82] = T686[86] & notSigSum[125];
  assign T219[81] = T686[86] & notSigSum[124];
  assign T219[80] = T686[86] & notSigSum[123];
  assign T219[79] = T686[86] & notSigSum[122];
  assign T219[78] = T686[86] & notSigSum[121];
  assign T219[77] = T686[86] & notSigSum[120];
  assign T219[76] = T686[86] & notSigSum[119];
  assign T219[75] = T686[86] & notSigSum[118];
  assign T219[74] = T686[86] & notSigSum[117];
  assign T219[73] = T686[86] & notSigSum[116];
  assign T219[72] = T686[86] & notSigSum[115];
  assign T219[71] = T686[86] & notSigSum[114];
  assign T219[70] = T686[86] & notSigSum[113];
  assign T219[69] = T686[86] & notSigSum[112];
  assign T219[68] = T686[86] & notSigSum[111];
  assign T219[67] = T686[86] & notSigSum[110];
  assign T219[66] = T686[86] & notSigSum[109];
  assign T219[65] = T686[86] & notSigSum[108];
  assign T219[64] = T686[86] & notSigSum[107];
  assign T219[63] = T686[86] & notSigSum[106];
  assign T219[62] = T686[86] & notSigSum[105];
  assign T219[61] = T686[86] & notSigSum[104];
  assign T219[60] = T686[86] & notSigSum[103];
  assign T219[59] = T686[86] & notSigSum[102];
  assign T219[58] = T686[86] & notSigSum[101];
  assign T219[57] = T686[86] & notSigSum[100];
  assign T219[56] = T686[86] & notSigSum[99];
  assign T219[55] = T686[86] & notSigSum[98];
  assign T219[54] = T686[86] & notSigSum[97];
  assign T219[53] = T686[86] & notSigSum[96];
  assign T219[52] = T686[86] & notSigSum[95];
  assign T219[51] = T686[86] & notSigSum[94];
  assign T219[50] = T686[86] & notSigSum[93];
  assign T219[49] = T686[86] & notSigSum[92];
  assign T219[48] = T686[86] & notSigSum[91];
  assign T219[47] = T686[86] & notSigSum[90];
  assign T219[46] = T686[86] & notSigSum[89];
  assign T219[45] = T686[86] & notSigSum[88];
  assign T219[44] = T686[86] & notSigSum[87];
  assign T219[43] = T686[86] & notSigSum[86];
  assign T219[42] = T686[86] & notSigSum[85];
  assign T219[41] = T686[86] & notSigSum[84];
  assign T219[40] = T686[86] & notSigSum[83];
  assign T219[39] = T686[86] & notSigSum[82];
  assign T219[38] = T686[86] & notSigSum[81];
  assign T219[37] = T686[86] & notSigSum[80];
  assign T219[36] = T686[86] & notSigSum[79];
  assign T219[35] = T686[86] & notSigSum[78];
  assign T219[34] = T686[86] & notSigSum[77];
  assign T219[33] = T686[86] & notSigSum[76];
  assign T219[32] = T686[86] & notSigSum[75];
  assign T219[31] = T686[86] & notSigSum[74];
  assign T219[30] = T686[86] & notSigSum[73];
  assign T219[29] = T686[86] & notSigSum[72];
  assign T219[28] = T686[86] & notSigSum[71];
  assign T219[27] = T686[86] & notSigSum[70];
  assign T219[26] = T686[86] & notSigSum[69];
  assign T219[25] = T686[86] & notSigSum[68];
  assign T219[24] = T686[86] & notSigSum[67];
  assign T219[23] = T686[86] & notSigSum[66];
  assign T219[22] = T686[86] & notSigSum[65];
  assign T219[21] = T686[86] & notSigSum[64];
  assign T219[20] = T686[86] & notSigSum[63];
  assign T219[19] = T686[86] & notSigSum[62];
  assign T219[18] = T686[86] & notSigSum[61];
  assign T219[17] = T686[86] & notSigSum[60];
  assign T219[16] = T686[86] & notSigSum[59];
  assign T219[15] = T686[86] & notSigSum[58];
  assign T219[14] = T686[86] & notSigSum[57];
  assign T219[13] = T686[86] & notSigSum[56];
  assign T219[12] = T686[86] & notSigSum[55];
  assign T219[11] = T686[86] & notSigSum[54];
  assign T219[10] = T686[86] & notSigSum[53];
  assign T219[9] = T686[86] & notSigSum[52];
  assign T219[8] = T686[86] & notSigSum[51];
  assign T219[7] = T686[86] & notSigSum[50];
  assign T219[6] = T686[86] & notSigSum[49];
  assign T219[5] = T686[86] & notSigSum[48];
  assign T219[4] = T686[86] & notSigSum[47];
  assign T219[3] = T686[86] & notSigSum[46];
  assign T219[2] = T686[86] & notSigSum[45];
  assign T219[1] = T686[86] & notSigSum[44];
  assign T219[0] = T686[86] & N811;
  assign T686[86] = T224;
  assign T224 = T682[0] & CDom_estNormDist[5];
  assign T227[86] = T237[86] | T228[86];
  assign T227[85] = T237[85] | T228[85];
  assign T227[84] = T237[84] | T228[84];
  assign T227[83] = T237[83] | T228[83];
  assign T227[82] = T237[82] | T228[82];
  assign T227[81] = T237[81] | T228[81];
  assign T227[80] = T237[80] | T228[80];
  assign T227[79] = T237[79] | T228[79];
  assign T227[78] = T237[78] | T228[78];
  assign T227[77] = T237[77] | T228[77];
  assign T227[76] = T237[76] | T228[76];
  assign T227[75] = T237[75] | T228[75];
  assign T227[74] = T237[74] | T228[74];
  assign T227[73] = T237[73] | T228[73];
  assign T227[72] = T237[72] | T228[72];
  assign T227[71] = T237[71] | T228[71];
  assign T227[70] = T237[70] | T228[70];
  assign T227[69] = T237[69] | T228[69];
  assign T227[68] = T237[68] | T228[68];
  assign T227[67] = T237[67] | T228[67];
  assign T227[66] = T237[66] | T228[66];
  assign T227[65] = T237[65] | T228[65];
  assign T227[64] = T237[64] | T228[64];
  assign T227[63] = T237[63] | T228[63];
  assign T227[62] = T237[62] | T228[62];
  assign T227[61] = T237[61] | T228[61];
  assign T227[60] = T237[60] | T228[60];
  assign T227[59] = T237[59] | T228[59];
  assign T227[58] = T237[58] | T228[58];
  assign T227[57] = T237[57] | T228[57];
  assign T227[56] = T237[56] | T228[56];
  assign T227[55] = T237[55] | T228[55];
  assign T227[54] = T237[54] | T228[54];
  assign T227[53] = T237[53] | T228[53];
  assign T227[52] = T237[52] | T228[52];
  assign T227[51] = T237[51] | T228[51];
  assign T227[50] = T237[50] | T228[50];
  assign T227[49] = T237[49] | T228[49];
  assign T227[48] = T237[48] | T228[48];
  assign T227[47] = T237[47] | T228[47];
  assign T227[46] = T237[46] | T228[46];
  assign T227[45] = T237[45] | T228[45];
  assign T227[44] = T237[44] | T228[44];
  assign T227[43] = T237[43] | T228[43];
  assign T227[42] = T237[42] | T228[42];
  assign T227[41] = T237[41] | T228[41];
  assign T227[40] = T237[40] | T228[40];
  assign T227[39] = T237[39] | T228[39];
  assign T227[38] = T237[38] | T228[38];
  assign T227[37] = T237[37] | T228[37];
  assign T227[36] = T237[36] | T228[36];
  assign T227[35] = T237[35] | T228[35];
  assign T227[34] = T237[34] | T228[34];
  assign T227[33] = T237[33] | T228[33];
  assign T227[32] = T237[32] | T228[32];
  assign T227[31] = T237[31] | T228[31];
  assign T227[30] = T237[30] | T228[30];
  assign T227[29] = T237[29] | T228[29];
  assign T227[28] = T237[28] | T228[28];
  assign T227[27] = T237[27] | T228[27];
  assign T227[26] = T237[26] | T228[26];
  assign T227[25] = T237[25] | T228[25];
  assign T227[24] = T237[24] | T228[24];
  assign T227[23] = T237[23] | T228[23];
  assign T227[22] = T237[22] | T228[22];
  assign T227[21] = T237[21] | T228[21];
  assign T227[20] = T237[20] | T228[20];
  assign T227[19] = T237[19] | T228[19];
  assign T227[18] = T237[18] | T228[18];
  assign T227[17] = T237[17] | T228[17];
  assign T227[16] = T237[16] | T228[16];
  assign T227[15] = T237[15] | T228[15];
  assign T227[14] = T237[14] | T228[14];
  assign T227[13] = T237[13] | T228[13];
  assign T227[12] = T237[12] | T228[12];
  assign T227[11] = T237[11] | T228[11];
  assign T227[10] = T237[10] | T228[10];
  assign T227[9] = T237[9] | T228[9];
  assign T227[8] = T237[8] | T228[8];
  assign T227[7] = T237[7] | T228[7];
  assign T227[6] = T237[6] | T228[6];
  assign T227[5] = T237[5] | T228[5];
  assign T227[4] = T237[4] | T228[4];
  assign T227[3] = T237[3] | T228[3];
  assign T227[2] = T237[2] | T228[2];
  assign T227[1] = T237[1] | T228[1];
  assign T227[0] = T237[0] | T228[0];
  assign T228[86] = T687[86] & notSigSum[161];
  assign T228[85] = T687[86] & notSigSum[160];
  assign T228[84] = T687[86] & notSigSum[159];
  assign T228[83] = T687[86] & notSigSum[158];
  assign T228[82] = T687[86] & notSigSum[157];
  assign T228[81] = T687[86] & notSigSum[156];
  assign T228[80] = T687[86] & notSigSum[155];
  assign T228[79] = T687[86] & notSigSum[154];
  assign T228[78] = T687[86] & notSigSum[153];
  assign T228[77] = T687[86] & notSigSum[152];
  assign T228[76] = T687[86] & notSigSum[151];
  assign T228[75] = T687[86] & notSigSum[150];
  assign T228[74] = T687[86] & notSigSum[149];
  assign T228[73] = T687[86] & notSigSum[148];
  assign T228[72] = T687[86] & notSigSum[147];
  assign T228[71] = T687[86] & notSigSum[146];
  assign T228[70] = T687[86] & notSigSum[145];
  assign T228[69] = T687[86] & notSigSum[144];
  assign T228[68] = T687[86] & notSigSum[143];
  assign T228[67] = T687[86] & notSigSum[142];
  assign T228[66] = T687[86] & notSigSum[141];
  assign T228[65] = T687[86] & notSigSum[140];
  assign T228[64] = T687[86] & notSigSum[139];
  assign T228[63] = T687[86] & notSigSum[138];
  assign T228[62] = T687[86] & notSigSum[137];
  assign T228[61] = T687[86] & notSigSum[136];
  assign T228[60] = T687[86] & notSigSum[135];
  assign T228[59] = T687[86] & notSigSum[134];
  assign T228[58] = T687[86] & notSigSum[133];
  assign T228[57] = T687[86] & notSigSum[132];
  assign T228[56] = T687[86] & notSigSum[131];
  assign T228[55] = T687[86] & notSigSum[130];
  assign T228[54] = T687[86] & notSigSum[129];
  assign T228[53] = T687[86] & notSigSum[128];
  assign T228[52] = T687[86] & notSigSum[127];
  assign T228[51] = T687[86] & notSigSum[126];
  assign T228[50] = T687[86] & notSigSum[125];
  assign T228[49] = T687[86] & notSigSum[124];
  assign T228[48] = T687[86] & notSigSum[123];
  assign T228[47] = T687[86] & notSigSum[122];
  assign T228[46] = T687[86] & notSigSum[121];
  assign T228[45] = T687[86] & notSigSum[120];
  assign T228[44] = T687[86] & notSigSum[119];
  assign T228[43] = T687[86] & notSigSum[118];
  assign T228[42] = T687[86] & notSigSum[117];
  assign T228[41] = T687[86] & notSigSum[116];
  assign T228[40] = T687[86] & notSigSum[115];
  assign T228[39] = T687[86] & notSigSum[114];
  assign T228[38] = T687[86] & notSigSum[113];
  assign T228[37] = T687[86] & notSigSum[112];
  assign T228[36] = T687[86] & notSigSum[111];
  assign T228[35] = T687[86] & notSigSum[110];
  assign T228[34] = T687[86] & notSigSum[109];
  assign T228[33] = T687[86] & notSigSum[108];
  assign T228[32] = T687[86] & notSigSum[107];
  assign T228[31] = T687[86] & notSigSum[106];
  assign T228[30] = T687[86] & notSigSum[105];
  assign T228[29] = T687[86] & notSigSum[104];
  assign T228[28] = T687[86] & notSigSum[103];
  assign T228[27] = T687[86] & notSigSum[102];
  assign T228[26] = T687[86] & notSigSum[101];
  assign T228[25] = T687[86] & notSigSum[100];
  assign T228[24] = T687[86] & notSigSum[99];
  assign T228[23] = T687[86] & notSigSum[98];
  assign T228[22] = T687[86] & notSigSum[97];
  assign T228[21] = T687[86] & notSigSum[96];
  assign T228[20] = T687[86] & notSigSum[95];
  assign T228[19] = T687[86] & notSigSum[94];
  assign T228[18] = T687[86] & notSigSum[93];
  assign T228[17] = T687[86] & notSigSum[92];
  assign T228[16] = T687[86] & notSigSum[91];
  assign T228[15] = T687[86] & notSigSum[90];
  assign T228[14] = T687[86] & notSigSum[89];
  assign T228[13] = T687[86] & notSigSum[88];
  assign T228[12] = T687[86] & notSigSum[87];
  assign T228[11] = T687[86] & notSigSum[86];
  assign T228[10] = T687[86] & notSigSum[85];
  assign T228[9] = T687[86] & notSigSum[84];
  assign T228[8] = T687[86] & notSigSum[83];
  assign T228[7] = T687[86] & notSigSum[82];
  assign T228[6] = T687[86] & notSigSum[81];
  assign T228[5] = T687[86] & notSigSum[80];
  assign T228[4] = T687[86] & notSigSum[79];
  assign T228[3] = T687[86] & notSigSum[78];
  assign T228[2] = T687[86] & notSigSum[77];
  assign T228[1] = T687[86] & notSigSum[76];
  assign T228[0] = T687[86] & N641;
  assign T687[86] = T233;
  assign T233 = T682[0] & T235;
  assign T235 = ~CDom_estNormDist[5];
  assign T237[86] = T247[86] | T238[86];
  assign T237[85] = T247[85] | T238[85];
  assign T237[84] = T247[84] | T238[84];
  assign T237[83] = T247[83] | T238[83];
  assign T237[82] = T247[82] | T238[82];
  assign T237[81] = T247[81] | T238[81];
  assign T237[80] = T247[80] | T238[80];
  assign T237[79] = T247[79] | T238[79];
  assign T237[78] = T247[78] | T238[78];
  assign T237[77] = T247[77] | T238[77];
  assign T237[76] = T247[76] | T238[76];
  assign T237[75] = T247[75] | T238[75];
  assign T237[74] = T247[74] | T238[74];
  assign T237[73] = T247[73] | T238[73];
  assign T237[72] = T247[72] | T238[72];
  assign T237[71] = T247[71] | T238[71];
  assign T237[70] = T247[70] | T238[70];
  assign T237[69] = T247[69] | T238[69];
  assign T237[68] = T247[68] | T238[68];
  assign T237[67] = T247[67] | T238[67];
  assign T237[66] = T247[66] | T238[66];
  assign T237[65] = T247[65] | T238[65];
  assign T237[64] = T247[64] | T238[64];
  assign T237[63] = T247[63] | T238[63];
  assign T237[62] = T247[62] | T238[62];
  assign T237[61] = T247[61] | T238[61];
  assign T237[60] = T247[60] | T238[60];
  assign T237[59] = T247[59] | T238[59];
  assign T237[58] = T247[58] | T238[58];
  assign T237[57] = T247[57] | T238[57];
  assign T237[56] = T247[56] | T238[56];
  assign T237[55] = T247[55] | T238[55];
  assign T237[54] = T247[54] | T238[54];
  assign T237[53] = T247[53] | T238[53];
  assign T237[52] = T247[52] | T238[52];
  assign T237[51] = T247[51] | T238[51];
  assign T237[50] = T247[50] | T238[50];
  assign T237[49] = T247[49] | T238[49];
  assign T237[48] = T247[48] | T238[48];
  assign T237[47] = T247[47] | T238[47];
  assign T237[46] = T247[46] | T238[46];
  assign T237[45] = T247[45] | T238[45];
  assign T237[44] = T247[44] | T238[44];
  assign T237[43] = T247[43] | T238[43];
  assign T237[42] = T247[42] | T238[42];
  assign T237[41] = T247[41] | T238[41];
  assign T237[40] = T247[40] | T238[40];
  assign T237[39] = T247[39] | T238[39];
  assign T237[38] = T247[38] | T238[38];
  assign T237[37] = T247[37] | T238[37];
  assign T237[36] = T247[36] | T238[36];
  assign T237[35] = T247[35] | T238[35];
  assign T237[34] = T247[34] | T238[34];
  assign T237[33] = T247[33] | T238[33];
  assign T237[32] = T247[32] | T238[32];
  assign T237[31] = T247[31] | T238[31];
  assign T237[30] = T247[30] | T238[30];
  assign T237[29] = T247[29] | T238[29];
  assign T237[28] = T247[28] | T238[28];
  assign T237[27] = T247[27] | T238[27];
  assign T237[26] = T247[26] | T238[26];
  assign T237[25] = T247[25] | T238[25];
  assign T237[24] = T247[24] | T238[24];
  assign T237[23] = T247[23] | T238[23];
  assign T237[22] = T247[22] | T238[22];
  assign T237[21] = T247[21] | T238[21];
  assign T237[20] = T247[20] | T238[20];
  assign T237[19] = T247[19] | T238[19];
  assign T237[18] = T247[18] | T238[18];
  assign T237[17] = T247[17] | T238[17];
  assign T237[16] = T247[16] | T238[16];
  assign T237[15] = T247[15] | T238[15];
  assign T237[14] = T247[14] | T238[14];
  assign T237[13] = T247[13] | T238[13];
  assign T237[12] = T247[12] | T238[12];
  assign T237[11] = T247[11] | T238[11];
  assign T237[10] = T247[10] | T238[10];
  assign T237[9] = T247[9] | T238[9];
  assign T237[8] = T247[8] | T238[8];
  assign T237[7] = T247[7] | T238[7];
  assign T237[6] = T247[6] | T238[6];
  assign T237[5] = T247[5] | T238[5];
  assign T237[4] = T247[4] | T238[4];
  assign T237[3] = T247[3] | T238[3];
  assign T237[2] = T247[2] | T238[2];
  assign T237[1] = T247[1] | T238[1];
  assign T237[0] = T247[0] | T238[0];
  assign T238[86] = T688[86] & sigSum[129];
  assign T238[85] = T688[86] & sigSum[128];
  assign T238[84] = T688[86] & sigSum[127];
  assign T238[83] = T688[86] & sigSum[126];
  assign T238[82] = T688[86] & sigSum[125];
  assign T238[81] = T688[86] & sigSum[124];
  assign T238[80] = T688[86] & sigSum[123];
  assign T238[79] = T688[86] & sigSum[122];
  assign T238[78] = T688[86] & sigSum[121];
  assign T238[77] = T688[86] & sigSum[120];
  assign T238[76] = T688[86] & sigSum[119];
  assign T238[75] = T688[86] & sigSum[118];
  assign T238[74] = T688[86] & sigSum[117];
  assign T238[73] = T688[86] & sigSum[116];
  assign T238[72] = T688[86] & sigSum[115];
  assign T238[71] = T688[86] & sigSum[114];
  assign T238[70] = T688[86] & sigSum[113];
  assign T238[69] = T688[86] & sigSum[112];
  assign T238[68] = T688[86] & sigSum[111];
  assign T238[67] = T688[86] & sigSum[110];
  assign T238[66] = T688[86] & sigSum[109];
  assign T238[65] = T688[86] & T25[108];
  assign T238[64] = T688[86] & T25[107];
  assign T238[63] = T688[86] & io_mulAddResult[105];
  assign T238[62] = T688[86] & io_mulAddResult[104];
  assign T238[61] = T688[86] & io_mulAddResult[103];
  assign T238[60] = T688[86] & io_mulAddResult[102];
  assign T238[59] = T688[86] & io_mulAddResult[101];
  assign T238[58] = T688[86] & io_mulAddResult[100];
  assign T238[57] = T688[86] & io_mulAddResult[99];
  assign T238[56] = T688[86] & io_mulAddResult[98];
  assign T238[55] = T688[86] & io_mulAddResult[97];
  assign T238[54] = T688[86] & io_mulAddResult[96];
  assign T238[53] = T688[86] & io_mulAddResult[95];
  assign T238[52] = T688[86] & io_mulAddResult[94];
  assign T238[51] = T688[86] & io_mulAddResult[93];
  assign T238[50] = T688[86] & io_mulAddResult[92];
  assign T238[49] = T688[86] & io_mulAddResult[91];
  assign T238[48] = T688[86] & io_mulAddResult[90];
  assign T238[47] = T688[86] & io_mulAddResult[89];
  assign T238[46] = T688[86] & io_mulAddResult[88];
  assign T238[45] = T688[86] & io_mulAddResult[87];
  assign T238[44] = T688[86] & io_mulAddResult[86];
  assign T238[43] = T688[86] & io_mulAddResult[85];
  assign T238[42] = T688[86] & io_mulAddResult[84];
  assign T238[41] = T688[86] & io_mulAddResult[83];
  assign T238[40] = T688[86] & io_mulAddResult[82];
  assign T238[39] = T688[86] & io_mulAddResult[81];
  assign T238[38] = T688[86] & io_mulAddResult[80];
  assign T238[37] = T688[86] & io_mulAddResult[79];
  assign T238[36] = T688[86] & io_mulAddResult[78];
  assign T238[35] = T688[86] & io_mulAddResult[77];
  assign T238[34] = T688[86] & io_mulAddResult[76];
  assign T238[33] = T688[86] & io_mulAddResult[75];
  assign T238[32] = T688[86] & io_mulAddResult[74];
  assign T238[31] = T688[86] & io_mulAddResult[73];
  assign T238[30] = T688[86] & io_mulAddResult[72];
  assign T238[29] = T688[86] & io_mulAddResult[71];
  assign T238[28] = T688[86] & io_mulAddResult[70];
  assign T238[27] = T688[86] & io_mulAddResult[69];
  assign T238[26] = T688[86] & io_mulAddResult[68];
  assign T238[25] = T688[86] & io_mulAddResult[67];
  assign T238[24] = T688[86] & io_mulAddResult[66];
  assign T238[23] = T688[86] & io_mulAddResult[65];
  assign T238[22] = T688[86] & io_mulAddResult[64];
  assign T238[21] = T688[86] & io_mulAddResult[63];
  assign T238[20] = T688[86] & io_mulAddResult[62];
  assign T238[19] = T688[86] & io_mulAddResult[61];
  assign T238[18] = T688[86] & io_mulAddResult[60];
  assign T238[17] = T688[86] & io_mulAddResult[59];
  assign T238[16] = T688[86] & io_mulAddResult[58];
  assign T238[15] = T688[86] & io_mulAddResult[57];
  assign T238[14] = T688[86] & io_mulAddResult[56];
  assign T238[13] = T688[86] & io_mulAddResult[55];
  assign T238[12] = T688[86] & io_mulAddResult[54];
  assign T238[11] = T688[86] & io_mulAddResult[53];
  assign T238[10] = T688[86] & io_mulAddResult[52];
  assign T238[9] = T688[86] & io_mulAddResult[51];
  assign T238[8] = T688[86] & io_mulAddResult[50];
  assign T238[7] = T688[86] & io_mulAddResult[49];
  assign T238[6] = T688[86] & io_mulAddResult[48];
  assign T238[5] = T688[86] & io_mulAddResult[47];
  assign T238[4] = T688[86] & io_mulAddResult[46];
  assign T238[3] = T688[86] & io_mulAddResult[45];
  assign T238[2] = T688[86] & io_mulAddResult[44];
  assign T238[1] = T688[86] & io_mulAddResult[43];
  assign T238[0] = T688[86] & N737;
  assign T688[86] = T243;
  assign T243 = T246 & CDom_estNormDist[5];
  assign T246 = ~T682[0];
  assign T247[86] = T689[86] & sigSum[161];
  assign T247[85] = T689[86] & sigSum[160];
  assign T247[84] = T689[86] & sigSum[159];
  assign T247[83] = T689[86] & sigSum[158];
  assign T247[82] = T689[86] & sigSum[157];
  assign T247[81] = T689[86] & sigSum[156];
  assign T247[80] = T689[86] & sigSum[155];
  assign T247[79] = T689[86] & sigSum[154];
  assign T247[78] = T689[86] & sigSum[153];
  assign T247[77] = T689[86] & sigSum[152];
  assign T247[76] = T689[86] & sigSum[151];
  assign T247[75] = T689[86] & sigSum[150];
  assign T247[74] = T689[86] & sigSum[149];
  assign T247[73] = T689[86] & sigSum[148];
  assign T247[72] = T689[86] & sigSum[147];
  assign T247[71] = T689[86] & sigSum[146];
  assign T247[70] = T689[86] & sigSum[145];
  assign T247[69] = T689[86] & sigSum[144];
  assign T247[68] = T689[86] & sigSum[143];
  assign T247[67] = T689[86] & sigSum[142];
  assign T247[66] = T689[86] & sigSum[141];
  assign T247[65] = T689[86] & sigSum[140];
  assign T247[64] = T689[86] & sigSum[139];
  assign T247[63] = T689[86] & sigSum[138];
  assign T247[62] = T689[86] & sigSum[137];
  assign T247[61] = T689[86] & sigSum[136];
  assign T247[60] = T689[86] & sigSum[135];
  assign T247[59] = T689[86] & sigSum[134];
  assign T247[58] = T689[86] & sigSum[133];
  assign T247[57] = T689[86] & sigSum[132];
  assign T247[56] = T689[86] & sigSum[131];
  assign T247[55] = T689[86] & sigSum[130];
  assign T247[54] = T689[86] & sigSum[129];
  assign T247[53] = T689[86] & sigSum[128];
  assign T247[52] = T689[86] & sigSum[127];
  assign T247[51] = T689[86] & sigSum[126];
  assign T247[50] = T689[86] & sigSum[125];
  assign T247[49] = T689[86] & sigSum[124];
  assign T247[48] = T689[86] & sigSum[123];
  assign T247[47] = T689[86] & sigSum[122];
  assign T247[46] = T689[86] & sigSum[121];
  assign T247[45] = T689[86] & sigSum[120];
  assign T247[44] = T689[86] & sigSum[119];
  assign T247[43] = T689[86] & sigSum[118];
  assign T247[42] = T689[86] & sigSum[117];
  assign T247[41] = T689[86] & sigSum[116];
  assign T247[40] = T689[86] & sigSum[115];
  assign T247[39] = T689[86] & sigSum[114];
  assign T247[38] = T689[86] & sigSum[113];
  assign T247[37] = T689[86] & sigSum[112];
  assign T247[36] = T689[86] & sigSum[111];
  assign T247[35] = T689[86] & sigSum[110];
  assign T247[34] = T689[86] & sigSum[109];
  assign T247[33] = T689[86] & T25[108];
  assign T247[32] = T689[86] & T25[107];
  assign T247[31] = T689[86] & io_mulAddResult[105];
  assign T247[30] = T689[86] & io_mulAddResult[104];
  assign T247[29] = T689[86] & io_mulAddResult[103];
  assign T247[28] = T689[86] & io_mulAddResult[102];
  assign T247[27] = T689[86] & io_mulAddResult[101];
  assign T247[26] = T689[86] & io_mulAddResult[100];
  assign T247[25] = T689[86] & io_mulAddResult[99];
  assign T247[24] = T689[86] & io_mulAddResult[98];
  assign T247[23] = T689[86] & io_mulAddResult[97];
  assign T247[22] = T689[86] & io_mulAddResult[96];
  assign T247[21] = T689[86] & io_mulAddResult[95];
  assign T247[20] = T689[86] & io_mulAddResult[94];
  assign T247[19] = T689[86] & io_mulAddResult[93];
  assign T247[18] = T689[86] & io_mulAddResult[92];
  assign T247[17] = T689[86] & io_mulAddResult[91];
  assign T247[16] = T689[86] & io_mulAddResult[90];
  assign T247[15] = T689[86] & io_mulAddResult[89];
  assign T247[14] = T689[86] & io_mulAddResult[88];
  assign T247[13] = T689[86] & io_mulAddResult[87];
  assign T247[12] = T689[86] & io_mulAddResult[86];
  assign T247[11] = T689[86] & io_mulAddResult[85];
  assign T247[10] = T689[86] & io_mulAddResult[84];
  assign T247[9] = T689[86] & io_mulAddResult[83];
  assign T247[8] = T689[86] & io_mulAddResult[82];
  assign T247[7] = T689[86] & io_mulAddResult[81];
  assign T247[6] = T689[86] & io_mulAddResult[80];
  assign T247[5] = T689[86] & io_mulAddResult[79];
  assign T247[4] = T689[86] & io_mulAddResult[78];
  assign T247[3] = T689[86] & io_mulAddResult[77];
  assign T247[2] = T689[86] & io_mulAddResult[76];
  assign T247[1] = T689[86] & io_mulAddResult[75];
  assign T247[0] = T689[86] & N663;
  assign T689[86] = T252;
  assign T252 = T256 & T254;
  assign T254 = ~CDom_estNormDist[5];
  assign T256 = ~T682[0];
  assign T279[31] = T280[31] & absSigSumExtraMask[31];
  assign T279[30] = T280[30] & absSigSumExtraMask[30];
  assign T279[29] = T280[29] & absSigSumExtraMask[29];
  assign T279[28] = T280[28] & absSigSumExtraMask[28];
  assign T279[27] = T280[27] & absSigSumExtraMask[27];
  assign T279[26] = T280[26] & absSigSumExtraMask[26];
  assign T279[25] = T280[25] & absSigSumExtraMask[25];
  assign T279[24] = T280[24] & absSigSumExtraMask[24];
  assign T279[23] = T280[23] & absSigSumExtraMask[23];
  assign T279[22] = T280[22] & absSigSumExtraMask[22];
  assign T279[21] = T280[21] & absSigSumExtraMask[21];
  assign T279[20] = T280[20] & absSigSumExtraMask[20];
  assign T279[19] = T280[19] & absSigSumExtraMask[19];
  assign T279[18] = T280[18] & absSigSumExtraMask[18];
  assign T279[17] = T280[17] & absSigSumExtraMask[17];
  assign T279[16] = T280[16] & absSigSumExtraMask[16];
  assign T279[15] = T280[15] & absSigSumExtraMask[15];
  assign T279[14] = T280[14] & absSigSumExtraMask[14];
  assign T279[13] = T280[13] & absSigSumExtraMask[13];
  assign T279[12] = T280[12] & absSigSumExtraMask[12];
  assign T279[11] = T280[11] & absSigSumExtraMask[11];
  assign T279[10] = T280[10] & absSigSumExtraMask[10];
  assign T279[9] = T280[9] & absSigSumExtraMask[9];
  assign T279[8] = T280[8] & absSigSumExtraMask[8];
  assign T279[7] = T280[7] & T116[0];
  assign T279[6] = T280[6] & T116[1];
  assign T279[5] = T280[5] & T116[2];
  assign T279[4] = T280[4] & T116[3];
  assign T279[3] = T280[3] & T115[0];
  assign T279[2] = T280[2] & T115[1];
  assign T279[1] = T280[1] & absSigSumExtraMask_1;
  assign T279[0] = T280[0] & 1'b1;
  assign T280[31] = ~T179[31];
  assign T280[30] = ~T179[30];
  assign T280[29] = ~T179[29];
  assign T280[28] = ~T179[28];
  assign T280[27] = ~T179[27];
  assign T280[26] = ~T179[26];
  assign T280[25] = ~T179[25];
  assign T280[24] = ~T179[24];
  assign T280[23] = ~T179[23];
  assign T280[22] = ~T179[22];
  assign T280[21] = ~T179[21];
  assign T280[20] = ~T179[20];
  assign T280[19] = ~T179[19];
  assign T280[18] = ~T179[18];
  assign T280[17] = ~T179[17];
  assign T280[16] = ~T179[16];
  assign T280[15] = ~T179[15];
  assign T280[14] = ~T179[14];
  assign T280[13] = ~T179[13];
  assign T280[12] = ~T179[12];
  assign T280[11] = ~T179[11];
  assign T280[10] = ~T179[10];
  assign T280[9] = ~T179[9];
  assign T280[8] = ~T179[8];
  assign T280[7] = ~T179[7];
  assign T280[6] = ~T179[6];
  assign T280[5] = ~T179[5];
  assign T280[4] = ~T179[4];
  assign T280[3] = ~T179[3];
  assign T280[2] = ~T179[2];
  assign T280[1] = ~T179[1];
  assign T280[0] = ~T179[0];
  assign T284[56] = sigX3_56 & 1'b0;
  assign T284[55] = T446[0] & T692[55];
  assign T284[54] = sigX3[54] & T692[54];
  assign T284[53] = sigX3[53] & T692[53];
  assign T284[52] = sigX3[52] & T692[52];
  assign T284[51] = sigX3[51] & T692[51];
  assign T284[50] = sigX3[50] & T692[50];
  assign T284[49] = sigX3[49] & T692[49];
  assign T284[48] = sigX3[48] & T692[48];
  assign T284[47] = sigX3[47] & T692[47];
  assign T284[46] = sigX3[46] & T692[46];
  assign T284[45] = sigX3[45] & T692[45];
  assign T284[44] = sigX3[44] & T692[44];
  assign T284[43] = sigX3[43] & T692[43];
  assign T284[42] = sigX3[42] & T692[42];
  assign T284[41] = sigX3[41] & T692[41];
  assign T284[40] = sigX3[40] & T692[40];
  assign T284[39] = sigX3[39] & T692[39];
  assign T284[38] = sigX3[38] & T692[38];
  assign T284[37] = sigX3[37] & T692[37];
  assign T284[36] = sigX3[36] & T692[36];
  assign T284[35] = sigX3[35] & T692[35];
  assign T284[34] = sigX3[34] & T692[34];
  assign T284[33] = sigX3[33] & T692[33];
  assign T284[32] = sigX3[32] & T692[32];
  assign T284[31] = sigX3[31] & T692[31];
  assign T284[30] = sigX3[30] & T692[30];
  assign T284[29] = sigX3[29] & T692[29];
  assign T284[28] = sigX3[28] & T692[28];
  assign T284[27] = sigX3[27] & T692[27];
  assign T284[26] = sigX3[26] & T692[26];
  assign T284[25] = sigX3[25] & T692[25];
  assign T284[24] = sigX3[24] & T692[24];
  assign T284[23] = sigX3[23] & T692[23];
  assign T284[22] = sigX3[22] & T692[22];
  assign T284[21] = sigX3[21] & T692[21];
  assign T284[20] = sigX3[20] & T692[20];
  assign T284[19] = sigX3[19] & T692[19];
  assign T284[18] = sigX3[18] & T692[18];
  assign T284[17] = sigX3[17] & T692[17];
  assign T284[16] = sigX3[16] & T692[16];
  assign T284[15] = sigX3[15] & T692[15];
  assign T284[14] = sigX3[14] & T692[14];
  assign T284[13] = sigX3[13] & T692[13];
  assign T284[12] = sigX3[12] & T692[12];
  assign T284[11] = sigX3[11] & T692[11];
  assign T284[10] = sigX3[10] & T692[10];
  assign T284[9] = sigX3[9] & T692[9];
  assign T284[8] = sigX3[8] & T692[8];
  assign T284[7] = sigX3[7] & T692[7];
  assign T284[6] = sigX3[6] & T692[6];
  assign T284[5] = sigX3[5] & T692[5];
  assign T284[4] = sigX3[4] & T692[4];
  assign T284[3] = sigX3[3] & T692[3];
  assign T284[2] = sigX3[2] & T692[2];
  assign T284[1] = sigX3[1] & T692[1];
  assign T284[0] = sigX3[0] & T692[0];
  assign T692[55] = 1'b0 & T445[54];
  assign T692[54] = T693[54] & T445[53];
  assign T692[53] = T693[53] & T445[52];
  assign T692[52] = T693[52] & T445[51];
  assign T692[51] = T693[51] & T445[50];
  assign T692[50] = T693[50] & T445[49];
  assign T692[49] = T693[49] & T445[48];
  assign T692[48] = T693[48] & T445[47];
  assign T692[47] = T693[47] & T445[46];
  assign T692[46] = T693[46] & T445[45];
  assign T692[45] = T693[45] & T445[44];
  assign T692[44] = T693[44] & T445[43];
  assign T692[43] = T693[43] & T445[42];
  assign T692[42] = T693[42] & T445[41];
  assign T692[41] = T693[41] & T445[40];
  assign T692[40] = T693[40] & T445[39];
  assign T692[39] = T693[39] & T445[38];
  assign T692[38] = T693[38] & T445[37];
  assign T692[37] = T693[37] & T445[36];
  assign T692[36] = T693[36] & T445[35];
  assign T692[35] = T693[35] & T445[34];
  assign T692[34] = T693[34] & T445[33];
  assign T692[33] = T693[33] & T445[32];
  assign T692[32] = T693[32] & T445[31];
  assign T692[31] = T693[31] & T445[30];
  assign T692[30] = T693[30] & T445[29];
  assign T692[29] = T693[29] & T445[28];
  assign T692[28] = T693[28] & T445[27];
  assign T692[27] = T693[27] & T445[26];
  assign T692[26] = T693[26] & T445[25];
  assign T692[25] = T693[25] & T445[24];
  assign T692[24] = T693[24] & T445[23];
  assign T692[23] = T693[23] & T445[22];
  assign T692[22] = T693[22] & T445[21];
  assign T692[21] = T693[21] & T445[20];
  assign T692[20] = T693[20] & T445[19];
  assign T692[19] = T693[19] & T445[18];
  assign T692[18] = T693[18] & T445[17];
  assign T692[17] = T693[17] & T445[16];
  assign T692[16] = T693[16] & T445[15];
  assign T692[15] = T693[15] & T445[14];
  assign T692[14] = T693[14] & T445[13];
  assign T692[13] = T693[13] & T445[12];
  assign T692[12] = T693[12] & T445[11];
  assign T692[11] = T693[11] & T445[10];
  assign T692[10] = T693[10] & T445[9];
  assign T692[9] = T693[9] & T445[8];
  assign T692[8] = T693[8] & T445[7];
  assign T692[7] = T693[7] & T445[6];
  assign T692[6] = T693[6] & T445[5];
  assign T692[5] = T693[5] & T445[4];
  assign T692[4] = T693[4] & T445[3];
  assign T692[3] = T693[3] & T445[2];
  assign T692[2] = T693[2] & T445[1];
  assign T692[1] = T693[1] & T445[0];
  assign T692[0] = T693[0] & roundMask[0];
  assign T693[54] = ~T445[54];
  assign T693[53] = ~T445[53];
  assign T693[52] = ~T445[52];
  assign T693[51] = ~T445[51];
  assign T693[50] = ~T445[50];
  assign T693[49] = ~T445[49];
  assign T693[48] = ~T445[48];
  assign T693[47] = ~T445[47];
  assign T693[46] = ~T445[46];
  assign T693[45] = ~T445[45];
  assign T693[44] = ~T445[44];
  assign T693[43] = ~T445[43];
  assign T693[42] = ~T445[42];
  assign T693[41] = ~T445[41];
  assign T693[40] = ~T445[40];
  assign T693[39] = ~T445[39];
  assign T693[38] = ~T445[38];
  assign T693[37] = ~T445[37];
  assign T693[36] = ~T445[36];
  assign T693[35] = ~T445[35];
  assign T693[34] = ~T445[34];
  assign T693[33] = ~T445[33];
  assign T693[32] = ~T445[32];
  assign T693[31] = ~T445[31];
  assign T693[30] = ~T445[30];
  assign T693[29] = ~T445[29];
  assign T693[28] = ~T445[28];
  assign T693[27] = ~T445[27];
  assign T693[26] = ~T445[26];
  assign T693[25] = ~T445[25];
  assign T693[24] = ~T445[24];
  assign T693[23] = ~T445[23];
  assign T693[22] = ~T445[22];
  assign T693[21] = ~T445[21];
  assign T693[20] = ~T445[20];
  assign T693[19] = ~T445[19];
  assign T693[18] = ~T445[18];
  assign T693[17] = ~T445[17];
  assign T693[16] = ~T445[16];
  assign T693[15] = ~T445[15];
  assign T693[14] = ~T445[14];
  assign T693[13] = ~T445[13];
  assign T693[12] = ~T445[12];
  assign T693[11] = ~T445[11];
  assign T693[10] = ~T445[10];
  assign T693[9] = ~T445[9];
  assign T693[8] = ~T445[8];
  assign T693[7] = ~T445[7];
  assign T693[6] = ~T445[6];
  assign T693[5] = ~T445[5];
  assign T693[4] = ~T445[4];
  assign T693[3] = ~T445[3];
  assign T693[2] = ~T445[2];
  assign T693[1] = ~T445[1];
  assign T693[0] = ~T445[0];
  assign T287 = ~allRound;
  assign allRound = N502 & N446;
  assign T288[56] = T290[56] & 1'b0;
  assign T288[55] = T290[55] & 1'b0;
  assign T288[54] = T290[54] & T445[54];
  assign T288[53] = T290[53] & T445[53];
  assign T288[52] = T290[52] & T445[52];
  assign T288[51] = T290[51] & T445[51];
  assign T288[50] = T290[50] & T445[50];
  assign T288[49] = T290[49] & T445[49];
  assign T288[48] = T290[48] & T445[48];
  assign T288[47] = T290[47] & T445[47];
  assign T288[46] = T290[46] & T445[46];
  assign T288[45] = T290[45] & T445[45];
  assign T288[44] = T290[44] & T445[44];
  assign T288[43] = T290[43] & T445[43];
  assign T288[42] = T290[42] & T445[42];
  assign T288[41] = T290[41] & T445[41];
  assign T288[40] = T290[40] & T445[40];
  assign T288[39] = T290[39] & T445[39];
  assign T288[38] = T290[38] & T445[38];
  assign T288[37] = T290[37] & T445[37];
  assign T288[36] = T290[36] & T445[36];
  assign T288[35] = T290[35] & T445[35];
  assign T288[34] = T290[34] & T445[34];
  assign T288[33] = T290[33] & T445[33];
  assign T288[32] = T290[32] & T445[32];
  assign T288[31] = T290[31] & T445[31];
  assign T288[30] = T290[30] & T445[30];
  assign T288[29] = T290[29] & T445[29];
  assign T288[28] = T290[28] & T445[28];
  assign T288[27] = T290[27] & T445[27];
  assign T288[26] = T290[26] & T445[26];
  assign T288[25] = T290[25] & T445[25];
  assign T288[24] = T290[24] & T445[24];
  assign T288[23] = T290[23] & T445[23];
  assign T288[22] = T290[22] & T445[22];
  assign T288[21] = T290[21] & T445[21];
  assign T288[20] = T290[20] & T445[20];
  assign T288[19] = T290[19] & T445[19];
  assign T288[18] = T290[18] & T445[18];
  assign T288[17] = T290[17] & T445[17];
  assign T288[16] = T290[16] & T445[16];
  assign T288[15] = T290[15] & T445[15];
  assign T288[14] = T290[14] & T445[14];
  assign T288[13] = T290[13] & T445[13];
  assign T288[12] = T290[12] & T445[12];
  assign T288[11] = T290[11] & T445[11];
  assign T288[10] = T290[10] & T445[10];
  assign T288[9] = T290[9] & T445[9];
  assign T288[8] = T290[8] & T445[8];
  assign T288[7] = T290[7] & T445[7];
  assign T288[6] = T290[6] & T445[6];
  assign T288[5] = T290[5] & T445[5];
  assign T288[4] = T290[4] & T445[4];
  assign T288[3] = T290[3] & T445[3];
  assign T288[2] = T290[2] & T445[2];
  assign T288[1] = T290[1] & T445[1];
  assign T288[0] = T290[0] & T445[0];
  assign T290[56] = ~sigX3_56;
  assign T290[55] = ~T446[0];
  assign T290[54] = ~sigX3[54];
  assign T290[53] = ~sigX3[53];
  assign T290[52] = ~sigX3[52];
  assign T290[51] = ~sigX3[51];
  assign T290[50] = ~sigX3[50];
  assign T290[49] = ~sigX3[49];
  assign T290[48] = ~sigX3[48];
  assign T290[47] = ~sigX3[47];
  assign T290[46] = ~sigX3[46];
  assign T290[45] = ~sigX3[45];
  assign T290[44] = ~sigX3[44];
  assign T290[43] = ~sigX3[43];
  assign T290[42] = ~sigX3[42];
  assign T290[41] = ~sigX3[41];
  assign T290[40] = ~sigX3[40];
  assign T290[39] = ~sigX3[39];
  assign T290[38] = ~sigX3[38];
  assign T290[37] = ~sigX3[37];
  assign T290[36] = ~sigX3[36];
  assign T290[35] = ~sigX3[35];
  assign T290[34] = ~sigX3[34];
  assign T290[33] = ~sigX3[33];
  assign T290[32] = ~sigX3[32];
  assign T290[31] = ~sigX3[31];
  assign T290[30] = ~sigX3[30];
  assign T290[29] = ~sigX3[29];
  assign T290[28] = ~sigX3[28];
  assign T290[27] = ~sigX3[27];
  assign T290[26] = ~sigX3[26];
  assign T290[25] = ~sigX3[25];
  assign T290[24] = ~sigX3[24];
  assign T290[23] = ~sigX3[23];
  assign T290[22] = ~sigX3[22];
  assign T290[21] = ~sigX3[21];
  assign T290[20] = ~sigX3[20];
  assign T290[19] = ~sigX3[19];
  assign T290[18] = ~sigX3[18];
  assign T290[17] = ~sigX3[17];
  assign T290[16] = ~sigX3[16];
  assign T290[15] = ~sigX3[15];
  assign T290[14] = ~sigX3[14];
  assign T290[13] = ~sigX3[13];
  assign T290[12] = ~sigX3[12];
  assign T290[11] = ~sigX3[11];
  assign T290[10] = ~sigX3[10];
  assign T290[9] = ~sigX3[9];
  assign T290[8] = ~sigX3[8];
  assign T290[7] = ~sigX3[7];
  assign T290[6] = ~sigX3[6];
  assign T290[5] = ~sigX3[5];
  assign T290[4] = ~sigX3[4];
  assign T290[3] = ~sigX3[3];
  assign T290[2] = ~sigX3[2];
  assign T290[1] = ~sigX3[1];
  assign T290[0] = ~sigX3[0];
  assign doIncrSig = T291 & T682[0];
  assign T291 = T293 & T292;
  assign T292 = ~sigSum[109];
  assign T293 = ~io_fromPreMul_isCDominant;
  assign commonCase = T295 & T294;
  assign T294 = ~notSpecial_addZeros;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & N630;
  assign T295 = ~addSpecial;
  assign addSpecial = mulSpecial | N385;
  assign mulSpecial = N386 | N387;
  assign io_exceptionFlags[1] = commonCase & underflowY;
  assign underflowY = inexactY & T299;
  assign T299 = sExpX3[13] | T300;
  assign N364 = ~sigX3Shift1;
  assign T695[1] = sigX3Shift1;
  assign T695[0] = N364;
  assign io_exceptionFlags[2] = commonCase & N384;
  assign T304[2] = T352[12] | T305[12];
  assign T304[1] = T352[11] | T305[11];
  assign T304[0] = T352[10] | T305[10];
  assign sExpY[9] = T352[9] | T305[9];
  assign sExpY[8] = T352[8] | T305[8];
  assign sExpY[7] = T352[7] | T305[7];
  assign sExpY[6] = T352[6] | T305[6];
  assign sExpY[5] = T352[5] | T305[5];
  assign sExpY[4] = T352[4] | T305[4];
  assign sExpY[3] = T352[3] | T305[3];
  assign sExpY[2] = T352[2] | T305[2];
  assign sExpY[1] = T352[1] | T305[1];
  assign sExpY[0] = T352[0] | T305[0];
  assign T308[1] = T322[54] | T309[54];
  assign T308[0] = T322[53] | T309[53];
  assign sigY3[52] = T322[52] | T309[52];
  assign sigY3[51] = T322[51] | T309[51];
  assign sigY3[50] = T322[50] | T309[50];
  assign sigY3[49] = T322[49] | T309[49];
  assign sigY3[48] = T322[48] | T309[48];
  assign sigY3[47] = T322[47] | T309[47];
  assign sigY3[46] = T322[46] | T309[46];
  assign sigY3[45] = T322[45] | T309[45];
  assign sigY3[44] = T322[44] | T309[44];
  assign sigY3[43] = T322[43] | T309[43];
  assign sigY3[42] = T322[42] | T309[42];
  assign sigY3[41] = T322[41] | T309[41];
  assign sigY3[40] = T322[40] | T309[40];
  assign sigY3[39] = T322[39] | T309[39];
  assign sigY3[38] = T322[38] | T309[38];
  assign sigY3[37] = T322[37] | T309[37];
  assign sigY3[36] = T322[36] | T309[36];
  assign sigY3[35] = T322[35] | T309[35];
  assign sigY3[34] = T322[34] | T309[34];
  assign sigY3[33] = T322[33] | T309[33];
  assign sigY3[32] = T322[32] | T309[32];
  assign sigY3[31] = T322[31] | T309[31];
  assign sigY3[30] = T322[30] | T309[30];
  assign sigY3[29] = T322[29] | T309[29];
  assign sigY3[28] = T322[28] | T309[28];
  assign sigY3[27] = T322[27] | T309[27];
  assign sigY3[26] = T322[26] | T309[26];
  assign sigY3[25] = T322[25] | T309[25];
  assign sigY3[24] = T322[24] | T309[24];
  assign sigY3[23] = T322[23] | T309[23];
  assign sigY3[22] = T322[22] | T309[22];
  assign sigY3[21] = T322[21] | T309[21];
  assign sigY3[20] = T322[20] | T309[20];
  assign sigY3[19] = T322[19] | T309[19];
  assign sigY3[18] = T322[18] | T309[18];
  assign sigY3[17] = T322[17] | T309[17];
  assign sigY3[16] = T322[16] | T309[16];
  assign sigY3[15] = T322[15] | T309[15];
  assign sigY3[14] = T322[14] | T309[14];
  assign sigY3[13] = T322[13] | T309[13];
  assign sigY3[12] = T322[12] | T309[12];
  assign sigY3[11] = T322[11] | T309[11];
  assign sigY3[10] = T322[10] | T309[10];
  assign sigY3[9] = T322[9] | T309[9];
  assign sigY3[8] = T322[8] | T309[8];
  assign sigY3[7] = T322[7] | T309[7];
  assign sigY3[6] = T322[6] | T309[6];
  assign sigY3[5] = T322[5] | T309[5];
  assign sigY3[4] = T322[4] | T309[4];
  assign sigY3[3] = T322[3] | T309[3];
  assign sigY3[2] = T322[2] | T309[2];
  assign sigY3[1] = T322[1] | T309[1];
  assign sigY3[0] = T322[0] | T309[0];
  assign N365 = ~roundEven;
  assign T310[54] = roundUp_sigY3[54] & T311[54];
  assign T310[53] = roundUp_sigY3[53] & T311[53];
  assign T310[52] = roundUp_sigY3[52] & T311[52];
  assign T310[51] = roundUp_sigY3[51] & T311[51];
  assign T310[50] = roundUp_sigY3[50] & T311[50];
  assign T310[49] = roundUp_sigY3[49] & T311[49];
  assign T310[48] = roundUp_sigY3[48] & T311[48];
  assign T310[47] = roundUp_sigY3[47] & T311[47];
  assign T310[46] = roundUp_sigY3[46] & T311[46];
  assign T310[45] = roundUp_sigY3[45] & T311[45];
  assign T310[44] = roundUp_sigY3[44] & T311[44];
  assign T310[43] = roundUp_sigY3[43] & T311[43];
  assign T310[42] = roundUp_sigY3[42] & T311[42];
  assign T310[41] = roundUp_sigY3[41] & T311[41];
  assign T310[40] = roundUp_sigY3[40] & T311[40];
  assign T310[39] = roundUp_sigY3[39] & T311[39];
  assign T310[38] = roundUp_sigY3[38] & T311[38];
  assign T310[37] = roundUp_sigY3[37] & T311[37];
  assign T310[36] = roundUp_sigY3[36] & T311[36];
  assign T310[35] = roundUp_sigY3[35] & T311[35];
  assign T310[34] = roundUp_sigY3[34] & T311[34];
  assign T310[33] = roundUp_sigY3[33] & T311[33];
  assign T310[32] = roundUp_sigY3[32] & T311[32];
  assign T310[31] = roundUp_sigY3[31] & T311[31];
  assign T310[30] = roundUp_sigY3[30] & T311[30];
  assign T310[29] = roundUp_sigY3[29] & T311[29];
  assign T310[28] = roundUp_sigY3[28] & T311[28];
  assign T310[27] = roundUp_sigY3[27] & T311[27];
  assign T310[26] = roundUp_sigY3[26] & T311[26];
  assign T310[25] = roundUp_sigY3[25] & T311[25];
  assign T310[24] = roundUp_sigY3[24] & T311[24];
  assign T310[23] = roundUp_sigY3[23] & T311[23];
  assign T310[22] = roundUp_sigY3[22] & T311[22];
  assign T310[21] = roundUp_sigY3[21] & T311[21];
  assign T310[20] = roundUp_sigY3[20] & T311[20];
  assign T310[19] = roundUp_sigY3[19] & T311[19];
  assign T310[18] = roundUp_sigY3[18] & T311[18];
  assign T310[17] = roundUp_sigY3[17] & T311[17];
  assign T310[16] = roundUp_sigY3[16] & T311[16];
  assign T310[15] = roundUp_sigY3[15] & T311[15];
  assign T310[14] = roundUp_sigY3[14] & T311[14];
  assign T310[13] = roundUp_sigY3[13] & T311[13];
  assign T310[12] = roundUp_sigY3[12] & T311[12];
  assign T310[11] = roundUp_sigY3[11] & T311[11];
  assign T310[10] = roundUp_sigY3[10] & T311[10];
  assign T310[9] = roundUp_sigY3[9] & T311[9];
  assign T310[8] = roundUp_sigY3[8] & T311[8];
  assign T310[7] = roundUp_sigY3[7] & T311[7];
  assign T310[6] = roundUp_sigY3[6] & T311[6];
  assign T310[5] = roundUp_sigY3[5] & T311[5];
  assign T310[4] = roundUp_sigY3[4] & T311[4];
  assign T310[3] = roundUp_sigY3[3] & T311[3];
  assign T310[2] = roundUp_sigY3[2] & T311[2];
  assign T310[1] = roundUp_sigY3[1] & T311[1];
  assign T310[0] = roundUp_sigY3[0] & T311[0];
  assign T311[54] = ~T445[54];
  assign T311[53] = ~T445[53];
  assign T311[52] = ~T445[52];
  assign T311[51] = ~T445[51];
  assign T311[50] = ~T445[50];
  assign T311[49] = ~T445[49];
  assign T311[48] = ~T445[48];
  assign T311[47] = ~T445[47];
  assign T311[46] = ~T445[46];
  assign T311[45] = ~T445[45];
  assign T311[44] = ~T445[44];
  assign T311[43] = ~T445[43];
  assign T311[42] = ~T445[42];
  assign T311[41] = ~T445[41];
  assign T311[40] = ~T445[40];
  assign T311[39] = ~T445[39];
  assign T311[38] = ~T445[38];
  assign T311[37] = ~T445[37];
  assign T311[36] = ~T445[36];
  assign T311[35] = ~T445[35];
  assign T311[34] = ~T445[34];
  assign T311[33] = ~T445[33];
  assign T311[32] = ~T445[32];
  assign T311[31] = ~T445[31];
  assign T311[30] = ~T445[30];
  assign T311[29] = ~T445[29];
  assign T311[28] = ~T445[28];
  assign T311[27] = ~T445[27];
  assign T311[26] = ~T445[26];
  assign T311[25] = ~T445[25];
  assign T311[24] = ~T445[24];
  assign T311[23] = ~T445[23];
  assign T311[22] = ~T445[22];
  assign T311[21] = ~T445[21];
  assign T311[20] = ~T445[20];
  assign T311[19] = ~T445[19];
  assign T311[18] = ~T445[18];
  assign T311[17] = ~T445[17];
  assign T311[16] = ~T445[16];
  assign T311[15] = ~T445[15];
  assign T311[14] = ~T445[14];
  assign T311[13] = ~T445[13];
  assign T311[12] = ~T445[12];
  assign T311[11] = ~T445[11];
  assign T311[10] = ~T445[10];
  assign T311[9] = ~T445[9];
  assign T311[8] = ~T445[8];
  assign T311[7] = ~T445[7];
  assign T311[6] = ~T445[6];
  assign T311[5] = ~T445[5];
  assign T311[4] = ~T445[4];
  assign T311[3] = ~T445[3];
  assign T311[2] = ~T445[2];
  assign T311[1] = ~T445[1];
  assign T311[0] = ~T445[0];
  assign T314[54] = sigX3_56 | 1'b0;
  assign T314[53] = T446[0] | T445[54];
  assign T314[52] = sigX3[54] | T445[53];
  assign T314[51] = sigX3[53] | T445[52];
  assign T314[50] = sigX3[52] | T445[51];
  assign T314[49] = sigX3[51] | T445[50];
  assign T314[48] = sigX3[50] | T445[49];
  assign T314[47] = sigX3[49] | T445[48];
  assign T314[46] = sigX3[48] | T445[47];
  assign T314[45] = sigX3[47] | T445[46];
  assign T314[44] = sigX3[46] | T445[45];
  assign T314[43] = sigX3[45] | T445[44];
  assign T314[42] = sigX3[44] | T445[43];
  assign T314[41] = sigX3[43] | T445[42];
  assign T314[40] = sigX3[42] | T445[41];
  assign T314[39] = sigX3[41] | T445[40];
  assign T314[38] = sigX3[40] | T445[39];
  assign T314[37] = sigX3[39] | T445[38];
  assign T314[36] = sigX3[38] | T445[37];
  assign T314[35] = sigX3[37] | T445[36];
  assign T314[34] = sigX3[36] | T445[35];
  assign T314[33] = sigX3[35] | T445[34];
  assign T314[32] = sigX3[34] | T445[33];
  assign T314[31] = sigX3[33] | T445[32];
  assign T314[30] = sigX3[32] | T445[31];
  assign T314[29] = sigX3[31] | T445[30];
  assign T314[28] = sigX3[30] | T445[29];
  assign T314[27] = sigX3[29] | T445[28];
  assign T314[26] = sigX3[28] | T445[27];
  assign T314[25] = sigX3[27] | T445[26];
  assign T314[24] = sigX3[26] | T445[25];
  assign T314[23] = sigX3[25] | T445[24];
  assign T314[22] = sigX3[24] | T445[23];
  assign T314[21] = sigX3[23] | T445[22];
  assign T314[20] = sigX3[22] | T445[21];
  assign T314[19] = sigX3[21] | T445[20];
  assign T314[18] = sigX3[20] | T445[19];
  assign T314[17] = sigX3[19] | T445[18];
  assign T314[16] = sigX3[18] | T445[17];
  assign T314[15] = sigX3[17] | T445[16];
  assign T314[14] = sigX3[16] | T445[15];
  assign T314[13] = sigX3[15] | T445[14];
  assign T314[12] = sigX3[14] | T445[13];
  assign T314[11] = sigX3[13] | T445[12];
  assign T314[10] = sigX3[12] | T445[11];
  assign T314[9] = sigX3[11] | T445[10];
  assign T314[8] = sigX3[10] | T445[9];
  assign T314[7] = sigX3[9] | T445[8];
  assign T314[6] = sigX3[8] | T445[7];
  assign T314[5] = sigX3[7] | T445[6];
  assign T314[4] = sigX3[6] | T445[5];
  assign T314[3] = sigX3[5] | T445[4];
  assign T314[2] = sigX3[4] | T445[3];
  assign T314[1] = sigX3[3] | T445[2];
  assign T314[0] = sigX3[2] | T445[1];
  assign T316 = T318 & T317;
  assign T317 = ~N558;
  assign T318 = N560 & N502;
  assign T319 = T320 & N446;
  assign T320 = N560 & T321;
  assign T321 = ~N502;
  assign T322[54] = T344[54] | T323[54];
  assign T322[53] = T344[53] | T323[53];
  assign T322[52] = T344[52] | T323[52];
  assign T322[51] = T344[51] | T323[51];
  assign T322[50] = T344[50] | T323[50];
  assign T322[49] = T344[49] | T323[49];
  assign T322[48] = T344[48] | T323[48];
  assign T322[47] = T344[47] | T323[47];
  assign T322[46] = T344[46] | T323[46];
  assign T322[45] = T344[45] | T323[45];
  assign T322[44] = T344[44] | T323[44];
  assign T322[43] = T344[43] | T323[43];
  assign T322[42] = T344[42] | T323[42];
  assign T322[41] = T344[41] | T323[41];
  assign T322[40] = T344[40] | T323[40];
  assign T322[39] = T344[39] | T323[39];
  assign T322[38] = T344[38] | T323[38];
  assign T322[37] = T344[37] | T323[37];
  assign T322[36] = T344[36] | T323[36];
  assign T322[35] = T344[35] | T323[35];
  assign T322[34] = T344[34] | T323[34];
  assign T322[33] = T344[33] | T323[33];
  assign T322[32] = T344[32] | T323[32];
  assign T322[31] = T344[31] | T323[31];
  assign T322[30] = T344[30] | T323[30];
  assign T322[29] = T344[29] | T323[29];
  assign T322[28] = T344[28] | T323[28];
  assign T322[27] = T344[27] | T323[27];
  assign T322[26] = T344[26] | T323[26];
  assign T322[25] = T344[25] | T323[25];
  assign T322[24] = T344[24] | T323[24];
  assign T322[23] = T344[23] | T323[23];
  assign T322[22] = T344[22] | T323[22];
  assign T322[21] = T344[21] | T323[21];
  assign T322[20] = T344[20] | T323[20];
  assign T322[19] = T344[19] | T323[19];
  assign T322[18] = T344[18] | T323[18];
  assign T322[17] = T344[17] | T323[17];
  assign T322[16] = T344[16] | T323[16];
  assign T322[15] = T344[15] | T323[15];
  assign T322[14] = T344[14] | T323[14];
  assign T322[13] = T344[13] | T323[13];
  assign T322[12] = T344[12] | T323[12];
  assign T322[11] = T344[11] | T323[11];
  assign T322[10] = T344[10] | T323[10];
  assign T322[9] = T344[9] | T323[9];
  assign T322[8] = T344[8] | T323[8];
  assign T322[7] = T344[7] | T323[7];
  assign T322[6] = T344[6] | T323[6];
  assign T322[5] = T344[5] | T323[5];
  assign T322[4] = T344[4] | T323[4];
  assign T322[3] = T344[3] | T323[3];
  assign T322[2] = T344[2] | T323[2];
  assign T322[1] = T344[1] | T323[1];
  assign T322[0] = T344[0] | T323[0];
  assign N366 = ~T324;
  assign T324 = T331 | T325;
  assign T325 = doIncrSig & roundDirectUp;
  assign N367 = ~signY;
  assign N368 = ~isZeroY;
  assign T327 = io_fromPreMul_signProd ^ doNegSignSum;
  assign N369 = ~io_fromPreMul_isCDominant;
  assign T328 = T682[0] & T329;
  assign T329 = ~N630;
  assign T331 = T334 | T332;
  assign T332 = T333 & N502;
  assign T333 = doIncrSig & N560;
  assign T334 = T336 | T335;
  assign T335 = doIncrSig & allRound;
  assign T336 = T340 | T337;
  assign T337 = T338 & anyRound;
  assign T338 = T339 & roundDirectUp;
  assign T339 = ~doIncrSig;
  assign T340 = T341 & N558;
  assign T341 = T342 & N502;
  assign T342 = T343 & N560;
  assign T343 = ~doIncrSig;
  assign N370 = ~T348;
  assign T345[54] = sigX3_56 & 1'b0;
  assign T345[53] = T446[0] & T697[55];
  assign T345[52] = sigX3[54] & T697[54];
  assign T345[51] = sigX3[53] & T697[53];
  assign T345[50] = sigX3[52] & T697[52];
  assign T345[49] = sigX3[51] & T697[51];
  assign T345[48] = sigX3[50] & T697[50];
  assign T345[47] = sigX3[49] & T697[49];
  assign T345[46] = sigX3[48] & T697[48];
  assign T345[45] = sigX3[47] & T697[47];
  assign T345[44] = sigX3[46] & T697[46];
  assign T345[43] = sigX3[45] & T697[45];
  assign T345[42] = sigX3[44] & T697[44];
  assign T345[41] = sigX3[43] & T697[43];
  assign T345[40] = sigX3[42] & T697[42];
  assign T345[39] = sigX3[41] & T697[41];
  assign T345[38] = sigX3[40] & T697[40];
  assign T345[37] = sigX3[39] & T697[39];
  assign T345[36] = sigX3[38] & T697[38];
  assign T345[35] = sigX3[37] & T697[37];
  assign T345[34] = sigX3[36] & T697[36];
  assign T345[33] = sigX3[35] & T697[35];
  assign T345[32] = sigX3[34] & T697[34];
  assign T345[31] = sigX3[33] & T697[33];
  assign T345[30] = sigX3[32] & T697[32];
  assign T345[29] = sigX3[31] & T697[31];
  assign T345[28] = sigX3[30] & T697[30];
  assign T345[27] = sigX3[29] & T697[29];
  assign T345[26] = sigX3[28] & T697[28];
  assign T345[25] = sigX3[27] & T697[27];
  assign T345[24] = sigX3[26] & T697[26];
  assign T345[23] = sigX3[25] & T697[25];
  assign T345[22] = sigX3[24] & T697[24];
  assign T345[21] = sigX3[23] & T697[23];
  assign T345[20] = sigX3[22] & T697[22];
  assign T345[19] = sigX3[21] & T697[21];
  assign T345[18] = sigX3[20] & T697[20];
  assign T345[17] = sigX3[19] & T697[19];
  assign T345[16] = sigX3[18] & T697[18];
  assign T345[15] = sigX3[17] & T697[17];
  assign T345[14] = sigX3[16] & T697[16];
  assign T345[13] = sigX3[15] & T697[15];
  assign T345[12] = sigX3[14] & T697[14];
  assign T345[11] = sigX3[13] & T697[13];
  assign T345[10] = sigX3[12] & T697[12];
  assign T345[9] = sigX3[11] & T697[11];
  assign T345[8] = sigX3[10] & T697[10];
  assign T345[7] = sigX3[9] & T697[9];
  assign T345[6] = sigX3[8] & T697[8];
  assign T345[5] = sigX3[7] & T697[7];
  assign T345[4] = sigX3[6] & T697[6];
  assign T345[3] = sigX3[5] & T697[5];
  assign T345[2] = sigX3[4] & T697[4];
  assign T345[1] = sigX3[3] & T697[3];
  assign T345[0] = sigX3[2] & T697[2];
  assign T697[55] = ~T445[54];
  assign T697[54] = ~T445[53];
  assign T697[53] = ~T445[52];
  assign T697[52] = ~T445[51];
  assign T697[51] = ~T445[50];
  assign T697[50] = ~T445[49];
  assign T697[49] = ~T445[48];
  assign T697[48] = ~T445[47];
  assign T697[47] = ~T445[46];
  assign T697[46] = ~T445[45];
  assign T697[45] = ~T445[44];
  assign T697[44] = ~T445[43];
  assign T697[43] = ~T445[42];
  assign T697[42] = ~T445[41];
  assign T697[41] = ~T445[40];
  assign T697[40] = ~T445[39];
  assign T697[39] = ~T445[38];
  assign T697[38] = ~T445[37];
  assign T697[37] = ~T445[36];
  assign T697[36] = ~T445[35];
  assign T697[35] = ~T445[34];
  assign T697[34] = ~T445[33];
  assign T697[33] = ~T445[32];
  assign T697[32] = ~T445[31];
  assign T697[31] = ~T445[30];
  assign T697[30] = ~T445[29];
  assign T697[29] = ~T445[28];
  assign T697[28] = ~T445[27];
  assign T697[27] = ~T445[26];
  assign T697[26] = ~T445[25];
  assign T697[25] = ~T445[24];
  assign T697[24] = ~T445[23];
  assign T697[23] = ~T445[22];
  assign T697[22] = ~T445[21];
  assign T697[21] = ~T445[20];
  assign T697[20] = ~T445[19];
  assign T697[19] = ~T445[18];
  assign T697[18] = ~T445[17];
  assign T697[17] = ~T445[16];
  assign T697[16] = ~T445[15];
  assign T697[15] = ~T445[14];
  assign T697[14] = ~T445[13];
  assign T697[13] = ~T445[12];
  assign T697[12] = ~T445[11];
  assign T697[11] = ~T445[10];
  assign T697[10] = ~T445[9];
  assign T697[9] = ~T445[8];
  assign T697[8] = ~T445[7];
  assign T697[7] = ~T445[6];
  assign T697[6] = ~T445[5];
  assign T697[5] = ~T445[4];
  assign T697[4] = ~T445[3];
  assign T697[3] = ~T445[2];
  assign T697[2] = ~T445[1];
  assign T348 = T351 & T350;
  assign T350 = ~roundEven;
  assign T351 = ~T324;
  assign T352[12] = T355[12] | T353[12];
  assign T352[11] = T355[11] | T353[11];
  assign T352[10] = T355[10] | T353[10];
  assign T352[9] = T355[9] | T353[9];
  assign T352[8] = T355[8] | T353[8];
  assign T352[7] = T355[7] | T353[7];
  assign T352[6] = T355[6] | T353[6];
  assign T352[5] = T355[5] | T353[5];
  assign T352[4] = T355[4] | T353[4];
  assign T352[3] = T355[3] | T353[3];
  assign T352[2] = T355[2] | T353[2];
  assign T352[1] = T355[1] | T353[1];
  assign T352[0] = T355[0] | T353[0];
  assign N371 = ~T308[0];
  assign N372 = ~T308[1];
  assign io_exceptionFlags[4] = T377 | notSigNaN_invalid;
  assign notSigNaN_invalid = T374 | T359;
  assign T359 = T360 & T682[0];
  assign T360 = T363 & isInfC;
  assign isInfC = N385 & T361;
  assign T361 = ~io_fromPreMul_highExpC[0];
  assign T363 = T369 & T364;
  assign T364 = isInfA | isInfB;
  assign isInfB = N387 & T365;
  assign T365 = ~io_fromPreMul_highExpB[0];
  assign isInfA = N386 & T367;
  assign T367 = ~io_fromPreMul_highExpA[0];
  assign T369 = T372 & T370;
  assign T370 = ~isNaNB;
  assign isNaNB = N387 & io_fromPreMul_highExpB[0];
  assign T372 = ~isNaNA;
  assign isNaNA = N386 & io_fromPreMul_highExpA[0];
  assign T374 = T376 | T375;
  assign T375 = N379 & isInfB;
  assign T376 = isInfA & N376;
  assign T377 = T380 | isSigNaNC;
  assign isSigNaNC = isNaNC & T378;
  assign T378 = ~io_fromPreMul_isNaN_isQuietNaNC;
  assign isNaNC = N385 & io_fromPreMul_highExpC[0];
  assign T380 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T381;
  assign T381 = ~io_fromPreMul_isNaN_isQuietNaNB;
  assign isSigNaNA = isNaNA & T382;
  assign T382 = ~io_fromPreMul_isNaN_isQuietNaNA;
  assign io_out[51] = T390[51] | T385[51];
  assign io_out[50] = T390[50] | T385[51];
  assign io_out[49] = T390[49] | T385[51];
  assign io_out[48] = T390[48] | T385[51];
  assign io_out[47] = T390[47] | T385[51];
  assign io_out[46] = T390[46] | T385[51];
  assign io_out[45] = T390[45] | T385[51];
  assign io_out[44] = T390[44] | T385[51];
  assign io_out[43] = T390[43] | T385[51];
  assign io_out[42] = T390[42] | T385[51];
  assign io_out[41] = T390[41] | T385[51];
  assign io_out[40] = T390[40] | T385[51];
  assign io_out[39] = T390[39] | T385[51];
  assign io_out[38] = T390[38] | T385[51];
  assign io_out[37] = T390[37] | T385[51];
  assign io_out[36] = T390[36] | T385[51];
  assign io_out[35] = T390[35] | T385[51];
  assign io_out[34] = T390[34] | T385[51];
  assign io_out[33] = T390[33] | T385[51];
  assign io_out[32] = T390[32] | T385[51];
  assign io_out[31] = T390[31] | T385[51];
  assign io_out[30] = T390[30] | T385[51];
  assign io_out[29] = T390[29] | T385[51];
  assign io_out[28] = T390[28] | T385[51];
  assign io_out[27] = T390[27] | T385[51];
  assign io_out[26] = T390[26] | T385[51];
  assign io_out[25] = T390[25] | T385[51];
  assign io_out[24] = T390[24] | T385[51];
  assign io_out[23] = T390[23] | T385[51];
  assign io_out[22] = T390[22] | T385[51];
  assign io_out[21] = T390[21] | T385[51];
  assign io_out[20] = T390[20] | T385[51];
  assign io_out[19] = T390[19] | T385[51];
  assign io_out[18] = T390[18] | T385[51];
  assign io_out[17] = T390[17] | T385[51];
  assign io_out[16] = T390[16] | T385[51];
  assign io_out[15] = T390[15] | T385[51];
  assign io_out[14] = T390[14] | T385[51];
  assign io_out[13] = T390[13] | T385[51];
  assign io_out[12] = T390[12] | T385[51];
  assign io_out[11] = T390[11] | T385[51];
  assign io_out[10] = T390[10] | T385[51];
  assign io_out[9] = T390[9] | T385[51];
  assign io_out[8] = T390[8] | T385[51];
  assign io_out[7] = T390[7] | T385[51];
  assign io_out[6] = T390[6] | T385[51];
  assign io_out[5] = T390[5] | T385[51];
  assign io_out[4] = T390[4] | T385[51];
  assign io_out[3] = T390[3] | T385[51];
  assign io_out[2] = T390[2] | T385[51];
  assign io_out[1] = T390[1] | T385[51];
  assign io_out[0] = T390[0] | T385_0;
  assign T698[0] = io_exceptionFlags[2] & T386;
  assign T386 = ~overflowY_roundMagUp;
  assign overflowY_roundMagUp = N560 | roundMagUp;
  assign roundMagUp = T389 | T387;
  assign T387 = N561 & T388;
  assign T388 = ~signY;
  assign T389 = N627 & signY;
  assign T390[51] = T394[51] | T391[51];
  assign T390[50] = T394[50] | 1'b0;
  assign T390[49] = T394[49] | 1'b0;
  assign T390[48] = T394[48] | 1'b0;
  assign T390[47] = T394[47] | 1'b0;
  assign T390[46] = T394[46] | 1'b0;
  assign T390[45] = T394[45] | 1'b0;
  assign T390[44] = T394[44] | 1'b0;
  assign T390[43] = T394[43] | 1'b0;
  assign T390[42] = T394[42] | 1'b0;
  assign T390[41] = T394[41] | 1'b0;
  assign T390[40] = T394[40] | 1'b0;
  assign T390[39] = T394[39] | 1'b0;
  assign T390[38] = T394[38] | 1'b0;
  assign T390[37] = T394[37] | 1'b0;
  assign T390[36] = T394[36] | 1'b0;
  assign T390[35] = T394[35] | 1'b0;
  assign T390[34] = T394[34] | 1'b0;
  assign T390[33] = T394[33] | 1'b0;
  assign T390[32] = T394[32] | 1'b0;
  assign T390[31] = T394[31] | 1'b0;
  assign T390[30] = T394[30] | 1'b0;
  assign T390[29] = T394[29] | 1'b0;
  assign T390[28] = T394[28] | 1'b0;
  assign T390[27] = T394[27] | 1'b0;
  assign T390[26] = T394[26] | 1'b0;
  assign T390[25] = T394[25] | 1'b0;
  assign T390[24] = T394[24] | 1'b0;
  assign T390[23] = T394[23] | 1'b0;
  assign T390[22] = T394[22] | 1'b0;
  assign T390[21] = T394[21] | 1'b0;
  assign T390[20] = T394[20] | 1'b0;
  assign T390[19] = T394[19] | 1'b0;
  assign T390[18] = T394[18] | 1'b0;
  assign T390[17] = T394[17] | 1'b0;
  assign T390[16] = T394[16] | 1'b0;
  assign T390[15] = T394[15] | 1'b0;
  assign T390[14] = T394[14] | 1'b0;
  assign T390[13] = T394[13] | 1'b0;
  assign T390[12] = T394[12] | 1'b0;
  assign T390[11] = T394[11] | 1'b0;
  assign T390[10] = T394[10] | 1'b0;
  assign T390[9] = T394[9] | 1'b0;
  assign T390[8] = T394[8] | 1'b0;
  assign T390[7] = T394[7] | 1'b0;
  assign T390[6] = T394[6] | 1'b0;
  assign T390[5] = T394[5] | 1'b0;
  assign T390[4] = T394[4] | 1'b0;
  assign T390[3] = T394[3] | 1'b0;
  assign T390[2] = T394[2] | 1'b0;
  assign T390[1] = T394[1] | 1'b0;
  assign T390[0] = T394[0] | 1'b0;
  assign T391[51] = T392 | notSigNaN_invalid;
  assign T392 = T393 | isNaNC;
  assign T393 = isNaNA | isNaNB;
  assign N373 = ~T397;
  assign T397 = T398 | T391[51];
  assign T398 = totalUnderflowY & roundMagUp;
  assign totalUnderflowY = T403 & T399;
  assign T399 = T304[2] | T400;
  assign T403 = ~isZeroY;
  assign io_out[63] = T405[11] | T404[11];
  assign io_out[62] = T405[10] | T404[11];
  assign io_out[61] = T405[9] | T404[11];
  assign io_out[60] = T405[8] | 1'b0;
  assign io_out[59] = T405[7] | 1'b0;
  assign io_out[58] = T405[6] | 1'b0;
  assign io_out[57] = T405[5] | 1'b0;
  assign io_out[56] = T405[4] | 1'b0;
  assign io_out[55] = T405[3] | 1'b0;
  assign io_out[54] = T405[2] | 1'b0;
  assign io_out[53] = T405[1] | 1'b0;
  assign io_out[52] = T405[0] | 1'b0;
  assign T404[11] = T391[51];
  assign T405[11] = T410[11] | T406[11];
  assign T405[10] = T410[10] | T406[11];
  assign T405[9] = T410[9] | 1'b0;
  assign T405[8] = T410[8] | 1'b0;
  assign T405[7] = T410[7] | 1'b0;
  assign T405[6] = T410[6] | 1'b0;
  assign T405[5] = T410[5] | 1'b0;
  assign T405[4] = T410[4] | 1'b0;
  assign T405[3] = T410[3] | 1'b0;
  assign T405[2] = T410[2] | 1'b0;
  assign T405[1] = T410[1] | 1'b0;
  assign T405[0] = T410[0] | 1'b0;
  assign T406[11] = notNaN_isInfOut;
  assign notNaN_isInfOut = T408 | T407;
  assign T407 = io_exceptionFlags[2] & overflowY_roundMagUp;
  assign T408 = T409 | isInfC;
  assign T409 = isInfA | isInfB;
  assign T410[11] = T412[11] | T411[11];
  assign T410[10] = T412[10] | 1'b0;
  assign T410[9] = T412[9] | T411[11];
  assign T410[8] = T412[8] | T411[11];
  assign T410[7] = T412[7] | T411[11];
  assign T410[6] = T412[6] | T411[11];
  assign T410[5] = T412[5] | T411[11];
  assign T410[4] = T412[4] | T411[11];
  assign T410[3] = T412[3] | T411[11];
  assign T410[2] = T412[2] | T411[11];
  assign T410[1] = T412[1] | T411[11];
  assign T410[0] = T412[0] | T411[11];
  assign T411[11] = T698[0];
  assign T412[11] = T415[11] | 1'b0;
  assign T412[10] = T415[10] | 1'b0;
  assign T412[9] = T415[9] | T413[9];
  assign T412[8] = T415[8] | T413[9];
  assign T412[7] = T415[7] | T413[9];
  assign T412[6] = T415[6] | T413[9];
  assign T412[5] = T415[5] | 1'b0;
  assign T412[4] = T415[4] | 1'b0;
  assign T412[3] = T415[3] | T413[9];
  assign T412[2] = T415[2] | T413[9];
  assign T412[1] = T415[1] | T413[9];
  assign T412[0] = T415[0] | 1'b0;
  assign T413[9] = pegMinFiniteMagOut;
  assign pegMinFiniteMagOut = T414 & roundMagUp;
  assign T414 = commonCase & totalUnderflowY;
  assign T415[11] = T418[11] & T416[11];
  assign T415[10] = T418[10] & T416[10];
  assign T415[9] = T418[9] & T416[9];
  assign T415[8] = T418[8] & T416[8];
  assign T415[7] = T418[7] & T416[7];
  assign T415[6] = T418[6] & T416[6];
  assign T415[5] = T418[5] & T416[5];
  assign T415[4] = T418[4] & T416[4];
  assign T415[3] = T418[3] & T416[3];
  assign T415[2] = T418[2] & T416[2];
  assign T415[1] = T418[1] & T416[1];
  assign T415[0] = T418[0] & T416[0];
  assign T416[11] = ~1'b0;
  assign T416[10] = ~1'b0;
  assign T416[9] = ~T417[9];
  assign T416[8] = ~1'b0;
  assign T416[7] = ~1'b0;
  assign T416[6] = ~1'b0;
  assign T416[5] = ~1'b0;
  assign T416[4] = ~1'b0;
  assign T416[3] = ~1'b0;
  assign T416[2] = ~1'b0;
  assign T416[1] = ~1'b0;
  assign T416[0] = ~1'b0;
  assign T417[9] = notNaN_isInfOut;
  assign T418[11] = T421[11] & T419[11];
  assign T418[10] = T421[10] & T419[10];
  assign T418[9] = T421[9] & T419[9];
  assign T418[8] = T421[8] & T419[8];
  assign T418[7] = T421[7] & T419[7];
  assign T418[6] = T421[6] & T419[6];
  assign T418[5] = T421[5] & T419[5];
  assign T418[4] = T421[4] & T419[4];
  assign T418[3] = T421[3] & T419[3];
  assign T418[2] = T421[2] & T419[2];
  assign T418[1] = T421[1] & T419[1];
  assign T418[0] = T421[0] & T419[0];
  assign T419[11] = ~1'b0;
  assign T419[10] = ~T420[10];
  assign T419[9] = ~1'b0;
  assign T419[8] = ~1'b0;
  assign T419[7] = ~1'b0;
  assign T419[6] = ~1'b0;
  assign T419[5] = ~1'b0;
  assign T419[4] = ~1'b0;
  assign T419[3] = ~1'b0;
  assign T419[2] = ~1'b0;
  assign T419[1] = ~1'b0;
  assign T419[0] = ~1'b0;
  assign T420[10] = T698[0];
  assign T421[11] = T424[11] & T422[11];
  assign T421[10] = T424[10] & T422[10];
  assign T421[9] = T424[9] & T422[9];
  assign T421[8] = T424[8] & T422[8];
  assign T421[7] = T424[7] & T422[7];
  assign T421[6] = T424[6] & T422[6];
  assign T421[5] = T424[5] & T422[5];
  assign T421[4] = T424[4] & T422[4];
  assign T421[3] = T424[3] & T422[3];
  assign T421[2] = T424[2] & T422[2];
  assign T421[1] = T424[1] & T422[1];
  assign T421[0] = T424[0] & T422[0];
  assign T422[11] = ~T423[11];
  assign T422[10] = ~T423[11];
  assign T422[9] = ~1'b0;
  assign T422[8] = ~1'b0;
  assign T422[7] = ~1'b0;
  assign T422[6] = ~1'b0;
  assign T422[5] = ~T423[11];
  assign T422[4] = ~T423[11];
  assign T422[3] = ~1'b0;
  assign T422[2] = ~1'b0;
  assign T422[1] = ~1'b0;
  assign T422[0] = ~T423[11];
  assign T423[11] = pegMinFiniteMagOut;
  assign T424[11] = T304[1] & T425[11];
  assign T424[10] = T304[0] & T425[10];
  assign T424[9] = sExpY[9] & T425[9];
  assign T424[8] = sExpY[8] & T425[8];
  assign T424[7] = sExpY[7] & T425[7];
  assign T424[6] = sExpY[6] & T425[6];
  assign T424[5] = sExpY[5] & T425[5];
  assign T424[4] = sExpY[4] & T425[4];
  assign T424[3] = sExpY[3] & T425[3];
  assign T424[2] = sExpY[2] & T425[2];
  assign T424[1] = sExpY[1] & T425[1];
  assign T424[0] = sExpY[0] & T425[0];
  assign T425[11] = ~T426[11];
  assign T425[10] = ~T426[11];
  assign T425[9] = ~T426[11];
  assign T425[8] = ~1'b0;
  assign T425[7] = ~1'b0;
  assign T425[6] = ~1'b0;
  assign T425[5] = ~1'b0;
  assign T425[4] = ~1'b0;
  assign T425[3] = ~1'b0;
  assign T425[2] = ~1'b0;
  assign T425[1] = ~1'b0;
  assign T425[0] = ~1'b0;
  assign T426[11] = notSpecial_isZeroOut;
  assign notSpecial_isZeroOut = T427 | totalUnderflowY;
  assign T427 = notSpecial_addZeros | isZeroY;
  assign io_out[64] = T429 | T428;
  assign T428 = commonCase & signY;
  assign T429 = T444 & uncommonCaseSignOut;
  assign uncommonCaseSignOut = T434 | T430;
  assign T430 = T431 & N627;
  assign T431 = T432 & T682[0];
  assign T432 = T433 & notSpecial_addZeros;
  assign T433 = ~mulSpecial;
  assign T434 = T438 | T435;
  assign T435 = T436 & io_fromPreMul_opSignC;
  assign T436 = T437 & N385;
  assign T437 = ~mulSpecial;
  assign T438 = T442 | T439;
  assign T439 = T440 & io_fromPreMul_signProd;
  assign T440 = mulSpecial & T441;
  assign T441 = ~N385;
  assign T442 = T443 & io_fromPreMul_opSignC;
  assign T443 = ~T682[0];
  assign T444 = ~T391[51];

endmodule