module fetch1_1e2926114d55612f17be0ce20b92717fa98c0d5f(clk, rst, stall_in, flush_in, inval_btc, stop_in, alt_reset_in, \w_in.redirect , \w_in.virt_mode , \w_in.priv_mode , \w_in.big_endian , \w_in.mode_32bit , \w_in.redirect_nia , \w_in.br_nia , \w_in.br_last , \w_in.br_taken , \d_in.redirect , \d_in.redirect_nia , \i_out.req , \i_out.virt_mode , \i_out.priv_mode , \i_out.big_endian , \i_out.stop_mark , \i_out.predicted , \i_out.pred_ntaken , \i_out.nia , log_out);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire [2:0] _04_;
  wire _05_;
  wire [65:0] _06_;
  wire [66:0] _07_;
  wire _08_;
  reg [70:0] _09_;
  reg [67:0] _10_;
  reg [42:0] _11_;
  wire [63:0] _12_;
  wire [31:0] _13_;
  wire [31:0] _14_;
  wire [63:0] _15_;
  wire [31:0] _16_;
  wire _17_;
  wire _18_;
  wire _19_;
  wire _20_;
  wire [1:0] _21_;
  wire _22_;
  wire _23_;
  wire [63:0] _24_;
  wire [2:0] _25_;
  wire [1:0] _26_;
  wire [63:0] _27_;
  wire [2:0] _28_;
  wire [2:0] _29_;
  wire [1:0] _30_;
  wire [63:0] _31_;
  wire _32_;
  wire [2:0] _33_;
  wire [2:0] _34_;
  wire [1:0] _35_;
  wire [63:0] _36_;
  wire _37_;
  wire [2:0] _38_;
  wire _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire advance_nia;
  input alt_reset_in;
  wire alt_reset_in;
  wire [114:0] btc_rd_data;
  wire btc_rd_valid;
  input clk;
  wire clk;
  input \d_in.redirect ;
  wire \d_in.redirect ;
  input [63:0] \d_in.redirect_nia ;
  wire [63:0] \d_in.redirect_nia ;
  input flush_in;
  wire flush_in;
  output \i_out.big_endian ;
  wire \i_out.big_endian ;
  output [63:0] \i_out.nia ;
  wire [63:0] \i_out.nia ;
  output \i_out.pred_ntaken ;
  wire \i_out.pred_ntaken ;
  output \i_out.predicted ;
  wire \i_out.predicted ;
  output \i_out.priv_mode ;
  wire \i_out.priv_mode ;
  output \i_out.req ;
  wire \i_out.req ;
  output \i_out.stop_mark ;
  wire \i_out.stop_mark ;
  output \i_out.virt_mode ;
  wire \i_out.virt_mode ;
  input inval_btc;
  wire inval_btc;
  wire [42:0] log_nia;
  output [42:0] log_out;
  wire [42:0] log_out;
  wire [70:0] r;
  wire [67:0] r_int;
  wire [70:0] r_next;
  wire [67:0] r_next_int;
  input rst;
  wire rst;
  input stall_in;
  wire stall_in;
  input stop_in;
  wire stop_in;
  input \w_in.big_endian ;
  wire \w_in.big_endian ;
  input \w_in.br_last ;
  wire \w_in.br_last ;
  input [63:0] \w_in.br_nia ;
  wire [63:0] \w_in.br_nia ;
  input \w_in.br_taken ;
  wire \w_in.br_taken ;
  input \w_in.mode_32bit ;
  wire \w_in.mode_32bit ;
  input \w_in.priv_mode ;
  wire \w_in.priv_mode ;
  input \w_in.redirect ;
  wire \w_in.redirect ;
  input [63:0] \w_in.redirect_nia ;
  wire [63:0] \w_in.redirect_nia ;
  input \w_in.virt_mode ;
  wire \w_in.virt_mode ;
  assign _00_ = rst | \w_in.redirect ;
  assign _01_ = _00_ | \d_in.redirect ;
  assign _02_ = ~ stall_in;
  assign _03_ = _01_ | _02_;
  assign _04_ = _03_ ? r_next[3:1] : r[3:1];
  assign _05_ = _03_ ? r_next_int[0] : r_int[0];
  assign _06_ = advance_nia ? r_next[70:5] : r[70:5];
  assign _07_ = advance_nia ? r_next_int[67:1] : r_int[67:1];
  assign _08_ = ~ rst;
  always @(posedge clk)
    _09_ <= { _06_, stop_in, _04_, _08_ };
  always @(posedge clk)
    _10_ <= { _07_, _05_ };
  always @(posedge clk)
    _11_ <= { r[70], r[50:9] };
  assign _12_ = alt_reset_in ? 64'hfffffffff0000000 : 64'h0000000000000000;
  assign _13_ = \w_in.mode_32bit  ? 32'd0 : \w_in.redirect_nia [63:32];
  assign _14_ = r_int[0] ? 32'd0 : \d_in.redirect_nia [63:32];
  assign _15_ = r[70:7] + 64'h0000000000000004;
  assign _16_ = r_int[0] ? 32'd0 : _15_[63:32];
  assign _17_ = btc_rd_valid & r_int[1];
  assign _18_ = btc_rd_data[113:62] == { _16_, _15_[31:12] };
  assign _19_ = _17_ & _18_;
  assign _20_ = ~ btc_rd_data[114];
  assign _21_ = _19_ ? { _20_, btc_rd_data[114] } : 2'h0;
  assign _22_ = r_int[2] ? 1'h1 : 1'h0;
  assign _23_ = r_int[2] ? 1'h0 : r_int[3];
  assign _24_ = r_int[2] ? r_int[67:4] : { _16_, _15_[31:0] };
  assign _25_ = r_int[2] ? 3'h0 : { _21_, 1'h1 };
  assign _26_ = \d_in.redirect  ? 2'h0 : { _23_, _22_ };
  assign _27_ = \d_in.redirect  ? { _14_, \d_in.redirect_nia [31:2], 2'h0 } : _24_;
  assign _28_ = \d_in.redirect  ? 3'h0 : _25_;
  assign _29_ = \w_in.redirect  ? { \w_in.big_endian , \w_in.priv_mode , \w_in.virt_mode  } : r[3:1];
  assign _30_ = \w_in.redirect  ? 2'h0 : _26_;
  assign _31_ = \w_in.redirect  ? { _13_, \w_in.redirect_nia [31:2], 2'h0 } : _27_;
  assign _32_ = \w_in.redirect  ? \w_in.mode_32bit  : r_int[0];
  assign _33_ = \w_in.redirect  ? 3'h0 : _28_;
  assign _34_ = rst ? 3'h2 : _29_;
  assign _35_ = rst ? 2'h0 : _30_;
  assign _36_ = rst ? _12_ : _31_;
  assign _37_ = rst ? 1'h0 : _32_;
  assign _38_ = rst ? 3'h0 : _33_;
  assign _39_ = rst | \w_in.redirect ;
  assign _40_ = _39_ | \d_in.redirect ;
  assign _41_ = ~ r[4];
  assign _42_ = ~ stall_in;
  assign _43_ = _41_ & _42_;
  assign _44_ = _40_ | _43_;
  assign r = _09_;
  assign r_next = { _36_, _35_, r[4], _34_, r[0] };
  assign r_int = _10_;
  assign r_next_int = { btc_rd_data[61:0], 2'h0, _38_, _37_ };
  assign advance_nia = _44_;
  assign log_nia = _11_;
  assign btc_rd_data = 115'h00000000000000000000000000000;
  assign btc_rd_valid = 1'h0;
  assign \i_out.req  = r[0];
  assign \i_out.virt_mode  = r[1];
  assign \i_out.priv_mode  = r[2];
  assign \i_out.big_endian  = r[3];
  assign \i_out.stop_mark  = r[4];
  assign \i_out.predicted  = r[5];
  assign \i_out.pred_ntaken  = r[6];
  assign \i_out.nia  = r[70:7];
  assign log_out = log_nia;
endmodule