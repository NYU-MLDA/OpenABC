module divider(clk, rst, \d_in.valid , \d_in.dividend , \d_in.divisor , \d_in.is_signed , \d_in.is_32bit , \d_in.is_extended , \d_in.is_modulus , \d_in.neg_result , \d_out.valid , \d_out.write_reg_data , \d_out.overflow );
  wire [128:0] _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire [63:0] _06_;
  wire [6:0] _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire _11_;
  wire [6:0] _12_;
  wire _13_;
  wire [6:0] _14_;
  wire [128:0] _15_;
  wire [63:0] _16_;
  wire [6:0] _17_;
  wire _18_;
  wire [128:0] _19_;
  wire [63:0] _20_;
  wire [6:0] _21_;
  wire _22_;
  wire [128:0] _23_;
  wire [63:0] _24_;
  wire _25_;
  wire [6:0] _26_;
  wire _27_;
  wire _28_;
  wire [128:0] _29_;
  wire [63:0] _30_;
  wire [63:0] _31_;
  wire _32_;
  wire [6:0] _33_;
  wire _34_;
  wire _35_;
  wire _36_;
  wire _37_;
  wire _38_;
  wire _39_;
  wire [128:0] _40_;
  wire [63:0] _41_;
  wire [63:0] _42_;
  wire _43_;
  wire [6:0] _44_;
  wire _45_;
  wire _46_;
  wire _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  reg [128:0] _51_;
  reg [63:0] _52_;
  reg [63:0] _53_;
  reg _54_;
  reg [6:0] _55_;
  reg _56_;
  reg _57_;
  reg _58_;
  reg _59_;
  reg _60_;
  reg _61_;
  wire [63:0] _62_;
  wire [64:0] _63_;
  wire [64:0] _64_;
  wire _65_;
  wire _66_;
  wire _67_;
  wire _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire [63:0] _76_;
  wire [63:0] _77_;
  wire _78_;
  wire _79_;
  reg [65:0] _80_;
  input clk;
  wire clk;
  wire [6:0] count;
  input [63:0] \d_in.dividend ;
  wire [63:0] \d_in.dividend ;
  input [63:0] \d_in.divisor ;
  wire [63:0] \d_in.divisor ;
  input \d_in.is_32bit ;
  wire \d_in.is_32bit ;
  input \d_in.is_extended ;
  wire \d_in.is_extended ;
  input \d_in.is_modulus ;
  wire \d_in.is_modulus ;
  input \d_in.is_signed ;
  wire \d_in.is_signed ;
  input \d_in.neg_result ;
  wire \d_in.neg_result ;
  input \d_in.valid ;
  wire \d_in.valid ;
  output \d_out.overflow ;
  wire \d_out.overflow ;
  output \d_out.valid ;
  wire \d_out.valid ;
  output [63:0] \d_out.write_reg_data ;
  wire [63:0] \d_out.write_reg_data ;
  wire [128:0] dend;
  wire did_ovf;
  wire [63:0] div;
  wire is_32bit;
  wire is_modulus;
  wire is_signed;
  wire neg_result;
  wire [63:0] oresult;
  wire overflow;
  wire ovf32;
  wire [63:0] quot;
  wire [63:0] result;
  input rst;
  wire rst;
  wire running;
  wire [64:0] sresult;
  assign _00_ = \d_in.is_extended  ? { 1'h0, \d_in.dividend , 64'h0000000000000000 } : { 65'h00000000000000000, \d_in.dividend  };
  assign _01_ = count == 7'h3f;
  assign _02_ = _25_ ? 1'h0 : running;
  assign _03_ = dend[127:64] >= div;
  assign _04_ = dend[128] | _03_;
  assign _05_ = ovf32 | quot[31];
  assign _06_ = dend[127:64] - div;
  assign _07_ = count + 7'h01;
  assign _08_ = dend[128:57] == 72'h000000000000000000;
  assign _09_ = count[6:3] != 4'h7;
  assign _10_ = _08_ & _09_;
  assign _11_ = | { ovf32, quot[31:24] };
  assign _12_ = count + 7'h08;
  assign _13_ = ovf32 | quot[31];
  assign _14_ = count + 7'h01;
  assign _15_ = _10_ ? { dend[120:0], 8'h00 } : { dend[127:0], 1'h0 };
  assign _16_ = _10_ ? { quot[55:0], 8'h00 } : { quot[62:0], 1'h0 };
  assign _17_ = _10_ ? _12_ : _14_;
  assign _18_ = _10_ ? _11_ : _13_;
  assign _19_ = _04_ ? { _06_, dend[63:0], 1'h0 } : _15_;
  assign _20_ = _04_ ? { quot[62:0], 1'h1 } : _16_;
  assign _21_ = _04_ ? _07_ : _17_;
  assign _22_ = _04_ ? _05_ : _18_;
  assign _23_ = running ? _19_ : dend;
  assign _24_ = running ? _20_ : quot;
  assign _25_ = running & _01_;
  assign _26_ = running ? _21_ : 7'h00;
  assign _27_ = running ? quot[63] : overflow;
  assign _28_ = running ? _22_ : ovf32;
  assign _29_ = \d_in.valid  ? _00_ : _23_;
  assign _30_ = \d_in.valid  ? \d_in.divisor  : div;
  assign _31_ = \d_in.valid  ? 64'h0000000000000000 : _24_;
  assign _32_ = \d_in.valid  ? 1'h1 : _02_;
  assign _33_ = \d_in.valid  ? 7'h7f : _26_;
  assign _34_ = \d_in.valid  ? \d_in.neg_result  : neg_result;
  assign _35_ = \d_in.valid  ? \d_in.is_modulus  : is_modulus;
  assign _36_ = \d_in.valid  ? \d_in.is_32bit  : is_32bit;
  assign _37_ = \d_in.valid  ? \d_in.is_signed  : is_signed;
  assign _38_ = \d_in.valid  ? 1'h0 : _27_;
  assign _39_ = \d_in.valid  ? 1'h0 : _28_;
  assign _40_ = rst ? 129'h000000000000000000000000000000000 : _29_;
  assign _41_ = rst ? 64'h0000000000000000 : _30_;
  assign _42_ = rst ? 64'h0000000000000000 : _31_;
  assign _43_ = rst ? 1'h0 : _32_;
  assign _44_ = rst ? 7'h00 : _33_;
  assign _45_ = rst ? neg_result : _34_;
  assign _46_ = rst ? is_modulus : _35_;
  assign _47_ = rst ? is_32bit : _36_;
  assign _48_ = rst ? is_signed : _37_;
  assign _49_ = rst ? overflow : _38_;
  assign _50_ = rst ? ovf32 : _39_;
  always @(posedge clk)
    _51_ <= _40_;
  always @(posedge clk)
    _52_ <= _41_;
  always @(posedge clk)
    _53_ <= _42_;
  always @(posedge clk)
    _54_ <= _43_;
  always @(posedge clk)
    _55_ <= _44_;
  always @(posedge clk)
    _56_ <= _45_;
  always @(posedge clk)
    _57_ <= _46_;
  always @(posedge clk)
    _58_ <= _47_;
  always @(posedge clk)
    _59_ <= _48_;
  always @(posedge clk)
    _60_ <= _49_;
  always @(posedge clk)
    _61_ <= _50_;
  assign _62_ = is_modulus ? dend[128:65] : quot;
  assign _63_ = - $signed({ 1'h0, result });
  assign _64_ = neg_result ? _63_ : { 1'h0, result };
  assign _65_ = ~ is_32bit;
  assign _66_ = sresult[64] ^ sresult[63];
  assign _67_ = is_signed & _66_;
  assign _68_ = overflow | _67_;
  assign _69_ = sresult[32] != sresult[31];
  assign _70_ = ovf32 | _69_;
  assign _71_ = _70_ ? 1'h1 : 1'h0;
  assign _72_ = is_signed ? _71_ : ovf32;
  assign _73_ = _65_ ? _68_ : _72_;
  assign _74_ = ~ is_modulus;
  assign _75_ = is_32bit & _74_;
  assign _76_ = _75_ ? { 32'h00000000, sresult[31:0] } : sresult[63:0];
  assign _77_ = did_ovf ? 64'h0000000000000000 : _76_;
  assign _78_ = count == 7'h40;
  assign _79_ = _78_ ? 1'h1 : 1'h0;
  always @(posedge clk)
    _80_ <= { did_ovf, oresult, _79_ };
  assign dend = _51_;
  assign div = _52_;
  assign quot = _53_;
  assign result = _62_;
  assign sresult = _64_;
  assign oresult = _77_;
  assign running = _54_;
  assign count = _55_;
  assign neg_result = _56_;
  assign is_modulus = _57_;
  assign is_32bit = _58_;
  assign is_signed = _59_;
  assign overflow = _60_;
  assign ovf32 = _61_;
  assign did_ovf = _73_;
  assign \d_out.valid  = _80_[0];
  assign \d_out.write_reg_data  = _80_[64:1];
  assign \d_out.overflow  = _80_[65];
endmodule