module bht_NR_ENTRIES128
(
  clk_i,
  rst_ni,
  flush_i,
  debug_mode_i,
  vpc_i,
  bht_update_i,
  bht_prediction_o_valid_,
  bht_prediction_o_taken_,
  bht_prediction_o_strongly_taken_
);

  input [63:0] vpc_i;
  input [66:0] bht_update_i;
  input clk_i;
  input rst_ni;
  input flush_i;
  input debug_mode_i;
  output bht_prediction_o_valid_;
  output bht_prediction_o_taken_;
  output bht_prediction_o_strongly_taken_;
  wire bht_prediction_o_valid_,bht_prediction_o_taken_,
  bht_prediction_o_strongly_taken_,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,
  N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,
  N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,
  N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,
  N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,
  N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,
  N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,
  N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,
  N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,
  N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,
  N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,
  N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,
  N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,
  N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,
  N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,
  N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,
  N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,
  N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,
  N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,
  N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,
  N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,
  N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,
  N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,
  N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,
  N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,
  N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,
  N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,
  N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,
  N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,
  N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,
  N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,
  N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,
  N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,
  N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,
  N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,
  N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,
  N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,
  N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,
  N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,
  N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,
  N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,
  N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,
  N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,
  N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,
  N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,
  N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,
  N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,
  N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,
  N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,
  N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,
  N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,
  N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,
  N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,
  N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,
  N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,
  N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,
  N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,
  N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,
  N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,
  N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,
  N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,
  N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,
  N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,
  N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,
  N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,
  N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,
  N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,
  N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,
  N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,
  N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,
  N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,
  N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,
  N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,
  N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,
  N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,
  N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,
  N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,
  N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,
  N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,
  N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,
  N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,
  N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,
  N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,
  N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,
  N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,
  N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,
  N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,
  N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,
  N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,
  N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,
  N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,
  N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,
  N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,
  N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,
  N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,
  N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,
  N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,
  N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,
  N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,
  N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,
  N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,
  N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,
  N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,
  N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,
  N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,
  N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,
  N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,
  N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,
  N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,
  N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,
  N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,
  N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,
  N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,
  N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,
  N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,
  N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,
  N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,
  N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,
  N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,
  N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3524,N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,
  N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,N3545,
  N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,
  N3560,N3561,N3562,N3563,N3564;
  reg [383:0] bht_q;
  assign bht_prediction_o_valid_ = (N276)? bht_q[2] : 
                                   (N278)? bht_q[5] : 
                                   (N280)? bht_q[8] : 
                                   (N282)? bht_q[11] : 
                                   (N284)? bht_q[14] : 
                                   (N286)? bht_q[17] : 
                                   (N288)? bht_q[20] : 
                                   (N290)? bht_q[23] : 
                                   (N292)? bht_q[26] : 
                                   (N294)? bht_q[29] : 
                                   (N296)? bht_q[32] : 
                                   (N298)? bht_q[35] : 
                                   (N300)? bht_q[38] : 
                                   (N302)? bht_q[41] : 
                                   (N304)? bht_q[44] : 
                                   (N306)? bht_q[47] : 
                                   (N308)? bht_q[50] : 
                                   (N310)? bht_q[53] : 
                                   (N312)? bht_q[56] : 
                                   (N314)? bht_q[59] : 
                                   (N316)? bht_q[62] : 
                                   (N318)? bht_q[65] : 
                                   (N320)? bht_q[68] : 
                                   (N322)? bht_q[71] : 
                                   (N324)? bht_q[74] : 
                                   (N326)? bht_q[77] : 
                                   (N328)? bht_q[80] : 
                                   (N330)? bht_q[83] : 
                                   (N332)? bht_q[86] : 
                                   (N334)? bht_q[89] : 
                                   (N336)? bht_q[92] : 
                                   (N338)? bht_q[95] : 
                                   (N340)? bht_q[98] : 
                                   (N342)? bht_q[101] : 
                                   (N344)? bht_q[104] : 
                                   (N346)? bht_q[107] : 
                                   (N348)? bht_q[110] : 
                                   (N350)? bht_q[113] : 
                                   (N352)? bht_q[116] : 
                                   (N354)? bht_q[119] : 
                                   (N356)? bht_q[122] : 
                                   (N358)? bht_q[125] : 
                                   (N360)? bht_q[128] : 
                                   (N362)? bht_q[131] : 
                                   (N364)? bht_q[134] : 
                                   (N366)? bht_q[137] : 
                                   (N368)? bht_q[140] : 
                                   (N370)? bht_q[143] : 
                                   (N372)? bht_q[146] : 
                                   (N374)? bht_q[149] : 
                                   (N376)? bht_q[152] : 
                                   (N378)? bht_q[155] : 
                                   (N380)? bht_q[158] : 
                                   (N382)? bht_q[161] : 
                                   (N384)? bht_q[164] : 
                                   (N386)? bht_q[167] : 
                                   (N388)? bht_q[170] : 
                                   (N390)? bht_q[173] : 
                                   (N392)? bht_q[176] : 
                                   (N394)? bht_q[179] : 
                                   (N396)? bht_q[182] : 
                                   (N398)? bht_q[185] : 
                                   (N400)? bht_q[188] : 
                                   (N402)? bht_q[191] : 
                                   (N277)? bht_q[194] : 
                                   (N279)? bht_q[197] : 
                                   (N281)? bht_q[200] : 
                                   (N283)? bht_q[203] : 
                                   (N285)? bht_q[206] : 
                                   (N287)? bht_q[209] : 
                                   (N289)? bht_q[212] : 
                                   (N291)? bht_q[215] : 
                                   (N293)? bht_q[218] : 
                                   (N295)? bht_q[221] : 
                                   (N297)? bht_q[224] : 
                                   (N299)? bht_q[227] : 
                                   (N301)? bht_q[230] : 
                                   (N303)? bht_q[233] : 
                                   (N305)? bht_q[236] : 
                                   (N307)? bht_q[239] : 
                                   (N309)? bht_q[242] : 
                                   (N311)? bht_q[245] : 
                                   (N313)? bht_q[248] : 
                                   (N315)? bht_q[251] : 
                                   (N317)? bht_q[254] : 
                                   (N319)? bht_q[257] : 
                                   (N321)? bht_q[260] : 
                                   (N323)? bht_q[263] : 
                                   (N325)? bht_q[266] : 
                                   (N327)? bht_q[269] : 
                                   (N329)? bht_q[272] : 
                                   (N331)? bht_q[275] : 
                                   (N333)? bht_q[278] : 
                                   (N335)? bht_q[281] : 
                                   (N337)? bht_q[284] : 
                                   (N339)? bht_q[287] : 
                                   (N341)? bht_q[290] : 
                                   (N343)? bht_q[293] : 
                                   (N345)? bht_q[296] : 
                                   (N347)? bht_q[299] : 
                                   (N349)? bht_q[302] : 
                                   (N351)? bht_q[305] : 
                                   (N353)? bht_q[308] : 
                                   (N355)? bht_q[311] : 
                                   (N357)? bht_q[314] : 
                                   (N359)? bht_q[317] : 
                                   (N361)? bht_q[320] : 
                                   (N363)? bht_q[323] : 
                                   (N365)? bht_q[326] : 
                                   (N367)? bht_q[329] : 
                                   (N369)? bht_q[332] : 
                                   (N371)? bht_q[335] : 
                                   (N373)? bht_q[338] : 
                                   (N375)? bht_q[341] : 
                                   (N377)? bht_q[344] : 
                                   (N379)? bht_q[347] : 
                                   (N381)? bht_q[350] : 
                                   (N383)? bht_q[353] : 
                                   (N385)? bht_q[356] : 
                                   (N387)? bht_q[359] : 
                                   (N389)? bht_q[362] : 
                                   (N391)? bht_q[365] : 
                                   (N393)? bht_q[368] : 
                                   (N395)? bht_q[371] : 
                                   (N397)? bht_q[374] : 
                                   (N399)? bht_q[377] : 
                                   (N401)? bht_q[380] : 
                                   (N403)? bht_q[383] : 1'b0;
  assign N468 = (N404)? bht_q[1] : 
                (N405)? bht_q[4] : 
                (N406)? bht_q[7] : 
                (N407)? bht_q[10] : 
                (N408)? bht_q[13] : 
                (N409)? bht_q[16] : 
                (N410)? bht_q[19] : 
                (N411)? bht_q[22] : 
                (N412)? bht_q[25] : 
                (N413)? bht_q[28] : 
                (N414)? bht_q[31] : 
                (N415)? bht_q[34] : 
                (N416)? bht_q[37] : 
                (N417)? bht_q[40] : 
                (N418)? bht_q[43] : 
                (N419)? bht_q[46] : 
                (N420)? bht_q[49] : 
                (N421)? bht_q[52] : 
                (N422)? bht_q[55] : 
                (N423)? bht_q[58] : 
                (N424)? bht_q[61] : 
                (N425)? bht_q[64] : 
                (N426)? bht_q[67] : 
                (N427)? bht_q[70] : 
                (N428)? bht_q[73] : 
                (N429)? bht_q[76] : 
                (N430)? bht_q[79] : 
                (N431)? bht_q[82] : 
                (N432)? bht_q[85] : 
                (N433)? bht_q[88] : 
                (N434)? bht_q[91] : 
                (N435)? bht_q[94] : 
                (N436)? bht_q[97] : 
                (N437)? bht_q[100] : 
                (N438)? bht_q[103] : 
                (N439)? bht_q[106] : 
                (N440)? bht_q[109] : 
                (N441)? bht_q[112] : 
                (N442)? bht_q[115] : 
                (N443)? bht_q[118] : 
                (N444)? bht_q[121] : 
                (N445)? bht_q[124] : 
                (N446)? bht_q[127] : 
                (N447)? bht_q[130] : 
                (N448)? bht_q[133] : 
                (N449)? bht_q[136] : 
                (N450)? bht_q[139] : 
                (N451)? bht_q[142] : 
                (N452)? bht_q[145] : 
                (N453)? bht_q[148] : 
                (N454)? bht_q[151] : 
                (N455)? bht_q[154] : 
                (N456)? bht_q[157] : 
                (N457)? bht_q[160] : 
                (N458)? bht_q[163] : 
                (N459)? bht_q[166] : 
                (N460)? bht_q[169] : 
                (N461)? bht_q[172] : 
                (N462)? bht_q[175] : 
                (N463)? bht_q[178] : 
                (N464)? bht_q[181] : 
                (N465)? bht_q[184] : 
                (N466)? bht_q[187] : 
                (N467)? bht_q[190] : 
                (N277)? bht_q[193] : 
                (N279)? bht_q[196] : 
                (N281)? bht_q[199] : 
                (N283)? bht_q[202] : 
                (N285)? bht_q[205] : 
                (N287)? bht_q[208] : 
                (N289)? bht_q[211] : 
                (N291)? bht_q[214] : 
                (N293)? bht_q[217] : 
                (N295)? bht_q[220] : 
                (N297)? bht_q[223] : 
                (N299)? bht_q[226] : 
                (N301)? bht_q[229] : 
                (N303)? bht_q[232] : 
                (N305)? bht_q[235] : 
                (N307)? bht_q[238] : 
                (N309)? bht_q[241] : 
                (N311)? bht_q[244] : 
                (N313)? bht_q[247] : 
                (N315)? bht_q[250] : 
                (N317)? bht_q[253] : 
                (N319)? bht_q[256] : 
                (N321)? bht_q[259] : 
                (N323)? bht_q[262] : 
                (N325)? bht_q[265] : 
                (N327)? bht_q[268] : 
                (N329)? bht_q[271] : 
                (N331)? bht_q[274] : 
                (N333)? bht_q[277] : 
                (N335)? bht_q[280] : 
                (N337)? bht_q[283] : 
                (N339)? bht_q[286] : 
                (N341)? bht_q[289] : 
                (N343)? bht_q[292] : 
                (N345)? bht_q[295] : 
                (N347)? bht_q[298] : 
                (N349)? bht_q[301] : 
                (N351)? bht_q[304] : 
                (N353)? bht_q[307] : 
                (N355)? bht_q[310] : 
                (N357)? bht_q[313] : 
                (N359)? bht_q[316] : 
                (N361)? bht_q[319] : 
                (N363)? bht_q[322] : 
                (N365)? bht_q[325] : 
                (N367)? bht_q[328] : 
                (N369)? bht_q[331] : 
                (N371)? bht_q[334] : 
                (N373)? bht_q[337] : 
                (N375)? bht_q[340] : 
                (N377)? bht_q[343] : 
                (N379)? bht_q[346] : 
                (N381)? bht_q[349] : 
                (N383)? bht_q[352] : 
                (N385)? bht_q[355] : 
                (N387)? bht_q[358] : 
                (N389)? bht_q[361] : 
                (N391)? bht_q[364] : 
                (N393)? bht_q[367] : 
                (N395)? bht_q[370] : 
                (N397)? bht_q[373] : 
                (N399)? bht_q[376] : 
                (N401)? bht_q[379] : 
                (N403)? bht_q[382] : 1'b0;
  assign N469 = (N404)? bht_q[0] : 
                (N405)? bht_q[3] : 
                (N406)? bht_q[6] : 
                (N407)? bht_q[9] : 
                (N408)? bht_q[12] : 
                (N409)? bht_q[15] : 
                (N410)? bht_q[18] : 
                (N411)? bht_q[21] : 
                (N412)? bht_q[24] : 
                (N413)? bht_q[27] : 
                (N414)? bht_q[30] : 
                (N415)? bht_q[33] : 
                (N416)? bht_q[36] : 
                (N417)? bht_q[39] : 
                (N418)? bht_q[42] : 
                (N419)? bht_q[45] : 
                (N420)? bht_q[48] : 
                (N421)? bht_q[51] : 
                (N422)? bht_q[54] : 
                (N423)? bht_q[57] : 
                (N424)? bht_q[60] : 
                (N425)? bht_q[63] : 
                (N426)? bht_q[66] : 
                (N427)? bht_q[69] : 
                (N428)? bht_q[72] : 
                (N429)? bht_q[75] : 
                (N430)? bht_q[78] : 
                (N431)? bht_q[81] : 
                (N432)? bht_q[84] : 
                (N433)? bht_q[87] : 
                (N434)? bht_q[90] : 
                (N435)? bht_q[93] : 
                (N436)? bht_q[96] : 
                (N437)? bht_q[99] : 
                (N438)? bht_q[102] : 
                (N439)? bht_q[105] : 
                (N440)? bht_q[108] : 
                (N441)? bht_q[111] : 
                (N442)? bht_q[114] : 
                (N443)? bht_q[117] : 
                (N444)? bht_q[120] : 
                (N445)? bht_q[123] : 
                (N446)? bht_q[126] : 
                (N447)? bht_q[129] : 
                (N448)? bht_q[132] : 
                (N449)? bht_q[135] : 
                (N450)? bht_q[138] : 
                (N451)? bht_q[141] : 
                (N452)? bht_q[144] : 
                (N453)? bht_q[147] : 
                (N454)? bht_q[150] : 
                (N455)? bht_q[153] : 
                (N456)? bht_q[156] : 
                (N457)? bht_q[159] : 
                (N458)? bht_q[162] : 
                (N459)? bht_q[165] : 
                (N460)? bht_q[168] : 
                (N461)? bht_q[171] : 
                (N462)? bht_q[174] : 
                (N463)? bht_q[177] : 
                (N464)? bht_q[180] : 
                (N465)? bht_q[183] : 
                (N466)? bht_q[186] : 
                (N467)? bht_q[189] : 
                (N277)? bht_q[192] : 
                (N279)? bht_q[195] : 
                (N281)? bht_q[198] : 
                (N283)? bht_q[201] : 
                (N285)? bht_q[204] : 
                (N287)? bht_q[207] : 
                (N289)? bht_q[210] : 
                (N291)? bht_q[213] : 
                (N293)? bht_q[216] : 
                (N295)? bht_q[219] : 
                (N297)? bht_q[222] : 
                (N299)? bht_q[225] : 
                (N301)? bht_q[228] : 
                (N303)? bht_q[231] : 
                (N305)? bht_q[234] : 
                (N307)? bht_q[237] : 
                (N309)? bht_q[240] : 
                (N311)? bht_q[243] : 
                (N313)? bht_q[246] : 
                (N315)? bht_q[249] : 
                (N317)? bht_q[252] : 
                (N319)? bht_q[255] : 
                (N321)? bht_q[258] : 
                (N323)? bht_q[261] : 
                (N325)? bht_q[264] : 
                (N327)? bht_q[267] : 
                (N329)? bht_q[270] : 
                (N331)? bht_q[273] : 
                (N333)? bht_q[276] : 
                (N335)? bht_q[279] : 
                (N337)? bht_q[282] : 
                (N339)? bht_q[285] : 
                (N341)? bht_q[288] : 
                (N343)? bht_q[291] : 
                (N345)? bht_q[294] : 
                (N347)? bht_q[297] : 
                (N349)? bht_q[300] : 
                (N351)? bht_q[303] : 
                (N353)? bht_q[306] : 
                (N355)? bht_q[309] : 
                (N357)? bht_q[312] : 
                (N359)? bht_q[315] : 
                (N361)? bht_q[318] : 
                (N363)? bht_q[321] : 
                (N365)? bht_q[324] : 
                (N367)? bht_q[327] : 
                (N369)? bht_q[330] : 
                (N371)? bht_q[333] : 
                (N373)? bht_q[336] : 
                (N375)? bht_q[339] : 
                (N377)? bht_q[342] : 
                (N379)? bht_q[345] : 
                (N381)? bht_q[348] : 
                (N383)? bht_q[351] : 
                (N385)? bht_q[354] : 
                (N387)? bht_q[357] : 
                (N389)? bht_q[360] : 
                (N391)? bht_q[363] : 
                (N393)? bht_q[366] : 
                (N395)? bht_q[369] : 
                (N397)? bht_q[372] : 
                (N399)? bht_q[375] : 
                (N401)? bht_q[378] : 
                (N403)? bht_q[381] : 1'b0;
  assign N534 = (N470)? bht_q[1] : 
                (N471)? bht_q[4] : 
                (N472)? bht_q[7] : 
                (N473)? bht_q[10] : 
                (N474)? bht_q[13] : 
                (N475)? bht_q[16] : 
                (N476)? bht_q[19] : 
                (N477)? bht_q[22] : 
                (N478)? bht_q[25] : 
                (N479)? bht_q[28] : 
                (N480)? bht_q[31] : 
                (N481)? bht_q[34] : 
                (N482)? bht_q[37] : 
                (N483)? bht_q[40] : 
                (N484)? bht_q[43] : 
                (N485)? bht_q[46] : 
                (N486)? bht_q[49] : 
                (N487)? bht_q[52] : 
                (N488)? bht_q[55] : 
                (N489)? bht_q[58] : 
                (N490)? bht_q[61] : 
                (N491)? bht_q[64] : 
                (N492)? bht_q[67] : 
                (N493)? bht_q[70] : 
                (N494)? bht_q[73] : 
                (N495)? bht_q[76] : 
                (N496)? bht_q[79] : 
                (N497)? bht_q[82] : 
                (N498)? bht_q[85] : 
                (N499)? bht_q[88] : 
                (N500)? bht_q[91] : 
                (N501)? bht_q[94] : 
                (N502)? bht_q[97] : 
                (N503)? bht_q[100] : 
                (N504)? bht_q[103] : 
                (N505)? bht_q[106] : 
                (N506)? bht_q[109] : 
                (N507)? bht_q[112] : 
                (N508)? bht_q[115] : 
                (N509)? bht_q[118] : 
                (N510)? bht_q[121] : 
                (N511)? bht_q[124] : 
                (N512)? bht_q[127] : 
                (N513)? bht_q[130] : 
                (N514)? bht_q[133] : 
                (N515)? bht_q[136] : 
                (N516)? bht_q[139] : 
                (N517)? bht_q[142] : 
                (N518)? bht_q[145] : 
                (N519)? bht_q[148] : 
                (N520)? bht_q[151] : 
                (N521)? bht_q[154] : 
                (N522)? bht_q[157] : 
                (N523)? bht_q[160] : 
                (N524)? bht_q[163] : 
                (N525)? bht_q[166] : 
                (N526)? bht_q[169] : 
                (N527)? bht_q[172] : 
                (N528)? bht_q[175] : 
                (N529)? bht_q[178] : 
                (N530)? bht_q[181] : 
                (N531)? bht_q[184] : 
                (N532)? bht_q[187] : 
                (N533)? bht_q[190] : 
                (N277)? bht_q[193] : 
                (N279)? bht_q[196] : 
                (N281)? bht_q[199] : 
                (N283)? bht_q[202] : 
                (N285)? bht_q[205] : 
                (N287)? bht_q[208] : 
                (N289)? bht_q[211] : 
                (N291)? bht_q[214] : 
                (N293)? bht_q[217] : 
                (N295)? bht_q[220] : 
                (N297)? bht_q[223] : 
                (N299)? bht_q[226] : 
                (N301)? bht_q[229] : 
                (N303)? bht_q[232] : 
                (N305)? bht_q[235] : 
                (N307)? bht_q[238] : 
                (N309)? bht_q[241] : 
                (N311)? bht_q[244] : 
                (N313)? bht_q[247] : 
                (N315)? bht_q[250] : 
                (N317)? bht_q[253] : 
                (N319)? bht_q[256] : 
                (N321)? bht_q[259] : 
                (N323)? bht_q[262] : 
                (N325)? bht_q[265] : 
                (N327)? bht_q[268] : 
                (N329)? bht_q[271] : 
                (N331)? bht_q[274] : 
                (N333)? bht_q[277] : 
                (N335)? bht_q[280] : 
                (N337)? bht_q[283] : 
                (N339)? bht_q[286] : 
                (N341)? bht_q[289] : 
                (N343)? bht_q[292] : 
                (N345)? bht_q[295] : 
                (N347)? bht_q[298] : 
                (N349)? bht_q[301] : 
                (N351)? bht_q[304] : 
                (N353)? bht_q[307] : 
                (N355)? bht_q[310] : 
                (N357)? bht_q[313] : 
                (N359)? bht_q[316] : 
                (N361)? bht_q[319] : 
                (N363)? bht_q[322] : 
                (N365)? bht_q[325] : 
                (N367)? bht_q[328] : 
                (N369)? bht_q[331] : 
                (N371)? bht_q[334] : 
                (N373)? bht_q[337] : 
                (N375)? bht_q[340] : 
                (N377)? bht_q[343] : 
                (N379)? bht_q[346] : 
                (N381)? bht_q[349] : 
                (N383)? bht_q[352] : 
                (N385)? bht_q[355] : 
                (N387)? bht_q[358] : 
                (N389)? bht_q[361] : 
                (N391)? bht_q[364] : 
                (N393)? bht_q[367] : 
                (N395)? bht_q[370] : 
                (N397)? bht_q[373] : 
                (N399)? bht_q[376] : 
                (N401)? bht_q[379] : 
                (N403)? bht_q[382] : 1'b0;
  assign N535 = (N470)? bht_q[0] : 
                (N471)? bht_q[3] : 
                (N472)? bht_q[6] : 
                (N473)? bht_q[9] : 
                (N474)? bht_q[12] : 
                (N475)? bht_q[15] : 
                (N476)? bht_q[18] : 
                (N477)? bht_q[21] : 
                (N478)? bht_q[24] : 
                (N479)? bht_q[27] : 
                (N480)? bht_q[30] : 
                (N481)? bht_q[33] : 
                (N482)? bht_q[36] : 
                (N483)? bht_q[39] : 
                (N484)? bht_q[42] : 
                (N485)? bht_q[45] : 
                (N486)? bht_q[48] : 
                (N487)? bht_q[51] : 
                (N488)? bht_q[54] : 
                (N489)? bht_q[57] : 
                (N490)? bht_q[60] : 
                (N491)? bht_q[63] : 
                (N492)? bht_q[66] : 
                (N493)? bht_q[69] : 
                (N494)? bht_q[72] : 
                (N495)? bht_q[75] : 
                (N496)? bht_q[78] : 
                (N497)? bht_q[81] : 
                (N498)? bht_q[84] : 
                (N499)? bht_q[87] : 
                (N500)? bht_q[90] : 
                (N501)? bht_q[93] : 
                (N502)? bht_q[96] : 
                (N503)? bht_q[99] : 
                (N504)? bht_q[102] : 
                (N505)? bht_q[105] : 
                (N506)? bht_q[108] : 
                (N507)? bht_q[111] : 
                (N508)? bht_q[114] : 
                (N509)? bht_q[117] : 
                (N510)? bht_q[120] : 
                (N511)? bht_q[123] : 
                (N512)? bht_q[126] : 
                (N513)? bht_q[129] : 
                (N514)? bht_q[132] : 
                (N515)? bht_q[135] : 
                (N516)? bht_q[138] : 
                (N517)? bht_q[141] : 
                (N518)? bht_q[144] : 
                (N519)? bht_q[147] : 
                (N520)? bht_q[150] : 
                (N521)? bht_q[153] : 
                (N522)? bht_q[156] : 
                (N523)? bht_q[159] : 
                (N524)? bht_q[162] : 
                (N525)? bht_q[165] : 
                (N526)? bht_q[168] : 
                (N527)? bht_q[171] : 
                (N528)? bht_q[174] : 
                (N529)? bht_q[177] : 
                (N530)? bht_q[180] : 
                (N531)? bht_q[183] : 
                (N532)? bht_q[186] : 
                (N533)? bht_q[189] : 
                (N277)? bht_q[192] : 
                (N279)? bht_q[195] : 
                (N281)? bht_q[198] : 
                (N283)? bht_q[201] : 
                (N285)? bht_q[204] : 
                (N287)? bht_q[207] : 
                (N289)? bht_q[210] : 
                (N291)? bht_q[213] : 
                (N293)? bht_q[216] : 
                (N295)? bht_q[219] : 
                (N297)? bht_q[222] : 
                (N299)? bht_q[225] : 
                (N301)? bht_q[228] : 
                (N303)? bht_q[231] : 
                (N305)? bht_q[234] : 
                (N307)? bht_q[237] : 
                (N309)? bht_q[240] : 
                (N311)? bht_q[243] : 
                (N313)? bht_q[246] : 
                (N315)? bht_q[249] : 
                (N317)? bht_q[252] : 
                (N319)? bht_q[255] : 
                (N321)? bht_q[258] : 
                (N323)? bht_q[261] : 
                (N325)? bht_q[264] : 
                (N327)? bht_q[267] : 
                (N329)? bht_q[270] : 
                (N331)? bht_q[273] : 
                (N333)? bht_q[276] : 
                (N335)? bht_q[279] : 
                (N337)? bht_q[282] : 
                (N339)? bht_q[285] : 
                (N341)? bht_q[288] : 
                (N343)? bht_q[291] : 
                (N345)? bht_q[294] : 
                (N347)? bht_q[297] : 
                (N349)? bht_q[300] : 
                (N351)? bht_q[303] : 
                (N353)? bht_q[306] : 
                (N355)? bht_q[309] : 
                (N357)? bht_q[312] : 
                (N359)? bht_q[315] : 
                (N361)? bht_q[318] : 
                (N363)? bht_q[321] : 
                (N365)? bht_q[324] : 
                (N367)? bht_q[327] : 
                (N369)? bht_q[330] : 
                (N371)? bht_q[333] : 
                (N373)? bht_q[336] : 
                (N375)? bht_q[339] : 
                (N377)? bht_q[342] : 
                (N379)? bht_q[345] : 
                (N381)? bht_q[348] : 
                (N383)? bht_q[351] : 
                (N385)? bht_q[354] : 
                (N387)? bht_q[357] : 
                (N389)? bht_q[360] : 
                (N391)? bht_q[363] : 
                (N393)? bht_q[366] : 
                (N395)? bht_q[369] : 
                (N397)? bht_q[372] : 
                (N399)? bht_q[375] : 
                (N401)? bht_q[378] : 
                (N403)? bht_q[381] : 1'b0;
  assign N795 = (N667)? bht_q[1] : 
                (N669)? bht_q[4] : 
                (N671)? bht_q[7] : 
                (N673)? bht_q[10] : 
                (N675)? bht_q[13] : 
                (N677)? bht_q[16] : 
                (N679)? bht_q[19] : 
                (N681)? bht_q[22] : 
                (N683)? bht_q[25] : 
                (N685)? bht_q[28] : 
                (N687)? bht_q[31] : 
                (N689)? bht_q[34] : 
                (N691)? bht_q[37] : 
                (N693)? bht_q[40] : 
                (N695)? bht_q[43] : 
                (N697)? bht_q[46] : 
                (N699)? bht_q[49] : 
                (N701)? bht_q[52] : 
                (N703)? bht_q[55] : 
                (N705)? bht_q[58] : 
                (N707)? bht_q[61] : 
                (N709)? bht_q[64] : 
                (N711)? bht_q[67] : 
                (N713)? bht_q[70] : 
                (N715)? bht_q[73] : 
                (N717)? bht_q[76] : 
                (N719)? bht_q[79] : 
                (N721)? bht_q[82] : 
                (N723)? bht_q[85] : 
                (N725)? bht_q[88] : 
                (N727)? bht_q[91] : 
                (N729)? bht_q[94] : 
                (N731)? bht_q[97] : 
                (N733)? bht_q[100] : 
                (N735)? bht_q[103] : 
                (N737)? bht_q[106] : 
                (N739)? bht_q[109] : 
                (N741)? bht_q[112] : 
                (N743)? bht_q[115] : 
                (N745)? bht_q[118] : 
                (N747)? bht_q[121] : 
                (N749)? bht_q[124] : 
                (N751)? bht_q[127] : 
                (N753)? bht_q[130] : 
                (N755)? bht_q[133] : 
                (N757)? bht_q[136] : 
                (N759)? bht_q[139] : 
                (N761)? bht_q[142] : 
                (N763)? bht_q[145] : 
                (N765)? bht_q[148] : 
                (N767)? bht_q[151] : 
                (N769)? bht_q[154] : 
                (N771)? bht_q[157] : 
                (N773)? bht_q[160] : 
                (N775)? bht_q[163] : 
                (N777)? bht_q[166] : 
                (N779)? bht_q[169] : 
                (N781)? bht_q[172] : 
                (N783)? bht_q[175] : 
                (N785)? bht_q[178] : 
                (N787)? bht_q[181] : 
                (N789)? bht_q[184] : 
                (N791)? bht_q[187] : 
                (N793)? bht_q[190] : 
                (N668)? bht_q[193] : 
                (N670)? bht_q[196] : 
                (N672)? bht_q[199] : 
                (N674)? bht_q[202] : 
                (N676)? bht_q[205] : 
                (N678)? bht_q[208] : 
                (N680)? bht_q[211] : 
                (N682)? bht_q[214] : 
                (N684)? bht_q[217] : 
                (N686)? bht_q[220] : 
                (N688)? bht_q[223] : 
                (N690)? bht_q[226] : 
                (N692)? bht_q[229] : 
                (N694)? bht_q[232] : 
                (N696)? bht_q[235] : 
                (N698)? bht_q[238] : 
                (N700)? bht_q[241] : 
                (N702)? bht_q[244] : 
                (N704)? bht_q[247] : 
                (N706)? bht_q[250] : 
                (N708)? bht_q[253] : 
                (N710)? bht_q[256] : 
                (N712)? bht_q[259] : 
                (N714)? bht_q[262] : 
                (N716)? bht_q[265] : 
                (N718)? bht_q[268] : 
                (N720)? bht_q[271] : 
                (N722)? bht_q[274] : 
                (N724)? bht_q[277] : 
                (N726)? bht_q[280] : 
                (N728)? bht_q[283] : 
                (N730)? bht_q[286] : 
                (N732)? bht_q[289] : 
                (N734)? bht_q[292] : 
                (N736)? bht_q[295] : 
                (N738)? bht_q[298] : 
                (N740)? bht_q[301] : 
                (N742)? bht_q[304] : 
                (N744)? bht_q[307] : 
                (N746)? bht_q[310] : 
                (N748)? bht_q[313] : 
                (N750)? bht_q[316] : 
                (N752)? bht_q[319] : 
                (N754)? bht_q[322] : 
                (N756)? bht_q[325] : 
                (N758)? bht_q[328] : 
                (N760)? bht_q[331] : 
                (N762)? bht_q[334] : 
                (N764)? bht_q[337] : 
                (N766)? bht_q[340] : 
                (N768)? bht_q[343] : 
                (N770)? bht_q[346] : 
                (N772)? bht_q[349] : 
                (N774)? bht_q[352] : 
                (N776)? bht_q[355] : 
                (N778)? bht_q[358] : 
                (N780)? bht_q[361] : 
                (N782)? bht_q[364] : 
                (N784)? bht_q[367] : 
                (N786)? bht_q[370] : 
                (N788)? bht_q[373] : 
                (N790)? bht_q[376] : 
                (N792)? bht_q[379] : 
                (N794)? bht_q[382] : 1'b0;
  assign N796 = (N667)? bht_q[0] : 
                (N669)? bht_q[3] : 
                (N671)? bht_q[6] : 
                (N673)? bht_q[9] : 
                (N675)? bht_q[12] : 
                (N677)? bht_q[15] : 
                (N679)? bht_q[18] : 
                (N681)? bht_q[21] : 
                (N683)? bht_q[24] : 
                (N685)? bht_q[27] : 
                (N687)? bht_q[30] : 
                (N689)? bht_q[33] : 
                (N691)? bht_q[36] : 
                (N693)? bht_q[39] : 
                (N695)? bht_q[42] : 
                (N697)? bht_q[45] : 
                (N699)? bht_q[48] : 
                (N701)? bht_q[51] : 
                (N703)? bht_q[54] : 
                (N705)? bht_q[57] : 
                (N707)? bht_q[60] : 
                (N709)? bht_q[63] : 
                (N711)? bht_q[66] : 
                (N713)? bht_q[69] : 
                (N715)? bht_q[72] : 
                (N717)? bht_q[75] : 
                (N719)? bht_q[78] : 
                (N721)? bht_q[81] : 
                (N723)? bht_q[84] : 
                (N725)? bht_q[87] : 
                (N727)? bht_q[90] : 
                (N729)? bht_q[93] : 
                (N731)? bht_q[96] : 
                (N733)? bht_q[99] : 
                (N735)? bht_q[102] : 
                (N737)? bht_q[105] : 
                (N739)? bht_q[108] : 
                (N741)? bht_q[111] : 
                (N743)? bht_q[114] : 
                (N745)? bht_q[117] : 
                (N747)? bht_q[120] : 
                (N749)? bht_q[123] : 
                (N751)? bht_q[126] : 
                (N753)? bht_q[129] : 
                (N755)? bht_q[132] : 
                (N757)? bht_q[135] : 
                (N759)? bht_q[138] : 
                (N761)? bht_q[141] : 
                (N763)? bht_q[144] : 
                (N765)? bht_q[147] : 
                (N767)? bht_q[150] : 
                (N769)? bht_q[153] : 
                (N771)? bht_q[156] : 
                (N773)? bht_q[159] : 
                (N775)? bht_q[162] : 
                (N777)? bht_q[165] : 
                (N779)? bht_q[168] : 
                (N781)? bht_q[171] : 
                (N783)? bht_q[174] : 
                (N785)? bht_q[177] : 
                (N787)? bht_q[180] : 
                (N789)? bht_q[183] : 
                (N791)? bht_q[186] : 
                (N793)? bht_q[189] : 
                (N668)? bht_q[192] : 
                (N670)? bht_q[195] : 
                (N672)? bht_q[198] : 
                (N674)? bht_q[201] : 
                (N676)? bht_q[204] : 
                (N678)? bht_q[207] : 
                (N680)? bht_q[210] : 
                (N682)? bht_q[213] : 
                (N684)? bht_q[216] : 
                (N686)? bht_q[219] : 
                (N688)? bht_q[222] : 
                (N690)? bht_q[225] : 
                (N692)? bht_q[228] : 
                (N694)? bht_q[231] : 
                (N696)? bht_q[234] : 
                (N698)? bht_q[237] : 
                (N700)? bht_q[240] : 
                (N702)? bht_q[243] : 
                (N704)? bht_q[246] : 
                (N706)? bht_q[249] : 
                (N708)? bht_q[252] : 
                (N710)? bht_q[255] : 
                (N712)? bht_q[258] : 
                (N714)? bht_q[261] : 
                (N716)? bht_q[264] : 
                (N718)? bht_q[267] : 
                (N720)? bht_q[270] : 
                (N722)? bht_q[273] : 
                (N724)? bht_q[276] : 
                (N726)? bht_q[279] : 
                (N728)? bht_q[282] : 
                (N730)? bht_q[285] : 
                (N732)? bht_q[288] : 
                (N734)? bht_q[291] : 
                (N736)? bht_q[294] : 
                (N738)? bht_q[297] : 
                (N740)? bht_q[300] : 
                (N742)? bht_q[303] : 
                (N744)? bht_q[306] : 
                (N746)? bht_q[309] : 
                (N748)? bht_q[312] : 
                (N750)? bht_q[315] : 
                (N752)? bht_q[318] : 
                (N754)? bht_q[321] : 
                (N756)? bht_q[324] : 
                (N758)? bht_q[327] : 
                (N760)? bht_q[330] : 
                (N762)? bht_q[333] : 
                (N764)? bht_q[336] : 
                (N766)? bht_q[339] : 
                (N768)? bht_q[342] : 
                (N770)? bht_q[345] : 
                (N772)? bht_q[348] : 
                (N774)? bht_q[351] : 
                (N776)? bht_q[354] : 
                (N778)? bht_q[357] : 
                (N780)? bht_q[360] : 
                (N782)? bht_q[363] : 
                (N784)? bht_q[366] : 
                (N786)? bht_q[369] : 
                (N788)? bht_q[372] : 
                (N790)? bht_q[375] : 
                (N792)? bht_q[378] : 
                (N794)? bht_q[381] : 1'b0;

  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[383] <= 1'b0;
    end else if(N3130) begin
      bht_q[383] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[382] <= 1'b0;
    end else if(N3132) begin
      bht_q[382] <= N3125;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[381] <= 1'b0;
    end else if(N3134) begin
      bht_q[381] <= N3124;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[380] <= 1'b0;
    end else if(N3139) begin
      bht_q[380] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[379] <= 1'b0;
    end else if(N3140) begin
      bht_q[379] <= N3123;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[378] <= 1'b0;
    end else if(N3140) begin
      bht_q[378] <= N3122;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[377] <= 1'b0;
    end else if(N3143) begin
      bht_q[377] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[376] <= 1'b0;
    end else if(N3140) begin
      bht_q[376] <= N3121;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[375] <= 1'b0;
    end else if(N3140) begin
      bht_q[375] <= N3120;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[374] <= 1'b0;
    end else if(N3146) begin
      bht_q[374] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[373] <= 1'b0;
    end else if(N3140) begin
      bht_q[373] <= N3119;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[372] <= 1'b0;
    end else if(N3140) begin
      bht_q[372] <= N3118;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[371] <= 1'b0;
    end else if(N3149) begin
      bht_q[371] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[370] <= 1'b0;
    end else if(N3140) begin
      bht_q[370] <= N3117;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[369] <= 1'b0;
    end else if(N3140) begin
      bht_q[369] <= N3116;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[368] <= 1'b0;
    end else if(N3152) begin
      bht_q[368] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[367] <= 1'b0;
    end else if(N3140) begin
      bht_q[367] <= N3115;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[366] <= 1'b0;
    end else if(N3140) begin
      bht_q[366] <= N3114;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[365] <= 1'b0;
    end else if(N3155) begin
      bht_q[365] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[364] <= 1'b0;
    end else if(N3140) begin
      bht_q[364] <= N3113;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[363] <= 1'b0;
    end else if(N3140) begin
      bht_q[363] <= N3112;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[362] <= 1'b0;
    end else if(N3158) begin
      bht_q[362] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[361] <= 1'b0;
    end else if(N3140) begin
      bht_q[361] <= N3111;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[360] <= 1'b0;
    end else if(N3140) begin
      bht_q[360] <= N3110;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[359] <= 1'b0;
    end else if(N3161) begin
      bht_q[359] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[358] <= 1'b0;
    end else if(N3140) begin
      bht_q[358] <= N3109;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[357] <= 1'b0;
    end else if(N3140) begin
      bht_q[357] <= N3108;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[356] <= 1'b0;
    end else if(N3164) begin
      bht_q[356] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[355] <= 1'b0;
    end else if(N3140) begin
      bht_q[355] <= N3107;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[354] <= 1'b0;
    end else if(N3140) begin
      bht_q[354] <= N3106;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[353] <= 1'b0;
    end else if(N3167) begin
      bht_q[353] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[352] <= 1'b0;
    end else if(N3140) begin
      bht_q[352] <= N3105;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[351] <= 1'b0;
    end else if(N3140) begin
      bht_q[351] <= N3104;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[350] <= 1'b0;
    end else if(N3170) begin
      bht_q[350] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[349] <= 1'b0;
    end else if(N3140) begin
      bht_q[349] <= N3103;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[348] <= 1'b0;
    end else if(N3140) begin
      bht_q[348] <= N3102;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[347] <= 1'b0;
    end else if(N3173) begin
      bht_q[347] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[346] <= 1'b0;
    end else if(N3140) begin
      bht_q[346] <= N3101;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[345] <= 1'b0;
    end else if(N3140) begin
      bht_q[345] <= N3100;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[344] <= 1'b0;
    end else if(N3176) begin
      bht_q[344] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[343] <= 1'b0;
    end else if(N3140) begin
      bht_q[343] <= N3099;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[342] <= 1'b0;
    end else if(N3140) begin
      bht_q[342] <= N3098;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[341] <= 1'b0;
    end else if(N3179) begin
      bht_q[341] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[340] <= 1'b0;
    end else if(N3140) begin
      bht_q[340] <= N3097;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[339] <= 1'b0;
    end else if(N3140) begin
      bht_q[339] <= N3096;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[338] <= 1'b0;
    end else if(N3182) begin
      bht_q[338] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[337] <= 1'b0;
    end else if(N3140) begin
      bht_q[337] <= N3095;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[336] <= 1'b0;
    end else if(N3140) begin
      bht_q[336] <= N3094;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[335] <= 1'b0;
    end else if(N3185) begin
      bht_q[335] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[334] <= 1'b0;
    end else if(N3140) begin
      bht_q[334] <= N3093;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[333] <= 1'b0;
    end else if(N3140) begin
      bht_q[333] <= N3092;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[332] <= 1'b0;
    end else if(N3188) begin
      bht_q[332] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[331] <= 1'b0;
    end else if(N3140) begin
      bht_q[331] <= N3091;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[330] <= 1'b0;
    end else if(N3140) begin
      bht_q[330] <= N3090;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[329] <= 1'b0;
    end else if(N3191) begin
      bht_q[329] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[328] <= 1'b0;
    end else if(N3140) begin
      bht_q[328] <= N3089;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[327] <= 1'b0;
    end else if(N3140) begin
      bht_q[327] <= N3088;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[326] <= 1'b0;
    end else if(N3194) begin
      bht_q[326] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[325] <= 1'b0;
    end else if(N3140) begin
      bht_q[325] <= N3087;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[324] <= 1'b0;
    end else if(N3140) begin
      bht_q[324] <= N3086;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[323] <= 1'b0;
    end else if(N3197) begin
      bht_q[323] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[322] <= 1'b0;
    end else if(N3140) begin
      bht_q[322] <= N3085;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[321] <= 1'b0;
    end else if(N3140) begin
      bht_q[321] <= N3084;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[320] <= 1'b0;
    end else if(N3200) begin
      bht_q[320] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[319] <= 1'b0;
    end else if(N3140) begin
      bht_q[319] <= N3083;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[318] <= 1'b0;
    end else if(N3140) begin
      bht_q[318] <= N3082;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[317] <= 1'b0;
    end else if(N3203) begin
      bht_q[317] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[316] <= 1'b0;
    end else if(N3140) begin
      bht_q[316] <= N3081;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[315] <= 1'b0;
    end else if(N3140) begin
      bht_q[315] <= N3080;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[314] <= 1'b0;
    end else if(N3206) begin
      bht_q[314] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[313] <= 1'b0;
    end else if(N3140) begin
      bht_q[313] <= N3079;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[312] <= 1'b0;
    end else if(N3140) begin
      bht_q[312] <= N3078;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[311] <= 1'b0;
    end else if(N3209) begin
      bht_q[311] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[310] <= 1'b0;
    end else if(N3140) begin
      bht_q[310] <= N3077;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[309] <= 1'b0;
    end else if(N3140) begin
      bht_q[309] <= N3076;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[308] <= 1'b0;
    end else if(N3212) begin
      bht_q[308] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[307] <= 1'b0;
    end else if(N3140) begin
      bht_q[307] <= N3075;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[306] <= 1'b0;
    end else if(N3140) begin
      bht_q[306] <= N3074;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[305] <= 1'b0;
    end else if(N3215) begin
      bht_q[305] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[304] <= 1'b0;
    end else if(N3140) begin
      bht_q[304] <= N3073;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[303] <= 1'b0;
    end else if(N3140) begin
      bht_q[303] <= N3072;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[302] <= 1'b0;
    end else if(N3218) begin
      bht_q[302] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[301] <= 1'b0;
    end else if(N3140) begin
      bht_q[301] <= N3071;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[300] <= 1'b0;
    end else if(N3140) begin
      bht_q[300] <= N3070;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[299] <= 1'b0;
    end else if(N3221) begin
      bht_q[299] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[298] <= 1'b0;
    end else if(N3140) begin
      bht_q[298] <= N3069;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[297] <= 1'b0;
    end else if(N3140) begin
      bht_q[297] <= N3068;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[296] <= 1'b0;
    end else if(N3224) begin
      bht_q[296] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[295] <= 1'b0;
    end else if(N3134) begin
      bht_q[295] <= N3067;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[294] <= 1'b0;
    end else if(N3134) begin
      bht_q[294] <= N3066;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[293] <= 1'b0;
    end else if(N3227) begin
      bht_q[293] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[292] <= 1'b0;
    end else if(N3134) begin
      bht_q[292] <= N3065;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[291] <= 1'b0;
    end else if(N3134) begin
      bht_q[291] <= N3064;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[290] <= 1'b0;
    end else if(N3230) begin
      bht_q[290] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[289] <= 1'b0;
    end else if(N3134) begin
      bht_q[289] <= N3063;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[288] <= 1'b0;
    end else if(N3134) begin
      bht_q[288] <= N3062;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[287] <= 1'b0;
    end else if(N3233) begin
      bht_q[287] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[286] <= 1'b0;
    end else if(N3134) begin
      bht_q[286] <= N3061;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[285] <= 1'b0;
    end else if(N3134) begin
      bht_q[285] <= N3060;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[284] <= 1'b0;
    end else if(N3236) begin
      bht_q[284] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[283] <= 1'b0;
    end else if(N3134) begin
      bht_q[283] <= N3059;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[282] <= 1'b0;
    end else if(N3134) begin
      bht_q[282] <= N3058;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[281] <= 1'b0;
    end else if(N3239) begin
      bht_q[281] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[280] <= 1'b0;
    end else if(N3134) begin
      bht_q[280] <= N3057;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[279] <= 1'b0;
    end else if(N3134) begin
      bht_q[279] <= N3056;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[278] <= 1'b0;
    end else if(N3242) begin
      bht_q[278] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[277] <= 1'b0;
    end else if(N3134) begin
      bht_q[277] <= N3055;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[276] <= 1'b0;
    end else if(N3134) begin
      bht_q[276] <= N3054;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[275] <= 1'b0;
    end else if(N3245) begin
      bht_q[275] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[274] <= 1'b0;
    end else if(N3134) begin
      bht_q[274] <= N3053;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[273] <= 1'b0;
    end else if(N3134) begin
      bht_q[273] <= N3052;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[272] <= 1'b0;
    end else if(N3248) begin
      bht_q[272] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[271] <= 1'b0;
    end else if(N3134) begin
      bht_q[271] <= N3051;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[270] <= 1'b0;
    end else if(N3134) begin
      bht_q[270] <= N3050;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[269] <= 1'b0;
    end else if(N3251) begin
      bht_q[269] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[268] <= 1'b0;
    end else if(N3134) begin
      bht_q[268] <= N3049;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[267] <= 1'b0;
    end else if(N3134) begin
      bht_q[267] <= N3048;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[266] <= 1'b0;
    end else if(N3254) begin
      bht_q[266] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[265] <= 1'b0;
    end else if(N3134) begin
      bht_q[265] <= N3047;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[264] <= 1'b0;
    end else if(N3134) begin
      bht_q[264] <= N3046;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[263] <= 1'b0;
    end else if(N3257) begin
      bht_q[263] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[262] <= 1'b0;
    end else if(N3134) begin
      bht_q[262] <= N3045;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[261] <= 1'b0;
    end else if(N3134) begin
      bht_q[261] <= N3044;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[260] <= 1'b0;
    end else if(N3260) begin
      bht_q[260] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[259] <= 1'b0;
    end else if(N3134) begin
      bht_q[259] <= N3043;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[258] <= 1'b0;
    end else if(N3134) begin
      bht_q[258] <= N3042;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[257] <= 1'b0;
    end else if(N3263) begin
      bht_q[257] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[256] <= 1'b0;
    end else if(N3134) begin
      bht_q[256] <= N3041;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[255] <= 1'b0;
    end else if(N3134) begin
      bht_q[255] <= N3040;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[254] <= 1'b0;
    end else if(N3266) begin
      bht_q[254] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[253] <= 1'b0;
    end else if(N3134) begin
      bht_q[253] <= N3039;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[252] <= 1'b0;
    end else if(N3134) begin
      bht_q[252] <= N3038;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[251] <= 1'b0;
    end else if(N3269) begin
      bht_q[251] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[250] <= 1'b0;
    end else if(N3134) begin
      bht_q[250] <= N3037;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[249] <= 1'b0;
    end else if(N3134) begin
      bht_q[249] <= N3036;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[248] <= 1'b0;
    end else if(N3272) begin
      bht_q[248] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[247] <= 1'b0;
    end else if(N3134) begin
      bht_q[247] <= N3035;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[246] <= 1'b0;
    end else if(N3134) begin
      bht_q[246] <= N3034;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[245] <= 1'b0;
    end else if(N3275) begin
      bht_q[245] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[244] <= 1'b0;
    end else if(N3134) begin
      bht_q[244] <= N3033;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[243] <= 1'b0;
    end else if(N3134) begin
      bht_q[243] <= N3032;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[242] <= 1'b0;
    end else if(N3278) begin
      bht_q[242] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[241] <= 1'b0;
    end else if(N3134) begin
      bht_q[241] <= N3031;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[240] <= 1'b0;
    end else if(N3134) begin
      bht_q[240] <= N3030;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[239] <= 1'b0;
    end else if(N3281) begin
      bht_q[239] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[238] <= 1'b0;
    end else if(N3134) begin
      bht_q[238] <= N3029;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[237] <= 1'b0;
    end else if(N3134) begin
      bht_q[237] <= N3028;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[236] <= 1'b0;
    end else if(N3284) begin
      bht_q[236] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[235] <= 1'b0;
    end else if(N3134) begin
      bht_q[235] <= N3027;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[234] <= 1'b0;
    end else if(N3134) begin
      bht_q[234] <= N3026;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[233] <= 1'b0;
    end else if(N3287) begin
      bht_q[233] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[232] <= 1'b0;
    end else if(N3134) begin
      bht_q[232] <= N3025;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[231] <= 1'b0;
    end else if(N3134) begin
      bht_q[231] <= N3024;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[230] <= 1'b0;
    end else if(N3290) begin
      bht_q[230] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[229] <= 1'b0;
    end else if(N3134) begin
      bht_q[229] <= N3023;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[228] <= 1'b0;
    end else if(N3134) begin
      bht_q[228] <= N3022;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[227] <= 1'b0;
    end else if(N3293) begin
      bht_q[227] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[226] <= 1'b0;
    end else if(N3134) begin
      bht_q[226] <= N3021;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[225] <= 1'b0;
    end else if(N3134) begin
      bht_q[225] <= N3020;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[224] <= 1'b0;
    end else if(N3296) begin
      bht_q[224] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[223] <= 1'b0;
    end else if(N3134) begin
      bht_q[223] <= N3019;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[222] <= 1'b0;
    end else if(N3134) begin
      bht_q[222] <= N3018;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[221] <= 1'b0;
    end else if(N3299) begin
      bht_q[221] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[220] <= 1'b0;
    end else if(N3134) begin
      bht_q[220] <= N3017;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[219] <= 1'b0;
    end else if(N3134) begin
      bht_q[219] <= N3016;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[218] <= 1'b0;
    end else if(N3302) begin
      bht_q[218] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[217] <= 1'b0;
    end else if(N3134) begin
      bht_q[217] <= N3015;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[216] <= 1'b0;
    end else if(N3134) begin
      bht_q[216] <= N3014;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[215] <= 1'b0;
    end else if(N3305) begin
      bht_q[215] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[214] <= 1'b0;
    end else if(N3134) begin
      bht_q[214] <= N3013;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[213] <= 1'b0;
    end else if(N3134) begin
      bht_q[213] <= N3012;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[212] <= 1'b0;
    end else if(N3308) begin
      bht_q[212] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[211] <= 1'b0;
    end else if(N3134) begin
      bht_q[211] <= N3011;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[210] <= 1'b0;
    end else if(N3134) begin
      bht_q[210] <= N3010;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[209] <= 1'b0;
    end else if(N3311) begin
      bht_q[209] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[208] <= 1'b0;
    end else if(N3134) begin
      bht_q[208] <= N3009;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[207] <= 1'b0;
    end else if(N3134) begin
      bht_q[207] <= N3008;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[206] <= 1'b0;
    end else if(N3314) begin
      bht_q[206] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[205] <= 1'b0;
    end else if(N3134) begin
      bht_q[205] <= N3007;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[204] <= 1'b0;
    end else if(N3134) begin
      bht_q[204] <= N3006;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[203] <= 1'b0;
    end else if(N3317) begin
      bht_q[203] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[202] <= 1'b0;
    end else if(N3134) begin
      bht_q[202] <= N3005;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[201] <= 1'b0;
    end else if(N3134) begin
      bht_q[201] <= N3004;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[200] <= 1'b0;
    end else if(N3320) begin
      bht_q[200] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[199] <= 1'b0;
    end else if(N3134) begin
      bht_q[199] <= N3003;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[198] <= 1'b0;
    end else if(N3134) begin
      bht_q[198] <= N3002;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[197] <= 1'b0;
    end else if(N3323) begin
      bht_q[197] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[196] <= 1'b0;
    end else if(N3132) begin
      bht_q[196] <= N3001;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[195] <= 1'b0;
    end else if(N3132) begin
      bht_q[195] <= N3000;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[194] <= 1'b0;
    end else if(N3326) begin
      bht_q[194] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[193] <= 1'b0;
    end else if(N3132) begin
      bht_q[193] <= N2999;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[192] <= 1'b0;
    end else if(N3132) begin
      bht_q[192] <= N2998;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[191] <= 1'b0;
    end else if(N3329) begin
      bht_q[191] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[190] <= 1'b0;
    end else if(N3132) begin
      bht_q[190] <= N2997;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[189] <= 1'b0;
    end else if(N3132) begin
      bht_q[189] <= N2996;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[188] <= 1'b0;
    end else if(N3332) begin
      bht_q[188] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[187] <= 1'b0;
    end else if(N3132) begin
      bht_q[187] <= N2995;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[186] <= 1'b0;
    end else if(N3132) begin
      bht_q[186] <= N2994;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[185] <= 1'b0;
    end else if(N3335) begin
      bht_q[185] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[184] <= 1'b0;
    end else if(N3132) begin
      bht_q[184] <= N2993;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[183] <= 1'b0;
    end else if(N3132) begin
      bht_q[183] <= N2992;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[182] <= 1'b0;
    end else if(N3338) begin
      bht_q[182] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[181] <= 1'b0;
    end else if(N3132) begin
      bht_q[181] <= N2991;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[180] <= 1'b0;
    end else if(N3132) begin
      bht_q[180] <= N2990;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[179] <= 1'b0;
    end else if(N3341) begin
      bht_q[179] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[178] <= 1'b0;
    end else if(N3132) begin
      bht_q[178] <= N2989;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[177] <= 1'b0;
    end else if(N3132) begin
      bht_q[177] <= N2988;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[176] <= 1'b0;
    end else if(N3344) begin
      bht_q[176] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[175] <= 1'b0;
    end else if(N3132) begin
      bht_q[175] <= N2987;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[174] <= 1'b0;
    end else if(N3132) begin
      bht_q[174] <= N2986;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[173] <= 1'b0;
    end else if(N3347) begin
      bht_q[173] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[172] <= 1'b0;
    end else if(N3132) begin
      bht_q[172] <= N2985;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[171] <= 1'b0;
    end else if(N3132) begin
      bht_q[171] <= N2984;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[170] <= 1'b0;
    end else if(N3350) begin
      bht_q[170] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[169] <= 1'b0;
    end else if(N3132) begin
      bht_q[169] <= N2983;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[168] <= 1'b0;
    end else if(N3132) begin
      bht_q[168] <= N2982;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[167] <= 1'b0;
    end else if(N3353) begin
      bht_q[167] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[166] <= 1'b0;
    end else if(N3132) begin
      bht_q[166] <= N2981;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[165] <= 1'b0;
    end else if(N3132) begin
      bht_q[165] <= N2980;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[164] <= 1'b0;
    end else if(N3356) begin
      bht_q[164] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[163] <= 1'b0;
    end else if(N3132) begin
      bht_q[163] <= N2979;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[162] <= 1'b0;
    end else if(N3132) begin
      bht_q[162] <= N2978;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[161] <= 1'b0;
    end else if(N3359) begin
      bht_q[161] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[160] <= 1'b0;
    end else if(N3132) begin
      bht_q[160] <= N2977;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[159] <= 1'b0;
    end else if(N3132) begin
      bht_q[159] <= N2976;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[158] <= 1'b0;
    end else if(N3362) begin
      bht_q[158] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[157] <= 1'b0;
    end else if(N3132) begin
      bht_q[157] <= N2975;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[156] <= 1'b0;
    end else if(N3132) begin
      bht_q[156] <= N2974;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[155] <= 1'b0;
    end else if(N3365) begin
      bht_q[155] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[154] <= 1'b0;
    end else if(N3132) begin
      bht_q[154] <= N2973;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[153] <= 1'b0;
    end else if(N3132) begin
      bht_q[153] <= N2972;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[152] <= 1'b0;
    end else if(N3368) begin
      bht_q[152] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[151] <= 1'b0;
    end else if(N3132) begin
      bht_q[151] <= N2971;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[150] <= 1'b0;
    end else if(N3132) begin
      bht_q[150] <= N2970;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[149] <= 1'b0;
    end else if(N3371) begin
      bht_q[149] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[148] <= 1'b0;
    end else if(N3132) begin
      bht_q[148] <= N2969;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[147] <= 1'b0;
    end else if(N3132) begin
      bht_q[147] <= N2968;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[146] <= 1'b0;
    end else if(N3374) begin
      bht_q[146] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[145] <= 1'b0;
    end else if(N3132) begin
      bht_q[145] <= N2967;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[144] <= 1'b0;
    end else if(N3132) begin
      bht_q[144] <= N2966;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[143] <= 1'b0;
    end else if(N3377) begin
      bht_q[143] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[142] <= 1'b0;
    end else if(N3132) begin
      bht_q[142] <= N2965;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[141] <= 1'b0;
    end else if(N3132) begin
      bht_q[141] <= N2964;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[140] <= 1'b0;
    end else if(N3380) begin
      bht_q[140] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[139] <= 1'b0;
    end else if(N3132) begin
      bht_q[139] <= N2963;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[138] <= 1'b0;
    end else if(N3132) begin
      bht_q[138] <= N2962;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[137] <= 1'b0;
    end else if(N3383) begin
      bht_q[137] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[136] <= 1'b0;
    end else if(N3132) begin
      bht_q[136] <= N2961;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[135] <= 1'b0;
    end else if(N3132) begin
      bht_q[135] <= N2960;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[134] <= 1'b0;
    end else if(N3386) begin
      bht_q[134] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[133] <= 1'b0;
    end else if(N3132) begin
      bht_q[133] <= N2959;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[132] <= 1'b0;
    end else if(N3132) begin
      bht_q[132] <= N2958;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[131] <= 1'b0;
    end else if(N3389) begin
      bht_q[131] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[130] <= 1'b0;
    end else if(N3132) begin
      bht_q[130] <= N2957;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[129] <= 1'b0;
    end else if(N3132) begin
      bht_q[129] <= N2956;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[128] <= 1'b0;
    end else if(N3392) begin
      bht_q[128] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[127] <= 1'b0;
    end else if(N3132) begin
      bht_q[127] <= N2955;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[126] <= 1'b0;
    end else if(N3132) begin
      bht_q[126] <= N2954;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[125] <= 1'b0;
    end else if(N3395) begin
      bht_q[125] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[124] <= 1'b0;
    end else if(N3132) begin
      bht_q[124] <= N2953;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[123] <= 1'b0;
    end else if(N3132) begin
      bht_q[123] <= N2952;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[122] <= 1'b0;
    end else if(N3398) begin
      bht_q[122] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[121] <= 1'b0;
    end else if(N3132) begin
      bht_q[121] <= N2951;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[120] <= 1'b0;
    end else if(N3132) begin
      bht_q[120] <= N2950;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[119] <= 1'b0;
    end else if(N3401) begin
      bht_q[119] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[118] <= 1'b0;
    end else if(N3132) begin
      bht_q[118] <= N2949;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[117] <= 1'b0;
    end else if(N3132) begin
      bht_q[117] <= N2948;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[116] <= 1'b0;
    end else if(N3404) begin
      bht_q[116] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[115] <= 1'b0;
    end else if(N3132) begin
      bht_q[115] <= N2947;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[114] <= 1'b0;
    end else if(N3132) begin
      bht_q[114] <= N2946;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[113] <= 1'b0;
    end else if(N3407) begin
      bht_q[113] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[112] <= 1'b0;
    end else if(N3132) begin
      bht_q[112] <= N2945;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[111] <= 1'b0;
    end else if(N3132) begin
      bht_q[111] <= N2944;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[110] <= 1'b0;
    end else if(N3410) begin
      bht_q[110] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[109] <= 1'b0;
    end else if(N3132) begin
      bht_q[109] <= N2943;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[108] <= 1'b0;
    end else if(N3132) begin
      bht_q[108] <= N2942;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[107] <= 1'b0;
    end else if(N3413) begin
      bht_q[107] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[106] <= 1'b0;
    end else if(N3132) begin
      bht_q[106] <= N2941;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[105] <= 1'b0;
    end else if(N3132) begin
      bht_q[105] <= N2940;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[104] <= 1'b0;
    end else if(N3416) begin
      bht_q[104] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[103] <= 1'b0;
    end else if(N3132) begin
      bht_q[103] <= N2939;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[102] <= 1'b0;
    end else if(N3132) begin
      bht_q[102] <= N2938;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[101] <= 1'b0;
    end else if(N3419) begin
      bht_q[101] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[100] <= 1'b0;
    end else if(N3132) begin
      bht_q[100] <= N2937;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[99] <= 1'b0;
    end else if(N3132) begin
      bht_q[99] <= N2936;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[98] <= 1'b0;
    end else if(N3422) begin
      bht_q[98] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[97] <= 1'b0;
    end else if(N3423) begin
      bht_q[97] <= N2935;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[96] <= 1'b0;
    end else if(N3423) begin
      bht_q[96] <= N2934;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[95] <= 1'b0;
    end else if(N3426) begin
      bht_q[95] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[94] <= 1'b0;
    end else if(N3423) begin
      bht_q[94] <= N2933;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[93] <= 1'b0;
    end else if(N3423) begin
      bht_q[93] <= N2932;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[92] <= 1'b0;
    end else if(N3429) begin
      bht_q[92] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[91] <= 1'b0;
    end else if(N3423) begin
      bht_q[91] <= N2931;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[90] <= 1'b0;
    end else if(N3423) begin
      bht_q[90] <= N2930;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[89] <= 1'b0;
    end else if(N3432) begin
      bht_q[89] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[88] <= 1'b0;
    end else if(N3423) begin
      bht_q[88] <= N2929;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[87] <= 1'b0;
    end else if(N3423) begin
      bht_q[87] <= N2928;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[86] <= 1'b0;
    end else if(N3435) begin
      bht_q[86] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[85] <= 1'b0;
    end else if(N3423) begin
      bht_q[85] <= N2927;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[84] <= 1'b0;
    end else if(N3423) begin
      bht_q[84] <= N2926;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[83] <= 1'b0;
    end else if(N3438) begin
      bht_q[83] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[82] <= 1'b0;
    end else if(N3423) begin
      bht_q[82] <= N2925;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[81] <= 1'b0;
    end else if(N3423) begin
      bht_q[81] <= N2924;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[80] <= 1'b0;
    end else if(N3441) begin
      bht_q[80] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[79] <= 1'b0;
    end else if(N3423) begin
      bht_q[79] <= N2923;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[78] <= 1'b0;
    end else if(N3423) begin
      bht_q[78] <= N2922;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[77] <= 1'b0;
    end else if(N3444) begin
      bht_q[77] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[76] <= 1'b0;
    end else if(N3423) begin
      bht_q[76] <= N2921;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[75] <= 1'b0;
    end else if(N3423) begin
      bht_q[75] <= N2920;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[74] <= 1'b0;
    end else if(N3447) begin
      bht_q[74] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[73] <= 1'b0;
    end else if(N3423) begin
      bht_q[73] <= N2919;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[72] <= 1'b0;
    end else if(N3423) begin
      bht_q[72] <= N2918;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[71] <= 1'b0;
    end else if(N3450) begin
      bht_q[71] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[70] <= 1'b0;
    end else if(N3423) begin
      bht_q[70] <= N2917;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[69] <= 1'b0;
    end else if(N3423) begin
      bht_q[69] <= N2916;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[68] <= 1'b0;
    end else if(N3453) begin
      bht_q[68] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[67] <= 1'b0;
    end else if(N3423) begin
      bht_q[67] <= N2915;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[66] <= 1'b0;
    end else if(N3423) begin
      bht_q[66] <= N2914;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[65] <= 1'b0;
    end else if(N3456) begin
      bht_q[65] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[64] <= 1'b0;
    end else if(N3423) begin
      bht_q[64] <= N2913;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[63] <= 1'b0;
    end else if(N3423) begin
      bht_q[63] <= N2912;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[62] <= 1'b0;
    end else if(N3459) begin
      bht_q[62] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[61] <= 1'b0;
    end else if(N3423) begin
      bht_q[61] <= N2911;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[60] <= 1'b0;
    end else if(N3423) begin
      bht_q[60] <= N2910;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[59] <= 1'b0;
    end else if(N3462) begin
      bht_q[59] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[58] <= 1'b0;
    end else if(N3423) begin
      bht_q[58] <= N2909;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[57] <= 1'b0;
    end else if(N3423) begin
      bht_q[57] <= N2908;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[56] <= 1'b0;
    end else if(N3465) begin
      bht_q[56] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[55] <= 1'b0;
    end else if(N3423) begin
      bht_q[55] <= N2907;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[54] <= 1'b0;
    end else if(N3423) begin
      bht_q[54] <= N2906;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[53] <= 1'b0;
    end else if(N3468) begin
      bht_q[53] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[52] <= 1'b0;
    end else if(N3423) begin
      bht_q[52] <= N2905;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[51] <= 1'b0;
    end else if(N3423) begin
      bht_q[51] <= N2904;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[50] <= 1'b0;
    end else if(N3471) begin
      bht_q[50] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[49] <= 1'b0;
    end else if(N3423) begin
      bht_q[49] <= N2903;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[48] <= 1'b0;
    end else if(N3423) begin
      bht_q[48] <= N2902;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[47] <= 1'b0;
    end else if(N3474) begin
      bht_q[47] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[46] <= 1'b0;
    end else if(N3423) begin
      bht_q[46] <= N2901;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[45] <= 1'b0;
    end else if(N3423) begin
      bht_q[45] <= N2900;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[44] <= 1'b0;
    end else if(N3477) begin
      bht_q[44] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[43] <= 1'b0;
    end else if(N3423) begin
      bht_q[43] <= N2899;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[42] <= 1'b0;
    end else if(N3423) begin
      bht_q[42] <= N2898;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[41] <= 1'b0;
    end else if(N3480) begin
      bht_q[41] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[40] <= 1'b0;
    end else if(N3423) begin
      bht_q[40] <= N2897;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[39] <= 1'b0;
    end else if(N3423) begin
      bht_q[39] <= N2896;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[38] <= 1'b0;
    end else if(N3483) begin
      bht_q[38] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[37] <= 1'b0;
    end else if(N3423) begin
      bht_q[37] <= N2895;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[36] <= 1'b0;
    end else if(N3423) begin
      bht_q[36] <= N2894;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[35] <= 1'b0;
    end else if(N3486) begin
      bht_q[35] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[34] <= 1'b0;
    end else if(N3423) begin
      bht_q[34] <= N2893;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[33] <= 1'b0;
    end else if(N3423) begin
      bht_q[33] <= N2892;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[32] <= 1'b0;
    end else if(N3489) begin
      bht_q[32] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[31] <= 1'b0;
    end else if(N3423) begin
      bht_q[31] <= N2891;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[30] <= 1'b0;
    end else if(N3423) begin
      bht_q[30] <= N2890;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[29] <= 1'b0;
    end else if(N3492) begin
      bht_q[29] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[28] <= 1'b0;
    end else if(N3423) begin
      bht_q[28] <= N2889;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[27] <= 1'b0;
    end else if(N3423) begin
      bht_q[27] <= N2888;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[26] <= 1'b0;
    end else if(N3495) begin
      bht_q[26] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[25] <= 1'b0;
    end else if(N3423) begin
      bht_q[25] <= N2887;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[24] <= 1'b0;
    end else if(N3423) begin
      bht_q[24] <= N2886;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[23] <= 1'b0;
    end else if(N3498) begin
      bht_q[23] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[22] <= 1'b0;
    end else if(N3423) begin
      bht_q[22] <= N2885;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[21] <= 1'b0;
    end else if(N3423) begin
      bht_q[21] <= N2884;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[20] <= 1'b0;
    end else if(N3501) begin
      bht_q[20] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[19] <= 1'b0;
    end else if(N3423) begin
      bht_q[19] <= N2883;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[18] <= 1'b0;
    end else if(N3423) begin
      bht_q[18] <= N2882;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[17] <= 1'b0;
    end else if(N3504) begin
      bht_q[17] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[16] <= 1'b0;
    end else if(N3423) begin
      bht_q[16] <= N2881;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[15] <= 1'b0;
    end else if(N3423) begin
      bht_q[15] <= N2880;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[14] <= 1'b0;
    end else if(N3507) begin
      bht_q[14] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[13] <= 1'b0;
    end else if(N3423) begin
      bht_q[13] <= N2879;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[12] <= 1'b0;
    end else if(N3423) begin
      bht_q[12] <= N2878;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[11] <= 1'b0;
    end else if(N3510) begin
      bht_q[11] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[10] <= 1'b0;
    end else if(N3423) begin
      bht_q[10] <= N2877;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[9] <= 1'b0;
    end else if(N3423) begin
      bht_q[9] <= N2876;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[8] <= 1'b0;
    end else if(N3513) begin
      bht_q[8] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[7] <= 1'b0;
    end else if(N3423) begin
      bht_q[7] <= N2875;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[6] <= 1'b0;
    end else if(N3423) begin
      bht_q[6] <= N2874;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[5] <= 1'b0;
    end else if(N3516) begin
      bht_q[5] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[4] <= 1'b0;
    end else if(N3423) begin
      bht_q[4] <= N2873;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[3] <= 1'b0;
    end else if(N3423) begin
      bht_q[3] <= N2872;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[2] <= 1'b0;
    end else if(N3519) begin
      bht_q[2] <= N2869;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[1] <= 1'b0;
    end else if(N3423) begin
      bht_q[1] <= N2871;
    end 
  end


  always @(posedge clk_i or posedge N2868) begin
    if(N2868) begin
      bht_q[0] <= 1'b0;
    end else if(N3423) begin
      bht_q[0] <= N2870;
    end 
  end

  assign N3520 = ~N468;
  assign N3521 = N469 | N3520;
  assign bht_prediction_o_taken_ = ~N3521;
  assign bht_prediction_o_strongly_taken_ = N535 & N534;
  assign N3524 = N796 & N795;
  assign N3525 = N796 | N795;
  assign N3526 = ~N3525;
  assign { N1062, N1061 } = { N795, N796 } - 1'b1;
  assign { N1578, N1577 } = { N795, N796 } + 1'b1;
  assign { N2351, N2350 } = { N795, N796 } - 1'b1;
  assign { N2093, N2092 } = { N795, N796 } + 1'b1;
  assign N3527 = ~bht_update_i[10];
  assign N3528 = bht_update_i[8] & bht_update_i[9];
  assign N3529 = N0 & bht_update_i[9];
  assign N0 = ~bht_update_i[8];
  assign N3530 = bht_update_i[8] & N1;
  assign N1 = ~bht_update_i[9];
  assign N3531 = N2 & N3;
  assign N2 = ~bht_update_i[8];
  assign N3 = ~bht_update_i[9];
  assign N3532 = bht_update_i[10] & N3528;
  assign N3533 = bht_update_i[10] & N3529;
  assign N3534 = bht_update_i[10] & N3530;
  assign N3535 = bht_update_i[10] & N3531;
  assign N3536 = N3527 & N3528;
  assign N3537 = N3527 & N3529;
  assign N3538 = N3527 & N3530;
  assign N3539 = N3527 & N3531;
  assign N3540 = bht_update_i[6] & bht_update_i[7];
  assign N3541 = N4 & bht_update_i[7];
  assign N4 = ~bht_update_i[6];
  assign N3542 = bht_update_i[6] & N5;
  assign N5 = ~bht_update_i[7];
  assign N3543 = N6 & N7;
  assign N6 = ~bht_update_i[6];
  assign N7 = ~bht_update_i[7];
  assign N3544 = bht_update_i[4] & bht_update_i[5];
  assign N3545 = N8 & bht_update_i[5];
  assign N8 = ~bht_update_i[4];
  assign N3546 = bht_update_i[4] & N9;
  assign N9 = ~bht_update_i[5];
  assign N3547 = N10 & N11;
  assign N10 = ~bht_update_i[4];
  assign N11 = ~bht_update_i[5];
  assign N3548 = N3540 & N3544;
  assign N3549 = N3540 & N3545;
  assign N3550 = N3540 & N3546;
  assign N3551 = N3540 & N3547;
  assign N3552 = N3541 & N3544;
  assign N3553 = N3541 & N3545;
  assign N3554 = N3541 & N3546;
  assign N3555 = N3541 & N3547;
  assign N3556 = N3542 & N3544;
  assign N3557 = N3542 & N3545;
  assign N3558 = N3542 & N3546;
  assign N3559 = N3542 & N3547;
  assign N3560 = N3543 & N3544;
  assign N3561 = N3543 & N3545;
  assign N3562 = N3543 & N3546;
  assign N3563 = N3543 & N3547;
  assign N927 = N3532 & N3548;
  assign N926 = N3532 & N3549;
  assign N925 = N3532 & N3550;
  assign N924 = N3532 & N3551;
  assign N923 = N3532 & N3552;
  assign N922 = N3532 & N3553;
  assign N921 = N3532 & N3554;
  assign N920 = N3532 & N3555;
  assign N919 = N3532 & N3556;
  assign N918 = N3532 & N3557;
  assign N917 = N3532 & N3558;
  assign N916 = N3532 & N3559;
  assign N915 = N3532 & N3560;
  assign N914 = N3532 & N3561;
  assign N913 = N3532 & N3562;
  assign N912 = N3532 & N3563;
  assign N911 = N3533 & N3548;
  assign N910 = N3533 & N3549;
  assign N909 = N3533 & N3550;
  assign N908 = N3533 & N3551;
  assign N907 = N3533 & N3552;
  assign N906 = N3533 & N3553;
  assign N905 = N3533 & N3554;
  assign N904 = N3533 & N3555;
  assign N903 = N3533 & N3556;
  assign N902 = N3533 & N3557;
  assign N901 = N3533 & N3558;
  assign N900 = N3533 & N3559;
  assign N899 = N3533 & N3560;
  assign N898 = N3533 & N3561;
  assign N897 = N3533 & N3562;
  assign N896 = N3533 & N3563;
  assign N895 = N3534 & N3548;
  assign N894 = N3534 & N3549;
  assign N893 = N3534 & N3550;
  assign N892 = N3534 & N3551;
  assign N891 = N3534 & N3552;
  assign N890 = N3534 & N3553;
  assign N889 = N3534 & N3554;
  assign N888 = N3534 & N3555;
  assign N887 = N3534 & N3556;
  assign N886 = N3534 & N3557;
  assign N885 = N3534 & N3558;
  assign N884 = N3534 & N3559;
  assign N883 = N3534 & N3560;
  assign N882 = N3534 & N3561;
  assign N881 = N3534 & N3562;
  assign N880 = N3534 & N3563;
  assign N879 = N3535 & N3548;
  assign N878 = N3535 & N3549;
  assign N877 = N3535 & N3550;
  assign N876 = N3535 & N3551;
  assign N875 = N3535 & N3552;
  assign N874 = N3535 & N3553;
  assign N873 = N3535 & N3554;
  assign N872 = N3535 & N3555;
  assign N871 = N3535 & N3556;
  assign N870 = N3535 & N3557;
  assign N869 = N3535 & N3558;
  assign N868 = N3535 & N3559;
  assign N867 = N3535 & N3560;
  assign N866 = N3535 & N3561;
  assign N865 = N3535 & N3562;
  assign N864 = N3535 & N3563;
  assign N863 = N3536 & N3548;
  assign N862 = N3536 & N3549;
  assign N861 = N3536 & N3550;
  assign N860 = N3536 & N3551;
  assign N859 = N3536 & N3552;
  assign N858 = N3536 & N3553;
  assign N857 = N3536 & N3554;
  assign N856 = N3536 & N3555;
  assign N855 = N3536 & N3556;
  assign N854 = N3536 & N3557;
  assign N853 = N3536 & N3558;
  assign N852 = N3536 & N3559;
  assign N851 = N3536 & N3560;
  assign N850 = N3536 & N3561;
  assign N849 = N3536 & N3562;
  assign N848 = N3536 & N3563;
  assign N847 = N3537 & N3548;
  assign N846 = N3537 & N3549;
  assign N845 = N3537 & N3550;
  assign N844 = N3537 & N3551;
  assign N843 = N3537 & N3552;
  assign N842 = N3537 & N3553;
  assign N841 = N3537 & N3554;
  assign N840 = N3537 & N3555;
  assign N839 = N3537 & N3556;
  assign N838 = N3537 & N3557;
  assign N837 = N3537 & N3558;
  assign N836 = N3537 & N3559;
  assign N835 = N3537 & N3560;
  assign N834 = N3537 & N3561;
  assign N833 = N3537 & N3562;
  assign N832 = N3537 & N3563;
  assign N831 = N3538 & N3548;
  assign N830 = N3538 & N3549;
  assign N829 = N3538 & N3550;
  assign N828 = N3538 & N3551;
  assign N827 = N3538 & N3552;
  assign N826 = N3538 & N3553;
  assign N825 = N3538 & N3554;
  assign N824 = N3538 & N3555;
  assign N823 = N3538 & N3556;
  assign N822 = N3538 & N3557;
  assign N821 = N3538 & N3558;
  assign N820 = N3538 & N3559;
  assign N819 = N3538 & N3560;
  assign N818 = N3538 & N3561;
  assign N817 = N3538 & N3562;
  assign N816 = N3538 & N3563;
  assign N815 = N3539 & N3548;
  assign N814 = N3539 & N3549;
  assign N813 = N3539 & N3550;
  assign N812 = N3539 & N3551;
  assign N811 = N3539 & N3552;
  assign N810 = N3539 & N3553;
  assign N809 = N3539 & N3554;
  assign N808 = N3539 & N3555;
  assign N807 = N3539 & N3556;
  assign N806 = N3539 & N3557;
  assign N805 = N3539 & N3558;
  assign N804 = N3539 & N3559;
  assign N803 = N3539 & N3560;
  assign N802 = N3539 & N3561;
  assign N801 = N3539 & N3562;
  assign N800 = N3539 & N3563;
  assign { N1064, N1063 } = (N12)? { N1062, N1061 } : 
                            (N928)? bht_q[1:0] : 1'b0;
  assign N12 = N800;
  assign { N1066, N1065 } = (N13)? { N1062, N1061 } : 
                            (N929)? bht_q[4:3] : 1'b0;
  assign N13 = N801;
  assign { N1068, N1067 } = (N14)? { N1062, N1061 } : 
                            (N930)? bht_q[7:6] : 1'b0;
  assign N14 = N802;
  assign { N1070, N1069 } = (N15)? { N1062, N1061 } : 
                            (N931)? bht_q[10:9] : 1'b0;
  assign N15 = N803;
  assign { N1072, N1071 } = (N16)? { N1062, N1061 } : 
                            (N932)? bht_q[13:12] : 1'b0;
  assign N16 = N804;
  assign { N1074, N1073 } = (N17)? { N1062, N1061 } : 
                            (N933)? bht_q[16:15] : 1'b0;
  assign N17 = N805;
  assign { N1076, N1075 } = (N18)? { N1062, N1061 } : 
                            (N934)? bht_q[19:18] : 1'b0;
  assign N18 = N806;
  assign { N1078, N1077 } = (N19)? { N1062, N1061 } : 
                            (N935)? bht_q[22:21] : 1'b0;
  assign N19 = N807;
  assign { N1080, N1079 } = (N20)? { N1062, N1061 } : 
                            (N936)? bht_q[25:24] : 1'b0;
  assign N20 = N808;
  assign { N1082, N1081 } = (N21)? { N1062, N1061 } : 
                            (N937)? bht_q[28:27] : 1'b0;
  assign N21 = N809;
  assign { N1084, N1083 } = (N22)? { N1062, N1061 } : 
                            (N938)? bht_q[31:30] : 1'b0;
  assign N22 = N810;
  assign { N1086, N1085 } = (N23)? { N1062, N1061 } : 
                            (N939)? bht_q[34:33] : 1'b0;
  assign N23 = N811;
  assign { N1088, N1087 } = (N24)? { N1062, N1061 } : 
                            (N940)? bht_q[37:36] : 1'b0;
  assign N24 = N812;
  assign { N1090, N1089 } = (N25)? { N1062, N1061 } : 
                            (N941)? bht_q[40:39] : 1'b0;
  assign N25 = N813;
  assign { N1092, N1091 } = (N26)? { N1062, N1061 } : 
                            (N942)? bht_q[43:42] : 1'b0;
  assign N26 = N814;
  assign { N1094, N1093 } = (N27)? { N1062, N1061 } : 
                            (N943)? bht_q[46:45] : 1'b0;
  assign N27 = N815;
  assign { N1096, N1095 } = (N28)? { N1062, N1061 } : 
                            (N944)? bht_q[49:48] : 1'b0;
  assign N28 = N816;
  assign { N1098, N1097 } = (N29)? { N1062, N1061 } : 
                            (N945)? bht_q[52:51] : 1'b0;
  assign N29 = N817;
  assign { N1100, N1099 } = (N30)? { N1062, N1061 } : 
                            (N946)? bht_q[55:54] : 1'b0;
  assign N30 = N818;
  assign { N1102, N1101 } = (N31)? { N1062, N1061 } : 
                            (N947)? bht_q[58:57] : 1'b0;
  assign N31 = N819;
  assign { N1104, N1103 } = (N32)? { N1062, N1061 } : 
                            (N948)? bht_q[61:60] : 1'b0;
  assign N32 = N820;
  assign { N1106, N1105 } = (N33)? { N1062, N1061 } : 
                            (N949)? bht_q[64:63] : 1'b0;
  assign N33 = N821;
  assign { N1108, N1107 } = (N34)? { N1062, N1061 } : 
                            (N950)? bht_q[67:66] : 1'b0;
  assign N34 = N822;
  assign { N1110, N1109 } = (N35)? { N1062, N1061 } : 
                            (N951)? bht_q[70:69] : 1'b0;
  assign N35 = N823;
  assign { N1112, N1111 } = (N36)? { N1062, N1061 } : 
                            (N952)? bht_q[73:72] : 1'b0;
  assign N36 = N824;
  assign { N1114, N1113 } = (N37)? { N1062, N1061 } : 
                            (N953)? bht_q[76:75] : 1'b0;
  assign N37 = N825;
  assign { N1116, N1115 } = (N38)? { N1062, N1061 } : 
                            (N954)? bht_q[79:78] : 1'b0;
  assign N38 = N826;
  assign { N1118, N1117 } = (N39)? { N1062, N1061 } : 
                            (N955)? bht_q[82:81] : 1'b0;
  assign N39 = N827;
  assign { N1120, N1119 } = (N40)? { N1062, N1061 } : 
                            (N956)? bht_q[85:84] : 1'b0;
  assign N40 = N828;
  assign { N1122, N1121 } = (N41)? { N1062, N1061 } : 
                            (N957)? bht_q[88:87] : 1'b0;
  assign N41 = N829;
  assign { N1124, N1123 } = (N42)? { N1062, N1061 } : 
                            (N958)? bht_q[91:90] : 1'b0;
  assign N42 = N830;
  assign { N1126, N1125 } = (N43)? { N1062, N1061 } : 
                            (N959)? bht_q[94:93] : 1'b0;
  assign N43 = N831;
  assign { N1128, N1127 } = (N44)? { N1062, N1061 } : 
                            (N960)? bht_q[97:96] : 1'b0;
  assign N44 = N832;
  assign { N1130, N1129 } = (N45)? { N1062, N1061 } : 
                            (N961)? bht_q[100:99] : 1'b0;
  assign N45 = N833;
  assign { N1132, N1131 } = (N46)? { N1062, N1061 } : 
                            (N962)? bht_q[103:102] : 1'b0;
  assign N46 = N834;
  assign { N1134, N1133 } = (N47)? { N1062, N1061 } : 
                            (N963)? bht_q[106:105] : 1'b0;
  assign N47 = N835;
  assign { N1136, N1135 } = (N48)? { N1062, N1061 } : 
                            (N964)? bht_q[109:108] : 1'b0;
  assign N48 = N836;
  assign { N1138, N1137 } = (N49)? { N1062, N1061 } : 
                            (N965)? bht_q[112:111] : 1'b0;
  assign N49 = N837;
  assign { N1140, N1139 } = (N50)? { N1062, N1061 } : 
                            (N966)? bht_q[115:114] : 1'b0;
  assign N50 = N838;
  assign { N1142, N1141 } = (N51)? { N1062, N1061 } : 
                            (N967)? bht_q[118:117] : 1'b0;
  assign N51 = N839;
  assign { N1144, N1143 } = (N52)? { N1062, N1061 } : 
                            (N968)? bht_q[121:120] : 1'b0;
  assign N52 = N840;
  assign { N1146, N1145 } = (N53)? { N1062, N1061 } : 
                            (N969)? bht_q[124:123] : 1'b0;
  assign N53 = N841;
  assign { N1148, N1147 } = (N54)? { N1062, N1061 } : 
                            (N970)? bht_q[127:126] : 1'b0;
  assign N54 = N842;
  assign { N1150, N1149 } = (N55)? { N1062, N1061 } : 
                            (N971)? bht_q[130:129] : 1'b0;
  assign N55 = N843;
  assign { N1152, N1151 } = (N56)? { N1062, N1061 } : 
                            (N972)? bht_q[133:132] : 1'b0;
  assign N56 = N844;
  assign { N1154, N1153 } = (N57)? { N1062, N1061 } : 
                            (N973)? bht_q[136:135] : 1'b0;
  assign N57 = N845;
  assign { N1156, N1155 } = (N58)? { N1062, N1061 } : 
                            (N974)? bht_q[139:138] : 1'b0;
  assign N58 = N846;
  assign { N1158, N1157 } = (N59)? { N1062, N1061 } : 
                            (N975)? bht_q[142:141] : 1'b0;
  assign N59 = N847;
  assign { N1160, N1159 } = (N60)? { N1062, N1061 } : 
                            (N976)? bht_q[145:144] : 1'b0;
  assign N60 = N848;
  assign { N1162, N1161 } = (N61)? { N1062, N1061 } : 
                            (N977)? bht_q[148:147] : 1'b0;
  assign N61 = N849;
  assign { N1164, N1163 } = (N62)? { N1062, N1061 } : 
                            (N978)? bht_q[151:150] : 1'b0;
  assign N62 = N850;
  assign { N1166, N1165 } = (N63)? { N1062, N1061 } : 
                            (N979)? bht_q[154:153] : 1'b0;
  assign N63 = N851;
  assign { N1168, N1167 } = (N64)? { N1062, N1061 } : 
                            (N980)? bht_q[157:156] : 1'b0;
  assign N64 = N852;
  assign { N1170, N1169 } = (N65)? { N1062, N1061 } : 
                            (N981)? bht_q[160:159] : 1'b0;
  assign N65 = N853;
  assign { N1172, N1171 } = (N66)? { N1062, N1061 } : 
                            (N982)? bht_q[163:162] : 1'b0;
  assign N66 = N854;
  assign { N1174, N1173 } = (N67)? { N1062, N1061 } : 
                            (N983)? bht_q[166:165] : 1'b0;
  assign N67 = N855;
  assign { N1176, N1175 } = (N68)? { N1062, N1061 } : 
                            (N984)? bht_q[169:168] : 1'b0;
  assign N68 = N856;
  assign { N1178, N1177 } = (N69)? { N1062, N1061 } : 
                            (N985)? bht_q[172:171] : 1'b0;
  assign N69 = N857;
  assign { N1180, N1179 } = (N70)? { N1062, N1061 } : 
                            (N986)? bht_q[175:174] : 1'b0;
  assign N70 = N858;
  assign { N1182, N1181 } = (N71)? { N1062, N1061 } : 
                            (N987)? bht_q[178:177] : 1'b0;
  assign N71 = N859;
  assign { N1184, N1183 } = (N72)? { N1062, N1061 } : 
                            (N988)? bht_q[181:180] : 1'b0;
  assign N72 = N860;
  assign { N1186, N1185 } = (N73)? { N1062, N1061 } : 
                            (N989)? bht_q[184:183] : 1'b0;
  assign N73 = N861;
  assign { N1188, N1187 } = (N74)? { N1062, N1061 } : 
                            (N990)? bht_q[187:186] : 1'b0;
  assign N74 = N862;
  assign { N1190, N1189 } = (N75)? { N1062, N1061 } : 
                            (N991)? bht_q[190:189] : 1'b0;
  assign N75 = N863;
  assign { N1192, N1191 } = (N76)? { N1062, N1061 } : 
                            (N992)? bht_q[193:192] : 1'b0;
  assign N76 = N864;
  assign { N1194, N1193 } = (N77)? { N1062, N1061 } : 
                            (N993)? bht_q[196:195] : 1'b0;
  assign N77 = N865;
  assign { N1196, N1195 } = (N78)? { N1062, N1061 } : 
                            (N994)? bht_q[199:198] : 1'b0;
  assign N78 = N866;
  assign { N1198, N1197 } = (N79)? { N1062, N1061 } : 
                            (N995)? bht_q[202:201] : 1'b0;
  assign N79 = N867;
  assign { N1200, N1199 } = (N80)? { N1062, N1061 } : 
                            (N996)? bht_q[205:204] : 1'b0;
  assign N80 = N868;
  assign { N1202, N1201 } = (N81)? { N1062, N1061 } : 
                            (N997)? bht_q[208:207] : 1'b0;
  assign N81 = N869;
  assign { N1204, N1203 } = (N82)? { N1062, N1061 } : 
                            (N998)? bht_q[211:210] : 1'b0;
  assign N82 = N870;
  assign { N1206, N1205 } = (N83)? { N1062, N1061 } : 
                            (N999)? bht_q[214:213] : 1'b0;
  assign N83 = N871;
  assign { N1208, N1207 } = (N84)? { N1062, N1061 } : 
                            (N1000)? bht_q[217:216] : 1'b0;
  assign N84 = N872;
  assign { N1210, N1209 } = (N85)? { N1062, N1061 } : 
                            (N1001)? bht_q[220:219] : 1'b0;
  assign N85 = N873;
  assign { N1212, N1211 } = (N86)? { N1062, N1061 } : 
                            (N1002)? bht_q[223:222] : 1'b0;
  assign N86 = N874;
  assign { N1214, N1213 } = (N87)? { N1062, N1061 } : 
                            (N1003)? bht_q[226:225] : 1'b0;
  assign N87 = N875;
  assign { N1216, N1215 } = (N88)? { N1062, N1061 } : 
                            (N1004)? bht_q[229:228] : 1'b0;
  assign N88 = N876;
  assign { N1218, N1217 } = (N89)? { N1062, N1061 } : 
                            (N1005)? bht_q[232:231] : 1'b0;
  assign N89 = N877;
  assign { N1220, N1219 } = (N90)? { N1062, N1061 } : 
                            (N1006)? bht_q[235:234] : 1'b0;
  assign N90 = N878;
  assign { N1222, N1221 } = (N91)? { N1062, N1061 } : 
                            (N1007)? bht_q[238:237] : 1'b0;
  assign N91 = N879;
  assign { N1224, N1223 } = (N92)? { N1062, N1061 } : 
                            (N1008)? bht_q[241:240] : 1'b0;
  assign N92 = N880;
  assign { N1226, N1225 } = (N93)? { N1062, N1061 } : 
                            (N1009)? bht_q[244:243] : 1'b0;
  assign N93 = N881;
  assign { N1228, N1227 } = (N94)? { N1062, N1061 } : 
                            (N1010)? bht_q[247:246] : 1'b0;
  assign N94 = N882;
  assign { N1230, N1229 } = (N95)? { N1062, N1061 } : 
                            (N1011)? bht_q[250:249] : 1'b0;
  assign N95 = N883;
  assign { N1232, N1231 } = (N96)? { N1062, N1061 } : 
                            (N1012)? bht_q[253:252] : 1'b0;
  assign N96 = N884;
  assign { N1234, N1233 } = (N97)? { N1062, N1061 } : 
                            (N1013)? bht_q[256:255] : 1'b0;
  assign N97 = N885;
  assign { N1236, N1235 } = (N98)? { N1062, N1061 } : 
                            (N1014)? bht_q[259:258] : 1'b0;
  assign N98 = N886;
  assign { N1238, N1237 } = (N99)? { N1062, N1061 } : 
                            (N1015)? bht_q[262:261] : 1'b0;
  assign N99 = N887;
  assign { N1240, N1239 } = (N100)? { N1062, N1061 } : 
                            (N1016)? bht_q[265:264] : 1'b0;
  assign N100 = N888;
  assign { N1242, N1241 } = (N101)? { N1062, N1061 } : 
                            (N1017)? bht_q[268:267] : 1'b0;
  assign N101 = N889;
  assign { N1244, N1243 } = (N102)? { N1062, N1061 } : 
                            (N1018)? bht_q[271:270] : 1'b0;
  assign N102 = N890;
  assign { N1246, N1245 } = (N103)? { N1062, N1061 } : 
                            (N1019)? bht_q[274:273] : 1'b0;
  assign N103 = N891;
  assign { N1248, N1247 } = (N104)? { N1062, N1061 } : 
                            (N1020)? bht_q[277:276] : 1'b0;
  assign N104 = N892;
  assign { N1250, N1249 } = (N105)? { N1062, N1061 } : 
                            (N1021)? bht_q[280:279] : 1'b0;
  assign N105 = N893;
  assign { N1252, N1251 } = (N106)? { N1062, N1061 } : 
                            (N1022)? bht_q[283:282] : 1'b0;
  assign N106 = N894;
  assign { N1254, N1253 } = (N107)? { N1062, N1061 } : 
                            (N1023)? bht_q[286:285] : 1'b0;
  assign N107 = N895;
  assign { N1256, N1255 } = (N108)? { N1062, N1061 } : 
                            (N1024)? bht_q[289:288] : 1'b0;
  assign N108 = N896;
  assign { N1258, N1257 } = (N109)? { N1062, N1061 } : 
                            (N1025)? bht_q[292:291] : 1'b0;
  assign N109 = N897;
  assign { N1260, N1259 } = (N110)? { N1062, N1061 } : 
                            (N1026)? bht_q[295:294] : 1'b0;
  assign N110 = N898;
  assign { N1262, N1261 } = (N111)? { N1062, N1061 } : 
                            (N1027)? bht_q[298:297] : 1'b0;
  assign N111 = N899;
  assign { N1264, N1263 } = (N112)? { N1062, N1061 } : 
                            (N1028)? bht_q[301:300] : 1'b0;
  assign N112 = N900;
  assign { N1266, N1265 } = (N113)? { N1062, N1061 } : 
                            (N1029)? bht_q[304:303] : 1'b0;
  assign N113 = N901;
  assign { N1268, N1267 } = (N114)? { N1062, N1061 } : 
                            (N1030)? bht_q[307:306] : 1'b0;
  assign N114 = N902;
  assign { N1270, N1269 } = (N115)? { N1062, N1061 } : 
                            (N1031)? bht_q[310:309] : 1'b0;
  assign N115 = N903;
  assign { N1272, N1271 } = (N116)? { N1062, N1061 } : 
                            (N1032)? bht_q[313:312] : 1'b0;
  assign N116 = N904;
  assign { N1274, N1273 } = (N117)? { N1062, N1061 } : 
                            (N1033)? bht_q[316:315] : 1'b0;
  assign N117 = N905;
  assign { N1276, N1275 } = (N118)? { N1062, N1061 } : 
                            (N1034)? bht_q[319:318] : 1'b0;
  assign N118 = N906;
  assign { N1278, N1277 } = (N119)? { N1062, N1061 } : 
                            (N1035)? bht_q[322:321] : 1'b0;
  assign N119 = N907;
  assign { N1280, N1279 } = (N120)? { N1062, N1061 } : 
                            (N1036)? bht_q[325:324] : 1'b0;
  assign N120 = N908;
  assign { N1282, N1281 } = (N121)? { N1062, N1061 } : 
                            (N1037)? bht_q[328:327] : 1'b0;
  assign N121 = N909;
  assign { N1284, N1283 } = (N122)? { N1062, N1061 } : 
                            (N1038)? bht_q[331:330] : 1'b0;
  assign N122 = N910;
  assign { N1286, N1285 } = (N123)? { N1062, N1061 } : 
                            (N1039)? bht_q[334:333] : 1'b0;
  assign N123 = N911;
  assign { N1288, N1287 } = (N124)? { N1062, N1061 } : 
                            (N1040)? bht_q[337:336] : 1'b0;
  assign N124 = N912;
  assign { N1290, N1289 } = (N125)? { N1062, N1061 } : 
                            (N1041)? bht_q[340:339] : 1'b0;
  assign N125 = N913;
  assign { N1292, N1291 } = (N126)? { N1062, N1061 } : 
                            (N1042)? bht_q[343:342] : 1'b0;
  assign N126 = N914;
  assign { N1294, N1293 } = (N127)? { N1062, N1061 } : 
                            (N1043)? bht_q[346:345] : 1'b0;
  assign N127 = N915;
  assign { N1296, N1295 } = (N128)? { N1062, N1061 } : 
                            (N1044)? bht_q[349:348] : 1'b0;
  assign N128 = N916;
  assign { N1298, N1297 } = (N129)? { N1062, N1061 } : 
                            (N1045)? bht_q[352:351] : 1'b0;
  assign N129 = N917;
  assign { N1300, N1299 } = (N130)? { N1062, N1061 } : 
                            (N1046)? bht_q[355:354] : 1'b0;
  assign N130 = N918;
  assign { N1302, N1301 } = (N131)? { N1062, N1061 } : 
                            (N1047)? bht_q[358:357] : 1'b0;
  assign N131 = N919;
  assign { N1304, N1303 } = (N132)? { N1062, N1061 } : 
                            (N1048)? bht_q[361:360] : 1'b0;
  assign N132 = N920;
  assign { N1306, N1305 } = (N133)? { N1062, N1061 } : 
                            (N1049)? bht_q[364:363] : 1'b0;
  assign N133 = N921;
  assign { N1308, N1307 } = (N134)? { N1062, N1061 } : 
                            (N1050)? bht_q[367:366] : 1'b0;
  assign N134 = N922;
  assign { N1310, N1309 } = (N135)? { N1062, N1061 } : 
                            (N1051)? bht_q[370:369] : 1'b0;
  assign N135 = N923;
  assign { N1312, N1311 } = (N136)? { N1062, N1061 } : 
                            (N1052)? bht_q[373:372] : 1'b0;
  assign N136 = N924;
  assign { N1314, N1313 } = (N137)? { N1062, N1061 } : 
                            (N1053)? bht_q[376:375] : 1'b0;
  assign N137 = N925;
  assign { N1316, N1315 } = (N138)? { N1062, N1061 } : 
                            (N1054)? bht_q[379:378] : 1'b0;
  assign N138 = N926;
  assign { N1318, N1317 } = (N139)? { N1062, N1061 } : 
                            (N1055)? bht_q[382:381] : 1'b0;
  assign N139 = N927;
  assign { N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319 } = (N140)? { N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N141)? { bht_q[382:381], bht_q[379:378], bht_q[376:375], bht_q[373:372], bht_q[370:369], bht_q[367:366], bht_q[364:363], bht_q[361:360], bht_q[358:357], bht_q[355:354], bht_q[352:351], bht_q[349:348], bht_q[346:345], bht_q[343:342], bht_q[340:339], bht_q[337:336], bht_q[334:333], bht_q[331:330], bht_q[328:327], bht_q[325:324], bht_q[322:321], bht_q[319:318], bht_q[316:315], bht_q[313:312], bht_q[310:309], bht_q[307:306], bht_q[304:303], bht_q[301:300], bht_q[298:297], bht_q[295:294], bht_q[292:291], bht_q[289:288], bht_q[286:285], bht_q[283:282], bht_q[280:279], bht_q[277:276], bht_q[274:273], bht_q[271:270], bht_q[268:267], bht_q[265:264], bht_q[262:261], bht_q[259:258], bht_q[256:255], bht_q[253:252], bht_q[250:249], bht_q[247:246], bht_q[244:243], bht_q[241:240], bht_q[238:237], bht_q[235:234], bht_q[232:231], bht_q[229:228], bht_q[226:225], bht_q[223:222], bht_q[220:219], bht_q[217:216], bht_q[214:213], bht_q[211:210], bht_q[208:207], bht_q[205:204], bht_q[202:201], bht_q[199:198], bht_q[196:195], bht_q[193:192], bht_q[190:189], bht_q[187:186], bht_q[184:183], bht_q[181:180], bht_q[178:177], bht_q[175:174], bht_q[172:171], bht_q[169:168], bht_q[166:165], bht_q[163:162], bht_q[160:159], bht_q[157:156], bht_q[154:153], bht_q[151:150], bht_q[148:147], bht_q[145:144], bht_q[142:141], bht_q[139:138], bht_q[136:135], bht_q[133:132], bht_q[130:129], bht_q[127:126], bht_q[124:123], bht_q[121:120], bht_q[118:117], bht_q[115:114], bht_q[112:111], bht_q[109:108], bht_q[106:105], bht_q[103:102], bht_q[100:99], bht_q[97:96], bht_q[94:93], bht_q[91:90], bht_q[88:87], bht_q[85:84], bht_q[82:81], bht_q[79:78], bht_q[76:75], bht_q[73:72], bht_q[70:69], bht_q[67:66], bht_q[64:63], bht_q[61:60], bht_q[58:57], bht_q[55:54], bht_q[52:51], bht_q[49:48], bht_q[46:45], bht_q[43:42], bht_q[40:39], bht_q[37:36], bht_q[34:33], bht_q[31:30], bht_q[28:27], bht_q[25:24], bht_q[22:21], bht_q[19:18], bht_q[16:15], bht_q[13:12], bht_q[10:9], bht_q[7:6], bht_q[4:3], bht_q[1:0] } : 1'b0;
  assign N140 = N1060;
  assign N141 = bht_update_i[0];
  assign { N1580, N1579 } = (N12)? { N1578, N1577 } : 
                            (N928)? bht_q[1:0] : 1'b0;
  assign { N1582, N1581 } = (N13)? { N1578, N1577 } : 
                            (N929)? bht_q[4:3] : 1'b0;
  assign { N1584, N1583 } = (N14)? { N1578, N1577 } : 
                            (N930)? bht_q[7:6] : 1'b0;
  assign { N1586, N1585 } = (N15)? { N1578, N1577 } : 
                            (N931)? bht_q[10:9] : 1'b0;
  assign { N1588, N1587 } = (N16)? { N1578, N1577 } : 
                            (N932)? bht_q[13:12] : 1'b0;
  assign { N1590, N1589 } = (N17)? { N1578, N1577 } : 
                            (N933)? bht_q[16:15] : 1'b0;
  assign { N1592, N1591 } = (N18)? { N1578, N1577 } : 
                            (N934)? bht_q[19:18] : 1'b0;
  assign { N1594, N1593 } = (N19)? { N1578, N1577 } : 
                            (N935)? bht_q[22:21] : 1'b0;
  assign { N1596, N1595 } = (N20)? { N1578, N1577 } : 
                            (N936)? bht_q[25:24] : 1'b0;
  assign { N1598, N1597 } = (N21)? { N1578, N1577 } : 
                            (N937)? bht_q[28:27] : 1'b0;
  assign { N1600, N1599 } = (N22)? { N1578, N1577 } : 
                            (N938)? bht_q[31:30] : 1'b0;
  assign { N1602, N1601 } = (N23)? { N1578, N1577 } : 
                            (N939)? bht_q[34:33] : 1'b0;
  assign { N1604, N1603 } = (N24)? { N1578, N1577 } : 
                            (N940)? bht_q[37:36] : 1'b0;
  assign { N1606, N1605 } = (N25)? { N1578, N1577 } : 
                            (N941)? bht_q[40:39] : 1'b0;
  assign { N1608, N1607 } = (N26)? { N1578, N1577 } : 
                            (N942)? bht_q[43:42] : 1'b0;
  assign { N1610, N1609 } = (N27)? { N1578, N1577 } : 
                            (N943)? bht_q[46:45] : 1'b0;
  assign { N1612, N1611 } = (N28)? { N1578, N1577 } : 
                            (N944)? bht_q[49:48] : 1'b0;
  assign { N1614, N1613 } = (N29)? { N1578, N1577 } : 
                            (N945)? bht_q[52:51] : 1'b0;
  assign { N1616, N1615 } = (N30)? { N1578, N1577 } : 
                            (N946)? bht_q[55:54] : 1'b0;
  assign { N1618, N1617 } = (N31)? { N1578, N1577 } : 
                            (N947)? bht_q[58:57] : 1'b0;
  assign { N1620, N1619 } = (N32)? { N1578, N1577 } : 
                            (N948)? bht_q[61:60] : 1'b0;
  assign { N1622, N1621 } = (N33)? { N1578, N1577 } : 
                            (N949)? bht_q[64:63] : 1'b0;
  assign { N1624, N1623 } = (N34)? { N1578, N1577 } : 
                            (N950)? bht_q[67:66] : 1'b0;
  assign { N1626, N1625 } = (N35)? { N1578, N1577 } : 
                            (N951)? bht_q[70:69] : 1'b0;
  assign { N1628, N1627 } = (N36)? { N1578, N1577 } : 
                            (N952)? bht_q[73:72] : 1'b0;
  assign { N1630, N1629 } = (N37)? { N1578, N1577 } : 
                            (N953)? bht_q[76:75] : 1'b0;
  assign { N1632, N1631 } = (N38)? { N1578, N1577 } : 
                            (N954)? bht_q[79:78] : 1'b0;
  assign { N1634, N1633 } = (N39)? { N1578, N1577 } : 
                            (N955)? bht_q[82:81] : 1'b0;
  assign { N1636, N1635 } = (N40)? { N1578, N1577 } : 
                            (N956)? bht_q[85:84] : 1'b0;
  assign { N1638, N1637 } = (N41)? { N1578, N1577 } : 
                            (N957)? bht_q[88:87] : 1'b0;
  assign { N1640, N1639 } = (N42)? { N1578, N1577 } : 
                            (N958)? bht_q[91:90] : 1'b0;
  assign { N1642, N1641 } = (N43)? { N1578, N1577 } : 
                            (N959)? bht_q[94:93] : 1'b0;
  assign { N1644, N1643 } = (N44)? { N1578, N1577 } : 
                            (N960)? bht_q[97:96] : 1'b0;
  assign { N1646, N1645 } = (N45)? { N1578, N1577 } : 
                            (N961)? bht_q[100:99] : 1'b0;
  assign { N1648, N1647 } = (N46)? { N1578, N1577 } : 
                            (N962)? bht_q[103:102] : 1'b0;
  assign { N1650, N1649 } = (N47)? { N1578, N1577 } : 
                            (N963)? bht_q[106:105] : 1'b0;
  assign { N1652, N1651 } = (N48)? { N1578, N1577 } : 
                            (N964)? bht_q[109:108] : 1'b0;
  assign { N1654, N1653 } = (N49)? { N1578, N1577 } : 
                            (N965)? bht_q[112:111] : 1'b0;
  assign { N1656, N1655 } = (N50)? { N1578, N1577 } : 
                            (N966)? bht_q[115:114] : 1'b0;
  assign { N1658, N1657 } = (N51)? { N1578, N1577 } : 
                            (N967)? bht_q[118:117] : 1'b0;
  assign { N1660, N1659 } = (N52)? { N1578, N1577 } : 
                            (N968)? bht_q[121:120] : 1'b0;
  assign { N1662, N1661 } = (N53)? { N1578, N1577 } : 
                            (N969)? bht_q[124:123] : 1'b0;
  assign { N1664, N1663 } = (N54)? { N1578, N1577 } : 
                            (N970)? bht_q[127:126] : 1'b0;
  assign { N1666, N1665 } = (N55)? { N1578, N1577 } : 
                            (N971)? bht_q[130:129] : 1'b0;
  assign { N1668, N1667 } = (N56)? { N1578, N1577 } : 
                            (N972)? bht_q[133:132] : 1'b0;
  assign { N1670, N1669 } = (N57)? { N1578, N1577 } : 
                            (N973)? bht_q[136:135] : 1'b0;
  assign { N1672, N1671 } = (N58)? { N1578, N1577 } : 
                            (N974)? bht_q[139:138] : 1'b0;
  assign { N1674, N1673 } = (N59)? { N1578, N1577 } : 
                            (N975)? bht_q[142:141] : 1'b0;
  assign { N1676, N1675 } = (N60)? { N1578, N1577 } : 
                            (N976)? bht_q[145:144] : 1'b0;
  assign { N1678, N1677 } = (N61)? { N1578, N1577 } : 
                            (N977)? bht_q[148:147] : 1'b0;
  assign { N1680, N1679 } = (N62)? { N1578, N1577 } : 
                            (N978)? bht_q[151:150] : 1'b0;
  assign { N1682, N1681 } = (N63)? { N1578, N1577 } : 
                            (N979)? bht_q[154:153] : 1'b0;
  assign { N1684, N1683 } = (N64)? { N1578, N1577 } : 
                            (N980)? bht_q[157:156] : 1'b0;
  assign { N1686, N1685 } = (N65)? { N1578, N1577 } : 
                            (N981)? bht_q[160:159] : 1'b0;
  assign { N1688, N1687 } = (N66)? { N1578, N1577 } : 
                            (N982)? bht_q[163:162] : 1'b0;
  assign { N1690, N1689 } = (N67)? { N1578, N1577 } : 
                            (N983)? bht_q[166:165] : 1'b0;
  assign { N1692, N1691 } = (N68)? { N1578, N1577 } : 
                            (N984)? bht_q[169:168] : 1'b0;
  assign { N1694, N1693 } = (N69)? { N1578, N1577 } : 
                            (N985)? bht_q[172:171] : 1'b0;
  assign { N1696, N1695 } = (N70)? { N1578, N1577 } : 
                            (N986)? bht_q[175:174] : 1'b0;
  assign { N1698, N1697 } = (N71)? { N1578, N1577 } : 
                            (N987)? bht_q[178:177] : 1'b0;
  assign { N1700, N1699 } = (N72)? { N1578, N1577 } : 
                            (N988)? bht_q[181:180] : 1'b0;
  assign { N1702, N1701 } = (N73)? { N1578, N1577 } : 
                            (N989)? bht_q[184:183] : 1'b0;
  assign { N1704, N1703 } = (N74)? { N1578, N1577 } : 
                            (N990)? bht_q[187:186] : 1'b0;
  assign { N1706, N1705 } = (N75)? { N1578, N1577 } : 
                            (N991)? bht_q[190:189] : 1'b0;
  assign { N1708, N1707 } = (N76)? { N1578, N1577 } : 
                            (N992)? bht_q[193:192] : 1'b0;
  assign { N1710, N1709 } = (N77)? { N1578, N1577 } : 
                            (N993)? bht_q[196:195] : 1'b0;
  assign { N1712, N1711 } = (N78)? { N1578, N1577 } : 
                            (N994)? bht_q[199:198] : 1'b0;
  assign { N1714, N1713 } = (N79)? { N1578, N1577 } : 
                            (N995)? bht_q[202:201] : 1'b0;
  assign { N1716, N1715 } = (N80)? { N1578, N1577 } : 
                            (N996)? bht_q[205:204] : 1'b0;
  assign { N1718, N1717 } = (N81)? { N1578, N1577 } : 
                            (N997)? bht_q[208:207] : 1'b0;
  assign { N1720, N1719 } = (N82)? { N1578, N1577 } : 
                            (N998)? bht_q[211:210] : 1'b0;
  assign { N1722, N1721 } = (N83)? { N1578, N1577 } : 
                            (N999)? bht_q[214:213] : 1'b0;
  assign { N1724, N1723 } = (N84)? { N1578, N1577 } : 
                            (N1000)? bht_q[217:216] : 1'b0;
  assign { N1726, N1725 } = (N85)? { N1578, N1577 } : 
                            (N1001)? bht_q[220:219] : 1'b0;
  assign { N1728, N1727 } = (N86)? { N1578, N1577 } : 
                            (N1002)? bht_q[223:222] : 1'b0;
  assign { N1730, N1729 } = (N87)? { N1578, N1577 } : 
                            (N1003)? bht_q[226:225] : 1'b0;
  assign { N1732, N1731 } = (N88)? { N1578, N1577 } : 
                            (N1004)? bht_q[229:228] : 1'b0;
  assign { N1734, N1733 } = (N89)? { N1578, N1577 } : 
                            (N1005)? bht_q[232:231] : 1'b0;
  assign { N1736, N1735 } = (N90)? { N1578, N1577 } : 
                            (N1006)? bht_q[235:234] : 1'b0;
  assign { N1738, N1737 } = (N91)? { N1578, N1577 } : 
                            (N1007)? bht_q[238:237] : 1'b0;
  assign { N1740, N1739 } = (N92)? { N1578, N1577 } : 
                            (N1008)? bht_q[241:240] : 1'b0;
  assign { N1742, N1741 } = (N93)? { N1578, N1577 } : 
                            (N1009)? bht_q[244:243] : 1'b0;
  assign { N1744, N1743 } = (N94)? { N1578, N1577 } : 
                            (N1010)? bht_q[247:246] : 1'b0;
  assign { N1746, N1745 } = (N95)? { N1578, N1577 } : 
                            (N1011)? bht_q[250:249] : 1'b0;
  assign { N1748, N1747 } = (N96)? { N1578, N1577 } : 
                            (N1012)? bht_q[253:252] : 1'b0;
  assign { N1750, N1749 } = (N97)? { N1578, N1577 } : 
                            (N1013)? bht_q[256:255] : 1'b0;
  assign { N1752, N1751 } = (N98)? { N1578, N1577 } : 
                            (N1014)? bht_q[259:258] : 1'b0;
  assign { N1754, N1753 } = (N99)? { N1578, N1577 } : 
                            (N1015)? bht_q[262:261] : 1'b0;
  assign { N1756, N1755 } = (N100)? { N1578, N1577 } : 
                            (N1016)? bht_q[265:264] : 1'b0;
  assign { N1758, N1757 } = (N101)? { N1578, N1577 } : 
                            (N1017)? bht_q[268:267] : 1'b0;
  assign { N1760, N1759 } = (N102)? { N1578, N1577 } : 
                            (N1018)? bht_q[271:270] : 1'b0;
  assign { N1762, N1761 } = (N103)? { N1578, N1577 } : 
                            (N1019)? bht_q[274:273] : 1'b0;
  assign { N1764, N1763 } = (N104)? { N1578, N1577 } : 
                            (N1020)? bht_q[277:276] : 1'b0;
  assign { N1766, N1765 } = (N105)? { N1578, N1577 } : 
                            (N1021)? bht_q[280:279] : 1'b0;
  assign { N1768, N1767 } = (N106)? { N1578, N1577 } : 
                            (N1022)? bht_q[283:282] : 1'b0;
  assign { N1770, N1769 } = (N107)? { N1578, N1577 } : 
                            (N1023)? bht_q[286:285] : 1'b0;
  assign { N1772, N1771 } = (N108)? { N1578, N1577 } : 
                            (N1024)? bht_q[289:288] : 1'b0;
  assign { N1774, N1773 } = (N109)? { N1578, N1577 } : 
                            (N1025)? bht_q[292:291] : 1'b0;
  assign { N1776, N1775 } = (N110)? { N1578, N1577 } : 
                            (N1026)? bht_q[295:294] : 1'b0;
  assign { N1778, N1777 } = (N111)? { N1578, N1577 } : 
                            (N1027)? bht_q[298:297] : 1'b0;
  assign { N1780, N1779 } = (N112)? { N1578, N1577 } : 
                            (N1028)? bht_q[301:300] : 1'b0;
  assign { N1782, N1781 } = (N113)? { N1578, N1577 } : 
                            (N1029)? bht_q[304:303] : 1'b0;
  assign { N1784, N1783 } = (N114)? { N1578, N1577 } : 
                            (N1030)? bht_q[307:306] : 1'b0;
  assign { N1786, N1785 } = (N115)? { N1578, N1577 } : 
                            (N1031)? bht_q[310:309] : 1'b0;
  assign { N1788, N1787 } = (N116)? { N1578, N1577 } : 
                            (N1032)? bht_q[313:312] : 1'b0;
  assign { N1790, N1789 } = (N117)? { N1578, N1577 } : 
                            (N1033)? bht_q[316:315] : 1'b0;
  assign { N1792, N1791 } = (N118)? { N1578, N1577 } : 
                            (N1034)? bht_q[319:318] : 1'b0;
  assign { N1794, N1793 } = (N119)? { N1578, N1577 } : 
                            (N1035)? bht_q[322:321] : 1'b0;
  assign { N1796, N1795 } = (N120)? { N1578, N1577 } : 
                            (N1036)? bht_q[325:324] : 1'b0;
  assign { N1798, N1797 } = (N121)? { N1578, N1577 } : 
                            (N1037)? bht_q[328:327] : 1'b0;
  assign { N1800, N1799 } = (N122)? { N1578, N1577 } : 
                            (N1038)? bht_q[331:330] : 1'b0;
  assign { N1802, N1801 } = (N123)? { N1578, N1577 } : 
                            (N1039)? bht_q[334:333] : 1'b0;
  assign { N1804, N1803 } = (N124)? { N1578, N1577 } : 
                            (N1040)? bht_q[337:336] : 1'b0;
  assign { N1806, N1805 } = (N125)? { N1578, N1577 } : 
                            (N1041)? bht_q[340:339] : 1'b0;
  assign { N1808, N1807 } = (N126)? { N1578, N1577 } : 
                            (N1042)? bht_q[343:342] : 1'b0;
  assign { N1810, N1809 } = (N127)? { N1578, N1577 } : 
                            (N1043)? bht_q[346:345] : 1'b0;
  assign { N1812, N1811 } = (N128)? { N1578, N1577 } : 
                            (N1044)? bht_q[349:348] : 1'b0;
  assign { N1814, N1813 } = (N129)? { N1578, N1577 } : 
                            (N1045)? bht_q[352:351] : 1'b0;
  assign { N1816, N1815 } = (N130)? { N1578, N1577 } : 
                            (N1046)? bht_q[355:354] : 1'b0;
  assign { N1818, N1817 } = (N131)? { N1578, N1577 } : 
                            (N1047)? bht_q[358:357] : 1'b0;
  assign { N1820, N1819 } = (N132)? { N1578, N1577 } : 
                            (N1048)? bht_q[361:360] : 1'b0;
  assign { N1822, N1821 } = (N133)? { N1578, N1577 } : 
                            (N1049)? bht_q[364:363] : 1'b0;
  assign { N1824, N1823 } = (N134)? { N1578, N1577 } : 
                            (N1050)? bht_q[367:366] : 1'b0;
  assign { N1826, N1825 } = (N135)? { N1578, N1577 } : 
                            (N1051)? bht_q[370:369] : 1'b0;
  assign { N1828, N1827 } = (N136)? { N1578, N1577 } : 
                            (N1052)? bht_q[373:372] : 1'b0;
  assign { N1830, N1829 } = (N137)? { N1578, N1577 } : 
                            (N1053)? bht_q[376:375] : 1'b0;
  assign { N1832, N1831 } = (N138)? { N1578, N1577 } : 
                            (N1054)? bht_q[379:378] : 1'b0;
  assign { N1834, N1833 } = (N139)? { N1578, N1577 } : 
                            (N1055)? bht_q[382:381] : 1'b0;
  assign { N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835 } = (N141)? { N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1576)? { bht_q[382:381], bht_q[379:378], bht_q[376:375], bht_q[373:372], bht_q[370:369], bht_q[367:366], bht_q[364:363], bht_q[361:360], bht_q[358:357], bht_q[355:354], bht_q[352:351], bht_q[349:348], bht_q[346:345], bht_q[343:342], bht_q[340:339], bht_q[337:336], bht_q[334:333], bht_q[331:330], bht_q[328:327], bht_q[325:324], bht_q[322:321], bht_q[319:318], bht_q[316:315], bht_q[313:312], bht_q[310:309], bht_q[307:306], bht_q[304:303], bht_q[301:300], bht_q[298:297], bht_q[295:294], bht_q[292:291], bht_q[289:288], bht_q[286:285], bht_q[283:282], bht_q[280:279], bht_q[277:276], bht_q[274:273], bht_q[271:270], bht_q[268:267], bht_q[265:264], bht_q[262:261], bht_q[259:258], bht_q[256:255], bht_q[253:252], bht_q[250:249], bht_q[247:246], bht_q[244:243], bht_q[241:240], bht_q[238:237], bht_q[235:234], bht_q[232:231], bht_q[229:228], bht_q[226:225], bht_q[223:222], bht_q[220:219], bht_q[217:216], bht_q[214:213], bht_q[211:210], bht_q[208:207], bht_q[205:204], bht_q[202:201], bht_q[199:198], bht_q[196:195], bht_q[193:192], bht_q[190:189], bht_q[187:186], bht_q[184:183], bht_q[181:180], bht_q[178:177], bht_q[175:174], bht_q[172:171], bht_q[169:168], bht_q[166:165], bht_q[163:162], bht_q[160:159], bht_q[157:156], bht_q[154:153], bht_q[151:150], bht_q[148:147], bht_q[145:144], bht_q[142:141], bht_q[139:138], bht_q[136:135], bht_q[133:132], bht_q[130:129], bht_q[127:126], bht_q[124:123], bht_q[121:120], bht_q[118:117], bht_q[115:114], bht_q[112:111], bht_q[109:108], bht_q[106:105], bht_q[103:102], bht_q[100:99], bht_q[97:96], bht_q[94:93], bht_q[91:90], bht_q[88:87], bht_q[85:84], bht_q[82:81], bht_q[79:78], bht_q[76:75], bht_q[73:72], bht_q[70:69], bht_q[67:66], bht_q[64:63], bht_q[61:60], bht_q[58:57], bht_q[55:54], bht_q[52:51], bht_q[49:48], bht_q[46:45], bht_q[43:42], bht_q[40:39], bht_q[37:36], bht_q[34:33], bht_q[31:30], bht_q[28:27], bht_q[25:24], bht_q[22:21], bht_q[19:18], bht_q[16:15], bht_q[13:12], bht_q[10:9], bht_q[7:6], bht_q[4:3], bht_q[1:0] } : 1'b0;
  assign { N2095, N2094 } = (N12)? { N2093, N2092 } : 
                            (N928)? bht_q[1:0] : 1'b0;
  assign { N2097, N2096 } = (N13)? { N2093, N2092 } : 
                            (N929)? bht_q[4:3] : 1'b0;
  assign { N2099, N2098 } = (N14)? { N2093, N2092 } : 
                            (N930)? bht_q[7:6] : 1'b0;
  assign { N2101, N2100 } = (N15)? { N2093, N2092 } : 
                            (N931)? bht_q[10:9] : 1'b0;
  assign { N2103, N2102 } = (N16)? { N2093, N2092 } : 
                            (N932)? bht_q[13:12] : 1'b0;
  assign { N2105, N2104 } = (N17)? { N2093, N2092 } : 
                            (N933)? bht_q[16:15] : 1'b0;
  assign { N2107, N2106 } = (N18)? { N2093, N2092 } : 
                            (N934)? bht_q[19:18] : 1'b0;
  assign { N2109, N2108 } = (N19)? { N2093, N2092 } : 
                            (N935)? bht_q[22:21] : 1'b0;
  assign { N2111, N2110 } = (N20)? { N2093, N2092 } : 
                            (N936)? bht_q[25:24] : 1'b0;
  assign { N2113, N2112 } = (N21)? { N2093, N2092 } : 
                            (N937)? bht_q[28:27] : 1'b0;
  assign { N2115, N2114 } = (N22)? { N2093, N2092 } : 
                            (N938)? bht_q[31:30] : 1'b0;
  assign { N2117, N2116 } = (N23)? { N2093, N2092 } : 
                            (N939)? bht_q[34:33] : 1'b0;
  assign { N2119, N2118 } = (N24)? { N2093, N2092 } : 
                            (N940)? bht_q[37:36] : 1'b0;
  assign { N2121, N2120 } = (N25)? { N2093, N2092 } : 
                            (N941)? bht_q[40:39] : 1'b0;
  assign { N2123, N2122 } = (N26)? { N2093, N2092 } : 
                            (N942)? bht_q[43:42] : 1'b0;
  assign { N2125, N2124 } = (N27)? { N2093, N2092 } : 
                            (N943)? bht_q[46:45] : 1'b0;
  assign { N2127, N2126 } = (N28)? { N2093, N2092 } : 
                            (N944)? bht_q[49:48] : 1'b0;
  assign { N2129, N2128 } = (N29)? { N2093, N2092 } : 
                            (N945)? bht_q[52:51] : 1'b0;
  assign { N2131, N2130 } = (N30)? { N2093, N2092 } : 
                            (N946)? bht_q[55:54] : 1'b0;
  assign { N2133, N2132 } = (N31)? { N2093, N2092 } : 
                            (N947)? bht_q[58:57] : 1'b0;
  assign { N2135, N2134 } = (N32)? { N2093, N2092 } : 
                            (N948)? bht_q[61:60] : 1'b0;
  assign { N2137, N2136 } = (N33)? { N2093, N2092 } : 
                            (N949)? bht_q[64:63] : 1'b0;
  assign { N2139, N2138 } = (N34)? { N2093, N2092 } : 
                            (N950)? bht_q[67:66] : 1'b0;
  assign { N2141, N2140 } = (N35)? { N2093, N2092 } : 
                            (N951)? bht_q[70:69] : 1'b0;
  assign { N2143, N2142 } = (N36)? { N2093, N2092 } : 
                            (N952)? bht_q[73:72] : 1'b0;
  assign { N2145, N2144 } = (N37)? { N2093, N2092 } : 
                            (N953)? bht_q[76:75] : 1'b0;
  assign { N2147, N2146 } = (N38)? { N2093, N2092 } : 
                            (N954)? bht_q[79:78] : 1'b0;
  assign { N2149, N2148 } = (N39)? { N2093, N2092 } : 
                            (N955)? bht_q[82:81] : 1'b0;
  assign { N2151, N2150 } = (N40)? { N2093, N2092 } : 
                            (N956)? bht_q[85:84] : 1'b0;
  assign { N2153, N2152 } = (N41)? { N2093, N2092 } : 
                            (N957)? bht_q[88:87] : 1'b0;
  assign { N2155, N2154 } = (N42)? { N2093, N2092 } : 
                            (N958)? bht_q[91:90] : 1'b0;
  assign { N2157, N2156 } = (N43)? { N2093, N2092 } : 
                            (N959)? bht_q[94:93] : 1'b0;
  assign { N2159, N2158 } = (N44)? { N2093, N2092 } : 
                            (N960)? bht_q[97:96] : 1'b0;
  assign { N2161, N2160 } = (N45)? { N2093, N2092 } : 
                            (N961)? bht_q[100:99] : 1'b0;
  assign { N2163, N2162 } = (N46)? { N2093, N2092 } : 
                            (N962)? bht_q[103:102] : 1'b0;
  assign { N2165, N2164 } = (N47)? { N2093, N2092 } : 
                            (N963)? bht_q[106:105] : 1'b0;
  assign { N2167, N2166 } = (N48)? { N2093, N2092 } : 
                            (N964)? bht_q[109:108] : 1'b0;
  assign { N2169, N2168 } = (N49)? { N2093, N2092 } : 
                            (N965)? bht_q[112:111] : 1'b0;
  assign { N2171, N2170 } = (N50)? { N2093, N2092 } : 
                            (N966)? bht_q[115:114] : 1'b0;
  assign { N2173, N2172 } = (N51)? { N2093, N2092 } : 
                            (N967)? bht_q[118:117] : 1'b0;
  assign { N2175, N2174 } = (N52)? { N2093, N2092 } : 
                            (N968)? bht_q[121:120] : 1'b0;
  assign { N2177, N2176 } = (N53)? { N2093, N2092 } : 
                            (N969)? bht_q[124:123] : 1'b0;
  assign { N2179, N2178 } = (N54)? { N2093, N2092 } : 
                            (N970)? bht_q[127:126] : 1'b0;
  assign { N2181, N2180 } = (N55)? { N2093, N2092 } : 
                            (N971)? bht_q[130:129] : 1'b0;
  assign { N2183, N2182 } = (N56)? { N2093, N2092 } : 
                            (N972)? bht_q[133:132] : 1'b0;
  assign { N2185, N2184 } = (N57)? { N2093, N2092 } : 
                            (N973)? bht_q[136:135] : 1'b0;
  assign { N2187, N2186 } = (N58)? { N2093, N2092 } : 
                            (N974)? bht_q[139:138] : 1'b0;
  assign { N2189, N2188 } = (N59)? { N2093, N2092 } : 
                            (N975)? bht_q[142:141] : 1'b0;
  assign { N2191, N2190 } = (N60)? { N2093, N2092 } : 
                            (N976)? bht_q[145:144] : 1'b0;
  assign { N2193, N2192 } = (N61)? { N2093, N2092 } : 
                            (N977)? bht_q[148:147] : 1'b0;
  assign { N2195, N2194 } = (N62)? { N2093, N2092 } : 
                            (N978)? bht_q[151:150] : 1'b0;
  assign { N2197, N2196 } = (N63)? { N2093, N2092 } : 
                            (N979)? bht_q[154:153] : 1'b0;
  assign { N2199, N2198 } = (N64)? { N2093, N2092 } : 
                            (N980)? bht_q[157:156] : 1'b0;
  assign { N2201, N2200 } = (N65)? { N2093, N2092 } : 
                            (N981)? bht_q[160:159] : 1'b0;
  assign { N2203, N2202 } = (N66)? { N2093, N2092 } : 
                            (N982)? bht_q[163:162] : 1'b0;
  assign { N2205, N2204 } = (N67)? { N2093, N2092 } : 
                            (N983)? bht_q[166:165] : 1'b0;
  assign { N2207, N2206 } = (N68)? { N2093, N2092 } : 
                            (N984)? bht_q[169:168] : 1'b0;
  assign { N2209, N2208 } = (N69)? { N2093, N2092 } : 
                            (N985)? bht_q[172:171] : 1'b0;
  assign { N2211, N2210 } = (N70)? { N2093, N2092 } : 
                            (N986)? bht_q[175:174] : 1'b0;
  assign { N2213, N2212 } = (N71)? { N2093, N2092 } : 
                            (N987)? bht_q[178:177] : 1'b0;
  assign { N2215, N2214 } = (N72)? { N2093, N2092 } : 
                            (N988)? bht_q[181:180] : 1'b0;
  assign { N2217, N2216 } = (N73)? { N2093, N2092 } : 
                            (N989)? bht_q[184:183] : 1'b0;
  assign { N2219, N2218 } = (N74)? { N2093, N2092 } : 
                            (N990)? bht_q[187:186] : 1'b0;
  assign { N2221, N2220 } = (N75)? { N2093, N2092 } : 
                            (N991)? bht_q[190:189] : 1'b0;
  assign { N2223, N2222 } = (N76)? { N2093, N2092 } : 
                            (N992)? bht_q[193:192] : 1'b0;
  assign { N2225, N2224 } = (N77)? { N2093, N2092 } : 
                            (N993)? bht_q[196:195] : 1'b0;
  assign { N2227, N2226 } = (N78)? { N2093, N2092 } : 
                            (N994)? bht_q[199:198] : 1'b0;
  assign { N2229, N2228 } = (N79)? { N2093, N2092 } : 
                            (N995)? bht_q[202:201] : 1'b0;
  assign { N2231, N2230 } = (N80)? { N2093, N2092 } : 
                            (N996)? bht_q[205:204] : 1'b0;
  assign { N2233, N2232 } = (N81)? { N2093, N2092 } : 
                            (N997)? bht_q[208:207] : 1'b0;
  assign { N2235, N2234 } = (N82)? { N2093, N2092 } : 
                            (N998)? bht_q[211:210] : 1'b0;
  assign { N2237, N2236 } = (N83)? { N2093, N2092 } : 
                            (N999)? bht_q[214:213] : 1'b0;
  assign { N2239, N2238 } = (N84)? { N2093, N2092 } : 
                            (N1000)? bht_q[217:216] : 1'b0;
  assign { N2241, N2240 } = (N85)? { N2093, N2092 } : 
                            (N1001)? bht_q[220:219] : 1'b0;
  assign { N2243, N2242 } = (N86)? { N2093, N2092 } : 
                            (N1002)? bht_q[223:222] : 1'b0;
  assign { N2245, N2244 } = (N87)? { N2093, N2092 } : 
                            (N1003)? bht_q[226:225] : 1'b0;
  assign { N2247, N2246 } = (N88)? { N2093, N2092 } : 
                            (N1004)? bht_q[229:228] : 1'b0;
  assign { N2249, N2248 } = (N89)? { N2093, N2092 } : 
                            (N1005)? bht_q[232:231] : 1'b0;
  assign { N2251, N2250 } = (N90)? { N2093, N2092 } : 
                            (N1006)? bht_q[235:234] : 1'b0;
  assign { N2253, N2252 } = (N91)? { N2093, N2092 } : 
                            (N1007)? bht_q[238:237] : 1'b0;
  assign { N2255, N2254 } = (N92)? { N2093, N2092 } : 
                            (N1008)? bht_q[241:240] : 1'b0;
  assign { N2257, N2256 } = (N93)? { N2093, N2092 } : 
                            (N1009)? bht_q[244:243] : 1'b0;
  assign { N2259, N2258 } = (N94)? { N2093, N2092 } : 
                            (N1010)? bht_q[247:246] : 1'b0;
  assign { N2261, N2260 } = (N95)? { N2093, N2092 } : 
                            (N1011)? bht_q[250:249] : 1'b0;
  assign { N2263, N2262 } = (N96)? { N2093, N2092 } : 
                            (N1012)? bht_q[253:252] : 1'b0;
  assign { N2265, N2264 } = (N97)? { N2093, N2092 } : 
                            (N1013)? bht_q[256:255] : 1'b0;
  assign { N2267, N2266 } = (N98)? { N2093, N2092 } : 
                            (N1014)? bht_q[259:258] : 1'b0;
  assign { N2269, N2268 } = (N99)? { N2093, N2092 } : 
                            (N1015)? bht_q[262:261] : 1'b0;
  assign { N2271, N2270 } = (N100)? { N2093, N2092 } : 
                            (N1016)? bht_q[265:264] : 1'b0;
  assign { N2273, N2272 } = (N101)? { N2093, N2092 } : 
                            (N1017)? bht_q[268:267] : 1'b0;
  assign { N2275, N2274 } = (N102)? { N2093, N2092 } : 
                            (N1018)? bht_q[271:270] : 1'b0;
  assign { N2277, N2276 } = (N103)? { N2093, N2092 } : 
                            (N1019)? bht_q[274:273] : 1'b0;
  assign { N2279, N2278 } = (N104)? { N2093, N2092 } : 
                            (N1020)? bht_q[277:276] : 1'b0;
  assign { N2281, N2280 } = (N105)? { N2093, N2092 } : 
                            (N1021)? bht_q[280:279] : 1'b0;
  assign { N2283, N2282 } = (N106)? { N2093, N2092 } : 
                            (N1022)? bht_q[283:282] : 1'b0;
  assign { N2285, N2284 } = (N107)? { N2093, N2092 } : 
                            (N1023)? bht_q[286:285] : 1'b0;
  assign { N2287, N2286 } = (N108)? { N2093, N2092 } : 
                            (N1024)? bht_q[289:288] : 1'b0;
  assign { N2289, N2288 } = (N109)? { N2093, N2092 } : 
                            (N1025)? bht_q[292:291] : 1'b0;
  assign { N2291, N2290 } = (N110)? { N2093, N2092 } : 
                            (N1026)? bht_q[295:294] : 1'b0;
  assign { N2293, N2292 } = (N111)? { N2093, N2092 } : 
                            (N1027)? bht_q[298:297] : 1'b0;
  assign { N2295, N2294 } = (N112)? { N2093, N2092 } : 
                            (N1028)? bht_q[301:300] : 1'b0;
  assign { N2297, N2296 } = (N113)? { N2093, N2092 } : 
                            (N1029)? bht_q[304:303] : 1'b0;
  assign { N2299, N2298 } = (N114)? { N2093, N2092 } : 
                            (N1030)? bht_q[307:306] : 1'b0;
  assign { N2301, N2300 } = (N115)? { N2093, N2092 } : 
                            (N1031)? bht_q[310:309] : 1'b0;
  assign { N2303, N2302 } = (N116)? { N2093, N2092 } : 
                            (N1032)? bht_q[313:312] : 1'b0;
  assign { N2305, N2304 } = (N117)? { N2093, N2092 } : 
                            (N1033)? bht_q[316:315] : 1'b0;
  assign { N2307, N2306 } = (N118)? { N2093, N2092 } : 
                            (N1034)? bht_q[319:318] : 1'b0;
  assign { N2309, N2308 } = (N119)? { N2093, N2092 } : 
                            (N1035)? bht_q[322:321] : 1'b0;
  assign { N2311, N2310 } = (N120)? { N2093, N2092 } : 
                            (N1036)? bht_q[325:324] : 1'b0;
  assign { N2313, N2312 } = (N121)? { N2093, N2092 } : 
                            (N1037)? bht_q[328:327] : 1'b0;
  assign { N2315, N2314 } = (N122)? { N2093, N2092 } : 
                            (N1038)? bht_q[331:330] : 1'b0;
  assign { N2317, N2316 } = (N123)? { N2093, N2092 } : 
                            (N1039)? bht_q[334:333] : 1'b0;
  assign { N2319, N2318 } = (N124)? { N2093, N2092 } : 
                            (N1040)? bht_q[337:336] : 1'b0;
  assign { N2321, N2320 } = (N125)? { N2093, N2092 } : 
                            (N1041)? bht_q[340:339] : 1'b0;
  assign { N2323, N2322 } = (N126)? { N2093, N2092 } : 
                            (N1042)? bht_q[343:342] : 1'b0;
  assign { N2325, N2324 } = (N127)? { N2093, N2092 } : 
                            (N1043)? bht_q[346:345] : 1'b0;
  assign { N2327, N2326 } = (N128)? { N2093, N2092 } : 
                            (N1044)? bht_q[349:348] : 1'b0;
  assign { N2329, N2328 } = (N129)? { N2093, N2092 } : 
                            (N1045)? bht_q[352:351] : 1'b0;
  assign { N2331, N2330 } = (N130)? { N2093, N2092 } : 
                            (N1046)? bht_q[355:354] : 1'b0;
  assign { N2333, N2332 } = (N131)? { N2093, N2092 } : 
                            (N1047)? bht_q[358:357] : 1'b0;
  assign { N2335, N2334 } = (N132)? { N2093, N2092 } : 
                            (N1048)? bht_q[361:360] : 1'b0;
  assign { N2337, N2336 } = (N133)? { N2093, N2092 } : 
                            (N1049)? bht_q[364:363] : 1'b0;
  assign { N2339, N2338 } = (N134)? { N2093, N2092 } : 
                            (N1050)? bht_q[367:366] : 1'b0;
  assign { N2341, N2340 } = (N135)? { N2093, N2092 } : 
                            (N1051)? bht_q[370:369] : 1'b0;
  assign { N2343, N2342 } = (N136)? { N2093, N2092 } : 
                            (N1052)? bht_q[373:372] : 1'b0;
  assign { N2345, N2344 } = (N137)? { N2093, N2092 } : 
                            (N1053)? bht_q[376:375] : 1'b0;
  assign { N2347, N2346 } = (N138)? { N2093, N2092 } : 
                            (N1054)? bht_q[379:378] : 1'b0;
  assign { N2349, N2348 } = (N139)? { N2093, N2092 } : 
                            (N1055)? bht_q[382:381] : 1'b0;
  assign { N2353, N2352 } = (N12)? { N2351, N2350 } : 
                            (N928)? bht_q[1:0] : 1'b0;
  assign { N2355, N2354 } = (N13)? { N2351, N2350 } : 
                            (N929)? bht_q[4:3] : 1'b0;
  assign { N2357, N2356 } = (N14)? { N2351, N2350 } : 
                            (N930)? bht_q[7:6] : 1'b0;
  assign { N2359, N2358 } = (N15)? { N2351, N2350 } : 
                            (N931)? bht_q[10:9] : 1'b0;
  assign { N2361, N2360 } = (N16)? { N2351, N2350 } : 
                            (N932)? bht_q[13:12] : 1'b0;
  assign { N2363, N2362 } = (N17)? { N2351, N2350 } : 
                            (N933)? bht_q[16:15] : 1'b0;
  assign { N2365, N2364 } = (N18)? { N2351, N2350 } : 
                            (N934)? bht_q[19:18] : 1'b0;
  assign { N2367, N2366 } = (N19)? { N2351, N2350 } : 
                            (N935)? bht_q[22:21] : 1'b0;
  assign { N2369, N2368 } = (N20)? { N2351, N2350 } : 
                            (N936)? bht_q[25:24] : 1'b0;
  assign { N2371, N2370 } = (N21)? { N2351, N2350 } : 
                            (N937)? bht_q[28:27] : 1'b0;
  assign { N2373, N2372 } = (N22)? { N2351, N2350 } : 
                            (N938)? bht_q[31:30] : 1'b0;
  assign { N2375, N2374 } = (N23)? { N2351, N2350 } : 
                            (N939)? bht_q[34:33] : 1'b0;
  assign { N2377, N2376 } = (N24)? { N2351, N2350 } : 
                            (N940)? bht_q[37:36] : 1'b0;
  assign { N2379, N2378 } = (N25)? { N2351, N2350 } : 
                            (N941)? bht_q[40:39] : 1'b0;
  assign { N2381, N2380 } = (N26)? { N2351, N2350 } : 
                            (N942)? bht_q[43:42] : 1'b0;
  assign { N2383, N2382 } = (N27)? { N2351, N2350 } : 
                            (N943)? bht_q[46:45] : 1'b0;
  assign { N2385, N2384 } = (N28)? { N2351, N2350 } : 
                            (N944)? bht_q[49:48] : 1'b0;
  assign { N2387, N2386 } = (N29)? { N2351, N2350 } : 
                            (N945)? bht_q[52:51] : 1'b0;
  assign { N2389, N2388 } = (N30)? { N2351, N2350 } : 
                            (N946)? bht_q[55:54] : 1'b0;
  assign { N2391, N2390 } = (N31)? { N2351, N2350 } : 
                            (N947)? bht_q[58:57] : 1'b0;
  assign { N2393, N2392 } = (N32)? { N2351, N2350 } : 
                            (N948)? bht_q[61:60] : 1'b0;
  assign { N2395, N2394 } = (N33)? { N2351, N2350 } : 
                            (N949)? bht_q[64:63] : 1'b0;
  assign { N2397, N2396 } = (N34)? { N2351, N2350 } : 
                            (N950)? bht_q[67:66] : 1'b0;
  assign { N2399, N2398 } = (N35)? { N2351, N2350 } : 
                            (N951)? bht_q[70:69] : 1'b0;
  assign { N2401, N2400 } = (N36)? { N2351, N2350 } : 
                            (N952)? bht_q[73:72] : 1'b0;
  assign { N2403, N2402 } = (N37)? { N2351, N2350 } : 
                            (N953)? bht_q[76:75] : 1'b0;
  assign { N2405, N2404 } = (N38)? { N2351, N2350 } : 
                            (N954)? bht_q[79:78] : 1'b0;
  assign { N2407, N2406 } = (N39)? { N2351, N2350 } : 
                            (N955)? bht_q[82:81] : 1'b0;
  assign { N2409, N2408 } = (N40)? { N2351, N2350 } : 
                            (N956)? bht_q[85:84] : 1'b0;
  assign { N2411, N2410 } = (N41)? { N2351, N2350 } : 
                            (N957)? bht_q[88:87] : 1'b0;
  assign { N2413, N2412 } = (N42)? { N2351, N2350 } : 
                            (N958)? bht_q[91:90] : 1'b0;
  assign { N2415, N2414 } = (N43)? { N2351, N2350 } : 
                            (N959)? bht_q[94:93] : 1'b0;
  assign { N2417, N2416 } = (N44)? { N2351, N2350 } : 
                            (N960)? bht_q[97:96] : 1'b0;
  assign { N2419, N2418 } = (N45)? { N2351, N2350 } : 
                            (N961)? bht_q[100:99] : 1'b0;
  assign { N2421, N2420 } = (N46)? { N2351, N2350 } : 
                            (N962)? bht_q[103:102] : 1'b0;
  assign { N2423, N2422 } = (N47)? { N2351, N2350 } : 
                            (N963)? bht_q[106:105] : 1'b0;
  assign { N2425, N2424 } = (N48)? { N2351, N2350 } : 
                            (N964)? bht_q[109:108] : 1'b0;
  assign { N2427, N2426 } = (N49)? { N2351, N2350 } : 
                            (N965)? bht_q[112:111] : 1'b0;
  assign { N2429, N2428 } = (N50)? { N2351, N2350 } : 
                            (N966)? bht_q[115:114] : 1'b0;
  assign { N2431, N2430 } = (N51)? { N2351, N2350 } : 
                            (N967)? bht_q[118:117] : 1'b0;
  assign { N2433, N2432 } = (N52)? { N2351, N2350 } : 
                            (N968)? bht_q[121:120] : 1'b0;
  assign { N2435, N2434 } = (N53)? { N2351, N2350 } : 
                            (N969)? bht_q[124:123] : 1'b0;
  assign { N2437, N2436 } = (N54)? { N2351, N2350 } : 
                            (N970)? bht_q[127:126] : 1'b0;
  assign { N2439, N2438 } = (N55)? { N2351, N2350 } : 
                            (N971)? bht_q[130:129] : 1'b0;
  assign { N2441, N2440 } = (N56)? { N2351, N2350 } : 
                            (N972)? bht_q[133:132] : 1'b0;
  assign { N2443, N2442 } = (N57)? { N2351, N2350 } : 
                            (N973)? bht_q[136:135] : 1'b0;
  assign { N2445, N2444 } = (N58)? { N2351, N2350 } : 
                            (N974)? bht_q[139:138] : 1'b0;
  assign { N2447, N2446 } = (N59)? { N2351, N2350 } : 
                            (N975)? bht_q[142:141] : 1'b0;
  assign { N2449, N2448 } = (N60)? { N2351, N2350 } : 
                            (N976)? bht_q[145:144] : 1'b0;
  assign { N2451, N2450 } = (N61)? { N2351, N2350 } : 
                            (N977)? bht_q[148:147] : 1'b0;
  assign { N2453, N2452 } = (N62)? { N2351, N2350 } : 
                            (N978)? bht_q[151:150] : 1'b0;
  assign { N2455, N2454 } = (N63)? { N2351, N2350 } : 
                            (N979)? bht_q[154:153] : 1'b0;
  assign { N2457, N2456 } = (N64)? { N2351, N2350 } : 
                            (N980)? bht_q[157:156] : 1'b0;
  assign { N2459, N2458 } = (N65)? { N2351, N2350 } : 
                            (N981)? bht_q[160:159] : 1'b0;
  assign { N2461, N2460 } = (N66)? { N2351, N2350 } : 
                            (N982)? bht_q[163:162] : 1'b0;
  assign { N2463, N2462 } = (N67)? { N2351, N2350 } : 
                            (N983)? bht_q[166:165] : 1'b0;
  assign { N2465, N2464 } = (N68)? { N2351, N2350 } : 
                            (N984)? bht_q[169:168] : 1'b0;
  assign { N2467, N2466 } = (N69)? { N2351, N2350 } : 
                            (N985)? bht_q[172:171] : 1'b0;
  assign { N2469, N2468 } = (N70)? { N2351, N2350 } : 
                            (N986)? bht_q[175:174] : 1'b0;
  assign { N2471, N2470 } = (N71)? { N2351, N2350 } : 
                            (N987)? bht_q[178:177] : 1'b0;
  assign { N2473, N2472 } = (N72)? { N2351, N2350 } : 
                            (N988)? bht_q[181:180] : 1'b0;
  assign { N2475, N2474 } = (N73)? { N2351, N2350 } : 
                            (N989)? bht_q[184:183] : 1'b0;
  assign { N2477, N2476 } = (N74)? { N2351, N2350 } : 
                            (N990)? bht_q[187:186] : 1'b0;
  assign { N2479, N2478 } = (N75)? { N2351, N2350 } : 
                            (N991)? bht_q[190:189] : 1'b0;
  assign { N2481, N2480 } = (N76)? { N2351, N2350 } : 
                            (N992)? bht_q[193:192] : 1'b0;
  assign { N2483, N2482 } = (N77)? { N2351, N2350 } : 
                            (N993)? bht_q[196:195] : 1'b0;
  assign { N2485, N2484 } = (N78)? { N2351, N2350 } : 
                            (N994)? bht_q[199:198] : 1'b0;
  assign { N2487, N2486 } = (N79)? { N2351, N2350 } : 
                            (N995)? bht_q[202:201] : 1'b0;
  assign { N2489, N2488 } = (N80)? { N2351, N2350 } : 
                            (N996)? bht_q[205:204] : 1'b0;
  assign { N2491, N2490 } = (N81)? { N2351, N2350 } : 
                            (N997)? bht_q[208:207] : 1'b0;
  assign { N2493, N2492 } = (N82)? { N2351, N2350 } : 
                            (N998)? bht_q[211:210] : 1'b0;
  assign { N2495, N2494 } = (N83)? { N2351, N2350 } : 
                            (N999)? bht_q[214:213] : 1'b0;
  assign { N2497, N2496 } = (N84)? { N2351, N2350 } : 
                            (N1000)? bht_q[217:216] : 1'b0;
  assign { N2499, N2498 } = (N85)? { N2351, N2350 } : 
                            (N1001)? bht_q[220:219] : 1'b0;
  assign { N2501, N2500 } = (N86)? { N2351, N2350 } : 
                            (N1002)? bht_q[223:222] : 1'b0;
  assign { N2503, N2502 } = (N87)? { N2351, N2350 } : 
                            (N1003)? bht_q[226:225] : 1'b0;
  assign { N2505, N2504 } = (N88)? { N2351, N2350 } : 
                            (N1004)? bht_q[229:228] : 1'b0;
  assign { N2507, N2506 } = (N89)? { N2351, N2350 } : 
                            (N1005)? bht_q[232:231] : 1'b0;
  assign { N2509, N2508 } = (N90)? { N2351, N2350 } : 
                            (N1006)? bht_q[235:234] : 1'b0;
  assign { N2511, N2510 } = (N91)? { N2351, N2350 } : 
                            (N1007)? bht_q[238:237] : 1'b0;
  assign { N2513, N2512 } = (N92)? { N2351, N2350 } : 
                            (N1008)? bht_q[241:240] : 1'b0;
  assign { N2515, N2514 } = (N93)? { N2351, N2350 } : 
                            (N1009)? bht_q[244:243] : 1'b0;
  assign { N2517, N2516 } = (N94)? { N2351, N2350 } : 
                            (N1010)? bht_q[247:246] : 1'b0;
  assign { N2519, N2518 } = (N95)? { N2351, N2350 } : 
                            (N1011)? bht_q[250:249] : 1'b0;
  assign { N2521, N2520 } = (N96)? { N2351, N2350 } : 
                            (N1012)? bht_q[253:252] : 1'b0;
  assign { N2523, N2522 } = (N97)? { N2351, N2350 } : 
                            (N1013)? bht_q[256:255] : 1'b0;
  assign { N2525, N2524 } = (N98)? { N2351, N2350 } : 
                            (N1014)? bht_q[259:258] : 1'b0;
  assign { N2527, N2526 } = (N99)? { N2351, N2350 } : 
                            (N1015)? bht_q[262:261] : 1'b0;
  assign { N2529, N2528 } = (N100)? { N2351, N2350 } : 
                            (N1016)? bht_q[265:264] : 1'b0;
  assign { N2531, N2530 } = (N101)? { N2351, N2350 } : 
                            (N1017)? bht_q[268:267] : 1'b0;
  assign { N2533, N2532 } = (N102)? { N2351, N2350 } : 
                            (N1018)? bht_q[271:270] : 1'b0;
  assign { N2535, N2534 } = (N103)? { N2351, N2350 } : 
                            (N1019)? bht_q[274:273] : 1'b0;
  assign { N2537, N2536 } = (N104)? { N2351, N2350 } : 
                            (N1020)? bht_q[277:276] : 1'b0;
  assign { N2539, N2538 } = (N105)? { N2351, N2350 } : 
                            (N1021)? bht_q[280:279] : 1'b0;
  assign { N2541, N2540 } = (N106)? { N2351, N2350 } : 
                            (N1022)? bht_q[283:282] : 1'b0;
  assign { N2543, N2542 } = (N107)? { N2351, N2350 } : 
                            (N1023)? bht_q[286:285] : 1'b0;
  assign { N2545, N2544 } = (N108)? { N2351, N2350 } : 
                            (N1024)? bht_q[289:288] : 1'b0;
  assign { N2547, N2546 } = (N109)? { N2351, N2350 } : 
                            (N1025)? bht_q[292:291] : 1'b0;
  assign { N2549, N2548 } = (N110)? { N2351, N2350 } : 
                            (N1026)? bht_q[295:294] : 1'b0;
  assign { N2551, N2550 } = (N111)? { N2351, N2350 } : 
                            (N1027)? bht_q[298:297] : 1'b0;
  assign { N2553, N2552 } = (N112)? { N2351, N2350 } : 
                            (N1028)? bht_q[301:300] : 1'b0;
  assign { N2555, N2554 } = (N113)? { N2351, N2350 } : 
                            (N1029)? bht_q[304:303] : 1'b0;
  assign { N2557, N2556 } = (N114)? { N2351, N2350 } : 
                            (N1030)? bht_q[307:306] : 1'b0;
  assign { N2559, N2558 } = (N115)? { N2351, N2350 } : 
                            (N1031)? bht_q[310:309] : 1'b0;
  assign { N2561, N2560 } = (N116)? { N2351, N2350 } : 
                            (N1032)? bht_q[313:312] : 1'b0;
  assign { N2563, N2562 } = (N117)? { N2351, N2350 } : 
                            (N1033)? bht_q[316:315] : 1'b0;
  assign { N2565, N2564 } = (N118)? { N2351, N2350 } : 
                            (N1034)? bht_q[319:318] : 1'b0;
  assign { N2567, N2566 } = (N119)? { N2351, N2350 } : 
                            (N1035)? bht_q[322:321] : 1'b0;
  assign { N2569, N2568 } = (N120)? { N2351, N2350 } : 
                            (N1036)? bht_q[325:324] : 1'b0;
  assign { N2571, N2570 } = (N121)? { N2351, N2350 } : 
                            (N1037)? bht_q[328:327] : 1'b0;
  assign { N2573, N2572 } = (N122)? { N2351, N2350 } : 
                            (N1038)? bht_q[331:330] : 1'b0;
  assign { N2575, N2574 } = (N123)? { N2351, N2350 } : 
                            (N1039)? bht_q[334:333] : 1'b0;
  assign { N2577, N2576 } = (N124)? { N2351, N2350 } : 
                            (N1040)? bht_q[337:336] : 1'b0;
  assign { N2579, N2578 } = (N125)? { N2351, N2350 } : 
                            (N1041)? bht_q[340:339] : 1'b0;
  assign { N2581, N2580 } = (N126)? { N2351, N2350 } : 
                            (N1042)? bht_q[343:342] : 1'b0;
  assign { N2583, N2582 } = (N127)? { N2351, N2350 } : 
                            (N1043)? bht_q[346:345] : 1'b0;
  assign { N2585, N2584 } = (N128)? { N2351, N2350 } : 
                            (N1044)? bht_q[349:348] : 1'b0;
  assign { N2587, N2586 } = (N129)? { N2351, N2350 } : 
                            (N1045)? bht_q[352:351] : 1'b0;
  assign { N2589, N2588 } = (N130)? { N2351, N2350 } : 
                            (N1046)? bht_q[355:354] : 1'b0;
  assign { N2591, N2590 } = (N131)? { N2351, N2350 } : 
                            (N1047)? bht_q[358:357] : 1'b0;
  assign { N2593, N2592 } = (N132)? { N2351, N2350 } : 
                            (N1048)? bht_q[361:360] : 1'b0;
  assign { N2595, N2594 } = (N133)? { N2351, N2350 } : 
                            (N1049)? bht_q[364:363] : 1'b0;
  assign { N2597, N2596 } = (N134)? { N2351, N2350 } : 
                            (N1050)? bht_q[367:366] : 1'b0;
  assign { N2599, N2598 } = (N135)? { N2351, N2350 } : 
                            (N1051)? bht_q[370:369] : 1'b0;
  assign { N2601, N2600 } = (N136)? { N2351, N2350 } : 
                            (N1052)? bht_q[373:372] : 1'b0;
  assign { N2603, N2602 } = (N137)? { N2351, N2350 } : 
                            (N1053)? bht_q[376:375] : 1'b0;
  assign { N2605, N2604 } = (N138)? { N2351, N2350 } : 
                            (N1054)? bht_q[379:378] : 1'b0;
  assign { N2607, N2606 } = (N139)? { N2351, N2350 } : 
                            (N1055)? bht_q[382:381] : 1'b0;
  assign { N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608 } = (N142)? { N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2865)? { N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2867)? { N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1058)? { N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352 } : 1'b0;
  assign N142 = N3524;
  assign { N3125, N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870 } = (N143)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N144)? { N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608 } : 1'b0;
  assign N143 = flush_i;
  assign N144 = N2869;
  assign N145 = ~vpc_i[2];
  assign N146 = ~vpc_i[3];
  assign N147 = N145 & N146;
  assign N148 = N145 & vpc_i[3];
  assign N149 = vpc_i[2] & N146;
  assign N150 = vpc_i[2] & vpc_i[3];
  assign N151 = ~vpc_i[4];
  assign N152 = N147 & N151;
  assign N153 = N147 & vpc_i[4];
  assign N154 = N149 & N151;
  assign N155 = N149 & vpc_i[4];
  assign N156 = N148 & N151;
  assign N157 = N148 & vpc_i[4];
  assign N158 = N150 & N151;
  assign N159 = N150 & vpc_i[4];
  assign N160 = ~vpc_i[5];
  assign N161 = N152 & N160;
  assign N162 = N152 & vpc_i[5];
  assign N163 = N154 & N160;
  assign N164 = N154 & vpc_i[5];
  assign N165 = N156 & N160;
  assign N166 = N156 & vpc_i[5];
  assign N167 = N158 & N160;
  assign N168 = N158 & vpc_i[5];
  assign N169 = N153 & N160;
  assign N170 = N153 & vpc_i[5];
  assign N171 = N155 & N160;
  assign N172 = N155 & vpc_i[5];
  assign N173 = N157 & N160;
  assign N174 = N157 & vpc_i[5];
  assign N175 = N159 & N160;
  assign N176 = N159 & vpc_i[5];
  assign N177 = ~vpc_i[6];
  assign N178 = N161 & N177;
  assign N179 = N161 & vpc_i[6];
  assign N180 = N163 & N177;
  assign N181 = N163 & vpc_i[6];
  assign N182 = N165 & N177;
  assign N183 = N165 & vpc_i[6];
  assign N184 = N167 & N177;
  assign N185 = N167 & vpc_i[6];
  assign N186 = N169 & N177;
  assign N187 = N169 & vpc_i[6];
  assign N188 = N171 & N177;
  assign N189 = N171 & vpc_i[6];
  assign N190 = N173 & N177;
  assign N191 = N173 & vpc_i[6];
  assign N192 = N175 & N177;
  assign N193 = N175 & vpc_i[6];
  assign N194 = N162 & N177;
  assign N195 = N162 & vpc_i[6];
  assign N196 = N164 & N177;
  assign N197 = N164 & vpc_i[6];
  assign N198 = N166 & N177;
  assign N199 = N166 & vpc_i[6];
  assign N200 = N168 & N177;
  assign N201 = N168 & vpc_i[6];
  assign N202 = N170 & N177;
  assign N203 = N170 & vpc_i[6];
  assign N204 = N172 & N177;
  assign N205 = N172 & vpc_i[6];
  assign N206 = N174 & N177;
  assign N207 = N174 & vpc_i[6];
  assign N208 = N176 & N177;
  assign N209 = N176 & vpc_i[6];
  assign N210 = ~vpc_i[7];
  assign N211 = N178 & N210;
  assign N212 = N178 & vpc_i[7];
  assign N213 = N180 & N210;
  assign N214 = N180 & vpc_i[7];
  assign N215 = N182 & N210;
  assign N216 = N182 & vpc_i[7];
  assign N217 = N184 & N210;
  assign N218 = N184 & vpc_i[7];
  assign N219 = N186 & N210;
  assign N220 = N186 & vpc_i[7];
  assign N221 = N188 & N210;
  assign N222 = N188 & vpc_i[7];
  assign N223 = N190 & N210;
  assign N224 = N190 & vpc_i[7];
  assign N225 = N192 & N210;
  assign N226 = N192 & vpc_i[7];
  assign N227 = N194 & N210;
  assign N228 = N194 & vpc_i[7];
  assign N229 = N196 & N210;
  assign N230 = N196 & vpc_i[7];
  assign N231 = N198 & N210;
  assign N232 = N198 & vpc_i[7];
  assign N233 = N200 & N210;
  assign N234 = N200 & vpc_i[7];
  assign N235 = N202 & N210;
  assign N236 = N202 & vpc_i[7];
  assign N237 = N204 & N210;
  assign N238 = N204 & vpc_i[7];
  assign N239 = N206 & N210;
  assign N240 = N206 & vpc_i[7];
  assign N241 = N208 & N210;
  assign N242 = N208 & vpc_i[7];
  assign N243 = N179 & N210;
  assign N244 = N179 & vpc_i[7];
  assign N245 = N181 & N210;
  assign N246 = N181 & vpc_i[7];
  assign N247 = N183 & N210;
  assign N248 = N183 & vpc_i[7];
  assign N249 = N185 & N210;
  assign N250 = N185 & vpc_i[7];
  assign N251 = N187 & N210;
  assign N252 = N187 & vpc_i[7];
  assign N253 = N189 & N210;
  assign N254 = N189 & vpc_i[7];
  assign N255 = N191 & N210;
  assign N256 = N191 & vpc_i[7];
  assign N257 = N193 & N210;
  assign N258 = N193 & vpc_i[7];
  assign N259 = N195 & N210;
  assign N260 = N195 & vpc_i[7];
  assign N261 = N197 & N210;
  assign N262 = N197 & vpc_i[7];
  assign N263 = N199 & N210;
  assign N264 = N199 & vpc_i[7];
  assign N265 = N201 & N210;
  assign N266 = N201 & vpc_i[7];
  assign N267 = N203 & N210;
  assign N268 = N203 & vpc_i[7];
  assign N269 = N205 & N210;
  assign N270 = N205 & vpc_i[7];
  assign N271 = N207 & N210;
  assign N272 = N207 & vpc_i[7];
  assign N273 = N209 & N210;
  assign N274 = N209 & vpc_i[7];
  assign N275 = ~vpc_i[8];
  assign N276 = N211 & N275;
  assign N277 = N211 & vpc_i[8];
  assign N278 = N213 & N275;
  assign N279 = N213 & vpc_i[8];
  assign N280 = N215 & N275;
  assign N281 = N215 & vpc_i[8];
  assign N282 = N217 & N275;
  assign N283 = N217 & vpc_i[8];
  assign N284 = N219 & N275;
  assign N285 = N219 & vpc_i[8];
  assign N286 = N221 & N275;
  assign N287 = N221 & vpc_i[8];
  assign N288 = N223 & N275;
  assign N289 = N223 & vpc_i[8];
  assign N290 = N225 & N275;
  assign N291 = N225 & vpc_i[8];
  assign N292 = N227 & N275;
  assign N293 = N227 & vpc_i[8];
  assign N294 = N229 & N275;
  assign N295 = N229 & vpc_i[8];
  assign N296 = N231 & N275;
  assign N297 = N231 & vpc_i[8];
  assign N298 = N233 & N275;
  assign N299 = N233 & vpc_i[8];
  assign N300 = N235 & N275;
  assign N301 = N235 & vpc_i[8];
  assign N302 = N237 & N275;
  assign N303 = N237 & vpc_i[8];
  assign N304 = N239 & N275;
  assign N305 = N239 & vpc_i[8];
  assign N306 = N241 & N275;
  assign N307 = N241 & vpc_i[8];
  assign N308 = N243 & N275;
  assign N309 = N243 & vpc_i[8];
  assign N310 = N245 & N275;
  assign N311 = N245 & vpc_i[8];
  assign N312 = N247 & N275;
  assign N313 = N247 & vpc_i[8];
  assign N314 = N249 & N275;
  assign N315 = N249 & vpc_i[8];
  assign N316 = N251 & N275;
  assign N317 = N251 & vpc_i[8];
  assign N318 = N253 & N275;
  assign N319 = N253 & vpc_i[8];
  assign N320 = N255 & N275;
  assign N321 = N255 & vpc_i[8];
  assign N322 = N257 & N275;
  assign N323 = N257 & vpc_i[8];
  assign N324 = N259 & N275;
  assign N325 = N259 & vpc_i[8];
  assign N326 = N261 & N275;
  assign N327 = N261 & vpc_i[8];
  assign N328 = N263 & N275;
  assign N329 = N263 & vpc_i[8];
  assign N330 = N265 & N275;
  assign N331 = N265 & vpc_i[8];
  assign N332 = N267 & N275;
  assign N333 = N267 & vpc_i[8];
  assign N334 = N269 & N275;
  assign N335 = N269 & vpc_i[8];
  assign N336 = N271 & N275;
  assign N337 = N271 & vpc_i[8];
  assign N338 = N273 & N275;
  assign N339 = N273 & vpc_i[8];
  assign N340 = N212 & N275;
  assign N341 = N212 & vpc_i[8];
  assign N342 = N214 & N275;
  assign N343 = N214 & vpc_i[8];
  assign N344 = N216 & N275;
  assign N345 = N216 & vpc_i[8];
  assign N346 = N218 & N275;
  assign N347 = N218 & vpc_i[8];
  assign N348 = N220 & N275;
  assign N349 = N220 & vpc_i[8];
  assign N350 = N222 & N275;
  assign N351 = N222 & vpc_i[8];
  assign N352 = N224 & N275;
  assign N353 = N224 & vpc_i[8];
  assign N354 = N226 & N275;
  assign N355 = N226 & vpc_i[8];
  assign N356 = N228 & N275;
  assign N357 = N228 & vpc_i[8];
  assign N358 = N230 & N275;
  assign N359 = N230 & vpc_i[8];
  assign N360 = N232 & N275;
  assign N361 = N232 & vpc_i[8];
  assign N362 = N234 & N275;
  assign N363 = N234 & vpc_i[8];
  assign N364 = N236 & N275;
  assign N365 = N236 & vpc_i[8];
  assign N366 = N238 & N275;
  assign N367 = N238 & vpc_i[8];
  assign N368 = N240 & N275;
  assign N369 = N240 & vpc_i[8];
  assign N370 = N242 & N275;
  assign N371 = N242 & vpc_i[8];
  assign N372 = N244 & N275;
  assign N373 = N244 & vpc_i[8];
  assign N374 = N246 & N275;
  assign N375 = N246 & vpc_i[8];
  assign N376 = N248 & N275;
  assign N377 = N248 & vpc_i[8];
  assign N378 = N250 & N275;
  assign N379 = N250 & vpc_i[8];
  assign N380 = N252 & N275;
  assign N381 = N252 & vpc_i[8];
  assign N382 = N254 & N275;
  assign N383 = N254 & vpc_i[8];
  assign N384 = N256 & N275;
  assign N385 = N256 & vpc_i[8];
  assign N386 = N258 & N275;
  assign N387 = N258 & vpc_i[8];
  assign N388 = N260 & N275;
  assign N389 = N260 & vpc_i[8];
  assign N390 = N262 & N275;
  assign N391 = N262 & vpc_i[8];
  assign N392 = N264 & N275;
  assign N393 = N264 & vpc_i[8];
  assign N394 = N266 & N275;
  assign N395 = N266 & vpc_i[8];
  assign N396 = N268 & N275;
  assign N397 = N268 & vpc_i[8];
  assign N398 = N270 & N275;
  assign N399 = N270 & vpc_i[8];
  assign N400 = N272 & N275;
  assign N401 = N272 & vpc_i[8];
  assign N402 = N274 & N275;
  assign N403 = N274 & vpc_i[8];
  assign N404 = N211 & N275;
  assign N405 = N213 & N275;
  assign N406 = N215 & N275;
  assign N407 = N217 & N275;
  assign N408 = N219 & N275;
  assign N409 = N221 & N275;
  assign N410 = N223 & N275;
  assign N411 = N225 & N275;
  assign N412 = N227 & N275;
  assign N413 = N229 & N275;
  assign N414 = N231 & N275;
  assign N415 = N233 & N275;
  assign N416 = N235 & N275;
  assign N417 = N237 & N275;
  assign N418 = N239 & N275;
  assign N419 = N241 & N275;
  assign N420 = N243 & N275;
  assign N421 = N245 & N275;
  assign N422 = N247 & N275;
  assign N423 = N249 & N275;
  assign N424 = N251 & N275;
  assign N425 = N253 & N275;
  assign N426 = N255 & N275;
  assign N427 = N257 & N275;
  assign N428 = N259 & N275;
  assign N429 = N261 & N275;
  assign N430 = N263 & N275;
  assign N431 = N265 & N275;
  assign N432 = N267 & N275;
  assign N433 = N269 & N275;
  assign N434 = N271 & N275;
  assign N435 = N273 & N275;
  assign N436 = N212 & N275;
  assign N437 = N214 & N275;
  assign N438 = N216 & N275;
  assign N439 = N218 & N275;
  assign N440 = N220 & N275;
  assign N441 = N222 & N275;
  assign N442 = N224 & N275;
  assign N443 = N226 & N275;
  assign N444 = N228 & N275;
  assign N445 = N230 & N275;
  assign N446 = N232 & N275;
  assign N447 = N234 & N275;
  assign N448 = N236 & N275;
  assign N449 = N238 & N275;
  assign N450 = N240 & N275;
  assign N451 = N242 & N275;
  assign N452 = N244 & N275;
  assign N453 = N246 & N275;
  assign N454 = N248 & N275;
  assign N455 = N250 & N275;
  assign N456 = N252 & N275;
  assign N457 = N254 & N275;
  assign N458 = N256 & N275;
  assign N459 = N258 & N275;
  assign N460 = N260 & N275;
  assign N461 = N262 & N275;
  assign N462 = N264 & N275;
  assign N463 = N266 & N275;
  assign N464 = N268 & N275;
  assign N465 = N270 & N275;
  assign N466 = N272 & N275;
  assign N467 = N274 & N275;
  assign N470 = N211 & N275;
  assign N471 = N213 & N275;
  assign N472 = N215 & N275;
  assign N473 = N217 & N275;
  assign N474 = N219 & N275;
  assign N475 = N221 & N275;
  assign N476 = N223 & N275;
  assign N477 = N225 & N275;
  assign N478 = N227 & N275;
  assign N479 = N229 & N275;
  assign N480 = N231 & N275;
  assign N481 = N233 & N275;
  assign N482 = N235 & N275;
  assign N483 = N237 & N275;
  assign N484 = N239 & N275;
  assign N485 = N241 & N275;
  assign N486 = N243 & N275;
  assign N487 = N245 & N275;
  assign N488 = N247 & N275;
  assign N489 = N249 & N275;
  assign N490 = N251 & N275;
  assign N491 = N253 & N275;
  assign N492 = N255 & N275;
  assign N493 = N257 & N275;
  assign N494 = N259 & N275;
  assign N495 = N261 & N275;
  assign N496 = N263 & N275;
  assign N497 = N265 & N275;
  assign N498 = N267 & N275;
  assign N499 = N269 & N275;
  assign N500 = N271 & N275;
  assign N501 = N273 & N275;
  assign N502 = N212 & N275;
  assign N503 = N214 & N275;
  assign N504 = N216 & N275;
  assign N505 = N218 & N275;
  assign N506 = N220 & N275;
  assign N507 = N222 & N275;
  assign N508 = N224 & N275;
  assign N509 = N226 & N275;
  assign N510 = N228 & N275;
  assign N511 = N230 & N275;
  assign N512 = N232 & N275;
  assign N513 = N234 & N275;
  assign N514 = N236 & N275;
  assign N515 = N238 & N275;
  assign N516 = N240 & N275;
  assign N517 = N242 & N275;
  assign N518 = N244 & N275;
  assign N519 = N246 & N275;
  assign N520 = N248 & N275;
  assign N521 = N250 & N275;
  assign N522 = N252 & N275;
  assign N523 = N254 & N275;
  assign N524 = N256 & N275;
  assign N525 = N258 & N275;
  assign N526 = N260 & N275;
  assign N527 = N262 & N275;
  assign N528 = N264 & N275;
  assign N529 = N266 & N275;
  assign N530 = N268 & N275;
  assign N531 = N270 & N275;
  assign N532 = N272 & N275;
  assign N533 = N274 & N275;
  assign N536 = ~bht_update_i[4];
  assign N537 = ~bht_update_i[5];
  assign N538 = N536 & N537;
  assign N539 = N536 & bht_update_i[5];
  assign N540 = bht_update_i[4] & N537;
  assign N541 = bht_update_i[4] & bht_update_i[5];
  assign N542 = ~bht_update_i[6];
  assign N543 = N538 & N542;
  assign N544 = N538 & bht_update_i[6];
  assign N545 = N540 & N542;
  assign N546 = N540 & bht_update_i[6];
  assign N547 = N539 & N542;
  assign N548 = N539 & bht_update_i[6];
  assign N549 = N541 & N542;
  assign N550 = N541 & bht_update_i[6];
  assign N551 = ~bht_update_i[7];
  assign N552 = N543 & N551;
  assign N553 = N543 & bht_update_i[7];
  assign N554 = N545 & N551;
  assign N555 = N545 & bht_update_i[7];
  assign N556 = N547 & N551;
  assign N557 = N547 & bht_update_i[7];
  assign N558 = N549 & N551;
  assign N559 = N549 & bht_update_i[7];
  assign N560 = N544 & N551;
  assign N561 = N544 & bht_update_i[7];
  assign N562 = N546 & N551;
  assign N563 = N546 & bht_update_i[7];
  assign N564 = N548 & N551;
  assign N565 = N548 & bht_update_i[7];
  assign N566 = N550 & N551;
  assign N567 = N550 & bht_update_i[7];
  assign N568 = ~bht_update_i[8];
  assign N569 = N552 & N568;
  assign N570 = N552 & bht_update_i[8];
  assign N571 = N554 & N568;
  assign N572 = N554 & bht_update_i[8];
  assign N573 = N556 & N568;
  assign N574 = N556 & bht_update_i[8];
  assign N575 = N558 & N568;
  assign N576 = N558 & bht_update_i[8];
  assign N577 = N560 & N568;
  assign N578 = N560 & bht_update_i[8];
  assign N579 = N562 & N568;
  assign N580 = N562 & bht_update_i[8];
  assign N581 = N564 & N568;
  assign N582 = N564 & bht_update_i[8];
  assign N583 = N566 & N568;
  assign N584 = N566 & bht_update_i[8];
  assign N585 = N553 & N568;
  assign N586 = N553 & bht_update_i[8];
  assign N587 = N555 & N568;
  assign N588 = N555 & bht_update_i[8];
  assign N589 = N557 & N568;
  assign N590 = N557 & bht_update_i[8];
  assign N591 = N559 & N568;
  assign N592 = N559 & bht_update_i[8];
  assign N593 = N561 & N568;
  assign N594 = N561 & bht_update_i[8];
  assign N595 = N563 & N568;
  assign N596 = N563 & bht_update_i[8];
  assign N597 = N565 & N568;
  assign N598 = N565 & bht_update_i[8];
  assign N599 = N567 & N568;
  assign N600 = N567 & bht_update_i[8];
  assign N601 = ~bht_update_i[9];
  assign N602 = N569 & N601;
  assign N603 = N569 & bht_update_i[9];
  assign N604 = N571 & N601;
  assign N605 = N571 & bht_update_i[9];
  assign N606 = N573 & N601;
  assign N607 = N573 & bht_update_i[9];
  assign N608 = N575 & N601;
  assign N609 = N575 & bht_update_i[9];
  assign N610 = N577 & N601;
  assign N611 = N577 & bht_update_i[9];
  assign N612 = N579 & N601;
  assign N613 = N579 & bht_update_i[9];
  assign N614 = N581 & N601;
  assign N615 = N581 & bht_update_i[9];
  assign N616 = N583 & N601;
  assign N617 = N583 & bht_update_i[9];
  assign N618 = N585 & N601;
  assign N619 = N585 & bht_update_i[9];
  assign N620 = N587 & N601;
  assign N621 = N587 & bht_update_i[9];
  assign N622 = N589 & N601;
  assign N623 = N589 & bht_update_i[9];
  assign N624 = N591 & N601;
  assign N625 = N591 & bht_update_i[9];
  assign N626 = N593 & N601;
  assign N627 = N593 & bht_update_i[9];
  assign N628 = N595 & N601;
  assign N629 = N595 & bht_update_i[9];
  assign N630 = N597 & N601;
  assign N631 = N597 & bht_update_i[9];
  assign N632 = N599 & N601;
  assign N633 = N599 & bht_update_i[9];
  assign N634 = N570 & N601;
  assign N635 = N570 & bht_update_i[9];
  assign N636 = N572 & N601;
  assign N637 = N572 & bht_update_i[9];
  assign N638 = N574 & N601;
  assign N639 = N574 & bht_update_i[9];
  assign N640 = N576 & N601;
  assign N641 = N576 & bht_update_i[9];
  assign N642 = N578 & N601;
  assign N643 = N578 & bht_update_i[9];
  assign N644 = N580 & N601;
  assign N645 = N580 & bht_update_i[9];
  assign N646 = N582 & N601;
  assign N647 = N582 & bht_update_i[9];
  assign N648 = N584 & N601;
  assign N649 = N584 & bht_update_i[9];
  assign N650 = N586 & N601;
  assign N651 = N586 & bht_update_i[9];
  assign N652 = N588 & N601;
  assign N653 = N588 & bht_update_i[9];
  assign N654 = N590 & N601;
  assign N655 = N590 & bht_update_i[9];
  assign N656 = N592 & N601;
  assign N657 = N592 & bht_update_i[9];
  assign N658 = N594 & N601;
  assign N659 = N594 & bht_update_i[9];
  assign N660 = N596 & N601;
  assign N661 = N596 & bht_update_i[9];
  assign N662 = N598 & N601;
  assign N663 = N598 & bht_update_i[9];
  assign N664 = N600 & N601;
  assign N665 = N600 & bht_update_i[9];
  assign N666 = ~bht_update_i[10];
  assign N667 = N602 & N666;
  assign N668 = N602 & bht_update_i[10];
  assign N669 = N604 & N666;
  assign N670 = N604 & bht_update_i[10];
  assign N671 = N606 & N666;
  assign N672 = N606 & bht_update_i[10];
  assign N673 = N608 & N666;
  assign N674 = N608 & bht_update_i[10];
  assign N675 = N610 & N666;
  assign N676 = N610 & bht_update_i[10];
  assign N677 = N612 & N666;
  assign N678 = N612 & bht_update_i[10];
  assign N679 = N614 & N666;
  assign N680 = N614 & bht_update_i[10];
  assign N681 = N616 & N666;
  assign N682 = N616 & bht_update_i[10];
  assign N683 = N618 & N666;
  assign N684 = N618 & bht_update_i[10];
  assign N685 = N620 & N666;
  assign N686 = N620 & bht_update_i[10];
  assign N687 = N622 & N666;
  assign N688 = N622 & bht_update_i[10];
  assign N689 = N624 & N666;
  assign N690 = N624 & bht_update_i[10];
  assign N691 = N626 & N666;
  assign N692 = N626 & bht_update_i[10];
  assign N693 = N628 & N666;
  assign N694 = N628 & bht_update_i[10];
  assign N695 = N630 & N666;
  assign N696 = N630 & bht_update_i[10];
  assign N697 = N632 & N666;
  assign N698 = N632 & bht_update_i[10];
  assign N699 = N634 & N666;
  assign N700 = N634 & bht_update_i[10];
  assign N701 = N636 & N666;
  assign N702 = N636 & bht_update_i[10];
  assign N703 = N638 & N666;
  assign N704 = N638 & bht_update_i[10];
  assign N705 = N640 & N666;
  assign N706 = N640 & bht_update_i[10];
  assign N707 = N642 & N666;
  assign N708 = N642 & bht_update_i[10];
  assign N709 = N644 & N666;
  assign N710 = N644 & bht_update_i[10];
  assign N711 = N646 & N666;
  assign N712 = N646 & bht_update_i[10];
  assign N713 = N648 & N666;
  assign N714 = N648 & bht_update_i[10];
  assign N715 = N650 & N666;
  assign N716 = N650 & bht_update_i[10];
  assign N717 = N652 & N666;
  assign N718 = N652 & bht_update_i[10];
  assign N719 = N654 & N666;
  assign N720 = N654 & bht_update_i[10];
  assign N721 = N656 & N666;
  assign N722 = N656 & bht_update_i[10];
  assign N723 = N658 & N666;
  assign N724 = N658 & bht_update_i[10];
  assign N725 = N660 & N666;
  assign N726 = N660 & bht_update_i[10];
  assign N727 = N662 & N666;
  assign N728 = N662 & bht_update_i[10];
  assign N729 = N664 & N666;
  assign N730 = N664 & bht_update_i[10];
  assign N731 = N603 & N666;
  assign N732 = N603 & bht_update_i[10];
  assign N733 = N605 & N666;
  assign N734 = N605 & bht_update_i[10];
  assign N735 = N607 & N666;
  assign N736 = N607 & bht_update_i[10];
  assign N737 = N609 & N666;
  assign N738 = N609 & bht_update_i[10];
  assign N739 = N611 & N666;
  assign N740 = N611 & bht_update_i[10];
  assign N741 = N613 & N666;
  assign N742 = N613 & bht_update_i[10];
  assign N743 = N615 & N666;
  assign N744 = N615 & bht_update_i[10];
  assign N745 = N617 & N666;
  assign N746 = N617 & bht_update_i[10];
  assign N747 = N619 & N666;
  assign N748 = N619 & bht_update_i[10];
  assign N749 = N621 & N666;
  assign N750 = N621 & bht_update_i[10];
  assign N751 = N623 & N666;
  assign N752 = N623 & bht_update_i[10];
  assign N753 = N625 & N666;
  assign N754 = N625 & bht_update_i[10];
  assign N755 = N627 & N666;
  assign N756 = N627 & bht_update_i[10];
  assign N757 = N629 & N666;
  assign N758 = N629 & bht_update_i[10];
  assign N759 = N631 & N666;
  assign N760 = N631 & bht_update_i[10];
  assign N761 = N633 & N666;
  assign N762 = N633 & bht_update_i[10];
  assign N763 = N635 & N666;
  assign N764 = N635 & bht_update_i[10];
  assign N765 = N637 & N666;
  assign N766 = N637 & bht_update_i[10];
  assign N767 = N639 & N666;
  assign N768 = N639 & bht_update_i[10];
  assign N769 = N641 & N666;
  assign N770 = N641 & bht_update_i[10];
  assign N771 = N643 & N666;
  assign N772 = N643 & bht_update_i[10];
  assign N773 = N645 & N666;
  assign N774 = N645 & bht_update_i[10];
  assign N775 = N647 & N666;
  assign N776 = N647 & bht_update_i[10];
  assign N777 = N649 & N666;
  assign N778 = N649 & bht_update_i[10];
  assign N779 = N651 & N666;
  assign N780 = N651 & bht_update_i[10];
  assign N781 = N653 & N666;
  assign N782 = N653 & bht_update_i[10];
  assign N783 = N655 & N666;
  assign N784 = N655 & bht_update_i[10];
  assign N785 = N657 & N666;
  assign N786 = N657 & bht_update_i[10];
  assign N787 = N659 & N666;
  assign N788 = N659 & bht_update_i[10];
  assign N789 = N661 & N666;
  assign N790 = N661 & bht_update_i[10];
  assign N791 = N663 & N666;
  assign N792 = N663 & bht_update_i[10];
  assign N793 = N665 & N666;
  assign N794 = N665 & bht_update_i[10];
  assign N797 = bht_update_i[66] & N3564;
  assign N3564 = ~debug_mode_i;
  assign N798 = ~N797;
  assign N799 = N797;
  assign N928 = ~N800;
  assign N929 = ~N801;
  assign N930 = ~N802;
  assign N931 = ~N803;
  assign N932 = ~N804;
  assign N933 = ~N805;
  assign N934 = ~N806;
  assign N935 = ~N807;
  assign N936 = ~N808;
  assign N937 = ~N809;
  assign N938 = ~N810;
  assign N939 = ~N811;
  assign N940 = ~N812;
  assign N941 = ~N813;
  assign N942 = ~N814;
  assign N943 = ~N815;
  assign N944 = ~N816;
  assign N945 = ~N817;
  assign N946 = ~N818;
  assign N947 = ~N819;
  assign N948 = ~N820;
  assign N949 = ~N821;
  assign N950 = ~N822;
  assign N951 = ~N823;
  assign N952 = ~N824;
  assign N953 = ~N825;
  assign N954 = ~N826;
  assign N955 = ~N827;
  assign N956 = ~N828;
  assign N957 = ~N829;
  assign N958 = ~N830;
  assign N959 = ~N831;
  assign N960 = ~N832;
  assign N961 = ~N833;
  assign N962 = ~N834;
  assign N963 = ~N835;
  assign N964 = ~N836;
  assign N965 = ~N837;
  assign N966 = ~N838;
  assign N967 = ~N839;
  assign N968 = ~N840;
  assign N969 = ~N841;
  assign N970 = ~N842;
  assign N971 = ~N843;
  assign N972 = ~N844;
  assign N973 = ~N845;
  assign N974 = ~N846;
  assign N975 = ~N847;
  assign N976 = ~N848;
  assign N977 = ~N849;
  assign N978 = ~N850;
  assign N979 = ~N851;
  assign N980 = ~N852;
  assign N981 = ~N853;
  assign N982 = ~N854;
  assign N983 = ~N855;
  assign N984 = ~N856;
  assign N985 = ~N857;
  assign N986 = ~N858;
  assign N987 = ~N859;
  assign N988 = ~N860;
  assign N989 = ~N861;
  assign N990 = ~N862;
  assign N991 = ~N863;
  assign N992 = ~N864;
  assign N993 = ~N865;
  assign N994 = ~N866;
  assign N995 = ~N867;
  assign N996 = ~N868;
  assign N997 = ~N869;
  assign N998 = ~N870;
  assign N999 = ~N871;
  assign N1000 = ~N872;
  assign N1001 = ~N873;
  assign N1002 = ~N874;
  assign N1003 = ~N875;
  assign N1004 = ~N876;
  assign N1005 = ~N877;
  assign N1006 = ~N878;
  assign N1007 = ~N879;
  assign N1008 = ~N880;
  assign N1009 = ~N881;
  assign N1010 = ~N882;
  assign N1011 = ~N883;
  assign N1012 = ~N884;
  assign N1013 = ~N885;
  assign N1014 = ~N886;
  assign N1015 = ~N887;
  assign N1016 = ~N888;
  assign N1017 = ~N889;
  assign N1018 = ~N890;
  assign N1019 = ~N891;
  assign N1020 = ~N892;
  assign N1021 = ~N893;
  assign N1022 = ~N894;
  assign N1023 = ~N895;
  assign N1024 = ~N896;
  assign N1025 = ~N897;
  assign N1026 = ~N898;
  assign N1027 = ~N899;
  assign N1028 = ~N900;
  assign N1029 = ~N901;
  assign N1030 = ~N902;
  assign N1031 = ~N903;
  assign N1032 = ~N904;
  assign N1033 = ~N905;
  assign N1034 = ~N906;
  assign N1035 = ~N907;
  assign N1036 = ~N908;
  assign N1037 = ~N909;
  assign N1038 = ~N910;
  assign N1039 = ~N911;
  assign N1040 = ~N912;
  assign N1041 = ~N913;
  assign N1042 = ~N914;
  assign N1043 = ~N915;
  assign N1044 = ~N916;
  assign N1045 = ~N917;
  assign N1046 = ~N918;
  assign N1047 = ~N919;
  assign N1048 = ~N920;
  assign N1049 = ~N921;
  assign N1050 = ~N922;
  assign N1051 = ~N923;
  assign N1052 = ~N924;
  assign N1053 = ~N925;
  assign N1054 = ~N926;
  assign N1055 = ~N927;
  assign N1056 = N3526 | N3524;
  assign N1057 = bht_update_i[0] | N1056;
  assign N1058 = ~N1057;
  assign N1059 = N799 & N3524;
  assign N1060 = ~bht_update_i[0];
  assign N1575 = N799 & N2865;
  assign N1576 = ~bht_update_i[0];
  assign N2091 = N799 & N2867;
  assign N2864 = ~N3524;
  assign N2865 = N3526 & N2864;
  assign N2866 = N2864 & N3525;
  assign N2867 = bht_update_i[0] & N2866;
  assign N2868 = ~rst_ni;
  assign N2869 = ~flush_i;
  assign N3126 = N797 & N2869;
  assign N3127 = N1055 & N3126;
  assign N3128 = N798 & N2869;
  assign N3129 = N3127 | N3128;
  assign N3130 = ~N3129;
  assign N3131 = N798 & N2869;
  assign N3132 = ~N3131;
  assign N3133 = N798 & N2869;
  assign N3134 = ~N3133;
  assign N3135 = N797 & N2869;
  assign N3136 = N1054 & N3135;
  assign N3137 = N798 & N2869;
  assign N3138 = N3136 | N3137;
  assign N3139 = ~N3138;
  assign N3140 = ~N3137;
  assign N3141 = N1053 & N3135;
  assign N3142 = N3141 | N3137;
  assign N3143 = ~N3142;
  assign N3144 = N1052 & N3135;
  assign N3145 = N3144 | N3137;
  assign N3146 = ~N3145;
  assign N3147 = N1051 & N3135;
  assign N3148 = N3147 | N3137;
  assign N3149 = ~N3148;
  assign N3150 = N1050 & N3135;
  assign N3151 = N3150 | N3137;
  assign N3152 = ~N3151;
  assign N3153 = N1049 & N3135;
  assign N3154 = N3153 | N3137;
  assign N3155 = ~N3154;
  assign N3156 = N1048 & N3135;
  assign N3157 = N3156 | N3137;
  assign N3158 = ~N3157;
  assign N3159 = N1047 & N3135;
  assign N3160 = N3159 | N3137;
  assign N3161 = ~N3160;
  assign N3162 = N1046 & N3135;
  assign N3163 = N3162 | N3137;
  assign N3164 = ~N3163;
  assign N3165 = N1045 & N3135;
  assign N3166 = N3165 | N3137;
  assign N3167 = ~N3166;
  assign N3168 = N1044 & N3135;
  assign N3169 = N3168 | N3137;
  assign N3170 = ~N3169;
  assign N3171 = N1043 & N3135;
  assign N3172 = N3171 | N3137;
  assign N3173 = ~N3172;
  assign N3174 = N1042 & N3135;
  assign N3175 = N3174 | N3137;
  assign N3176 = ~N3175;
  assign N3177 = N1041 & N3135;
  assign N3178 = N3177 | N3137;
  assign N3179 = ~N3178;
  assign N3180 = N1040 & N3135;
  assign N3181 = N3180 | N3137;
  assign N3182 = ~N3181;
  assign N3183 = N1039 & N3135;
  assign N3184 = N3183 | N3137;
  assign N3185 = ~N3184;
  assign N3186 = N1038 & N3135;
  assign N3187 = N3186 | N3137;
  assign N3188 = ~N3187;
  assign N3189 = N1037 & N3135;
  assign N3190 = N3189 | N3137;
  assign N3191 = ~N3190;
  assign N3192 = N1036 & N3135;
  assign N3193 = N3192 | N3137;
  assign N3194 = ~N3193;
  assign N3195 = N1035 & N3135;
  assign N3196 = N3195 | N3137;
  assign N3197 = ~N3196;
  assign N3198 = N1034 & N3135;
  assign N3199 = N3198 | N3137;
  assign N3200 = ~N3199;
  assign N3201 = N1033 & N3135;
  assign N3202 = N3201 | N3137;
  assign N3203 = ~N3202;
  assign N3204 = N1032 & N3135;
  assign N3205 = N3204 | N3137;
  assign N3206 = ~N3205;
  assign N3207 = N1031 & N3135;
  assign N3208 = N3207 | N3137;
  assign N3209 = ~N3208;
  assign N3210 = N1030 & N3135;
  assign N3211 = N3210 | N3137;
  assign N3212 = ~N3211;
  assign N3213 = N1029 & N3135;
  assign N3214 = N3213 | N3137;
  assign N3215 = ~N3214;
  assign N3216 = N1028 & N3135;
  assign N3217 = N3216 | N3137;
  assign N3218 = ~N3217;
  assign N3219 = N1027 & N3135;
  assign N3220 = N3219 | N3137;
  assign N3221 = ~N3220;
  assign N3222 = N1026 & N3126;
  assign N3223 = N3222 | N3133;
  assign N3224 = ~N3223;
  assign N3225 = N1025 & N3126;
  assign N3226 = N3225 | N3133;
  assign N3227 = ~N3226;
  assign N3228 = N1024 & N3126;
  assign N3229 = N3228 | N3133;
  assign N3230 = ~N3229;
  assign N3231 = N1023 & N3126;
  assign N3232 = N3231 | N3133;
  assign N3233 = ~N3232;
  assign N3234 = N1022 & N3126;
  assign N3235 = N3234 | N3133;
  assign N3236 = ~N3235;
  assign N3237 = N1021 & N3126;
  assign N3238 = N3237 | N3133;
  assign N3239 = ~N3238;
  assign N3240 = N1020 & N3126;
  assign N3241 = N3240 | N3133;
  assign N3242 = ~N3241;
  assign N3243 = N1019 & N3126;
  assign N3244 = N3243 | N3133;
  assign N3245 = ~N3244;
  assign N3246 = N1018 & N3126;
  assign N3247 = N3246 | N3133;
  assign N3248 = ~N3247;
  assign N3249 = N1017 & N3126;
  assign N3250 = N3249 | N3133;
  assign N3251 = ~N3250;
  assign N3252 = N1016 & N3126;
  assign N3253 = N3252 | N3133;
  assign N3254 = ~N3253;
  assign N3255 = N1015 & N3126;
  assign N3256 = N3255 | N3133;
  assign N3257 = ~N3256;
  assign N3258 = N1014 & N3126;
  assign N3259 = N3258 | N3133;
  assign N3260 = ~N3259;
  assign N3261 = N1013 & N3126;
  assign N3262 = N3261 | N3133;
  assign N3263 = ~N3262;
  assign N3264 = N1012 & N3126;
  assign N3265 = N3264 | N3133;
  assign N3266 = ~N3265;
  assign N3267 = N1011 & N3126;
  assign N3268 = N3267 | N3133;
  assign N3269 = ~N3268;
  assign N3270 = N1010 & N3126;
  assign N3271 = N3270 | N3133;
  assign N3272 = ~N3271;
  assign N3273 = N1009 & N3126;
  assign N3274 = N3273 | N3133;
  assign N3275 = ~N3274;
  assign N3276 = N1008 & N3126;
  assign N3277 = N3276 | N3133;
  assign N3278 = ~N3277;
  assign N3279 = N1007 & N3126;
  assign N3280 = N3279 | N3133;
  assign N3281 = ~N3280;
  assign N3282 = N1006 & N3126;
  assign N3283 = N3282 | N3133;
  assign N3284 = ~N3283;
  assign N3285 = N1005 & N3126;
  assign N3286 = N3285 | N3133;
  assign N3287 = ~N3286;
  assign N3288 = N1004 & N3126;
  assign N3289 = N3288 | N3133;
  assign N3290 = ~N3289;
  assign N3291 = N1003 & N3126;
  assign N3292 = N3291 | N3133;
  assign N3293 = ~N3292;
  assign N3294 = N1002 & N3126;
  assign N3295 = N3294 | N3133;
  assign N3296 = ~N3295;
  assign N3297 = N1001 & N3126;
  assign N3298 = N3297 | N3133;
  assign N3299 = ~N3298;
  assign N3300 = N1000 & N3126;
  assign N3301 = N3300 | N3133;
  assign N3302 = ~N3301;
  assign N3303 = N999 & N3126;
  assign N3304 = N3303 | N3133;
  assign N3305 = ~N3304;
  assign N3306 = N998 & N3126;
  assign N3307 = N3306 | N3133;
  assign N3308 = ~N3307;
  assign N3309 = N997 & N3126;
  assign N3310 = N3309 | N3133;
  assign N3311 = ~N3310;
  assign N3312 = N996 & N3126;
  assign N3313 = N3312 | N3133;
  assign N3314 = ~N3313;
  assign N3315 = N995 & N3126;
  assign N3316 = N3315 | N3133;
  assign N3317 = ~N3316;
  assign N3318 = N994 & N3126;
  assign N3319 = N3318 | N3133;
  assign N3320 = ~N3319;
  assign N3321 = N993 & N3126;
  assign N3322 = N3321 | N3131;
  assign N3323 = ~N3322;
  assign N3324 = N992 & N3126;
  assign N3325 = N3324 | N3131;
  assign N3326 = ~N3325;
  assign N3327 = N991 & N3126;
  assign N3328 = N3327 | N3131;
  assign N3329 = ~N3328;
  assign N3330 = N990 & N3126;
  assign N3331 = N3330 | N3131;
  assign N3332 = ~N3331;
  assign N3333 = N989 & N3126;
  assign N3334 = N3333 | N3131;
  assign N3335 = ~N3334;
  assign N3336 = N988 & N3126;
  assign N3337 = N3336 | N3131;
  assign N3338 = ~N3337;
  assign N3339 = N987 & N3126;
  assign N3340 = N3339 | N3131;
  assign N3341 = ~N3340;
  assign N3342 = N986 & N3126;
  assign N3343 = N3342 | N3131;
  assign N3344 = ~N3343;
  assign N3345 = N985 & N3126;
  assign N3346 = N3345 | N3131;
  assign N3347 = ~N3346;
  assign N3348 = N984 & N3126;
  assign N3349 = N3348 | N3131;
  assign N3350 = ~N3349;
  assign N3351 = N983 & N3126;
  assign N3352 = N3351 | N3131;
  assign N3353 = ~N3352;
  assign N3354 = N982 & N3126;
  assign N3355 = N3354 | N3131;
  assign N3356 = ~N3355;
  assign N3357 = N981 & N3126;
  assign N3358 = N3357 | N3131;
  assign N3359 = ~N3358;
  assign N3360 = N980 & N3126;
  assign N3361 = N3360 | N3131;
  assign N3362 = ~N3361;
  assign N3363 = N979 & N3126;
  assign N3364 = N3363 | N3131;
  assign N3365 = ~N3364;
  assign N3366 = N978 & N3126;
  assign N3367 = N3366 | N3131;
  assign N3368 = ~N3367;
  assign N3369 = N977 & N3126;
  assign N3370 = N3369 | N3131;
  assign N3371 = ~N3370;
  assign N3372 = N976 & N3126;
  assign N3373 = N3372 | N3131;
  assign N3374 = ~N3373;
  assign N3375 = N975 & N3126;
  assign N3376 = N3375 | N3131;
  assign N3377 = ~N3376;
  assign N3378 = N974 & N3126;
  assign N3379 = N3378 | N3131;
  assign N3380 = ~N3379;
  assign N3381 = N973 & N3126;
  assign N3382 = N3381 | N3131;
  assign N3383 = ~N3382;
  assign N3384 = N972 & N3126;
  assign N3385 = N3384 | N3131;
  assign N3386 = ~N3385;
  assign N3387 = N971 & N3126;
  assign N3388 = N3387 | N3131;
  assign N3389 = ~N3388;
  assign N3390 = N970 & N3126;
  assign N3391 = N3390 | N3131;
  assign N3392 = ~N3391;
  assign N3393 = N969 & N3126;
  assign N3394 = N3393 | N3131;
  assign N3395 = ~N3394;
  assign N3396 = N968 & N3126;
  assign N3397 = N3396 | N3131;
  assign N3398 = ~N3397;
  assign N3399 = N967 & N3126;
  assign N3400 = N3399 | N3131;
  assign N3401 = ~N3400;
  assign N3402 = N966 & N3126;
  assign N3403 = N3402 | N3131;
  assign N3404 = ~N3403;
  assign N3405 = N965 & N3126;
  assign N3406 = N3405 | N3131;
  assign N3407 = ~N3406;
  assign N3408 = N964 & N3126;
  assign N3409 = N3408 | N3131;
  assign N3410 = ~N3409;
  assign N3411 = N963 & N3126;
  assign N3412 = N3411 | N3131;
  assign N3413 = ~N3412;
  assign N3414 = N962 & N3126;
  assign N3415 = N3414 | N3131;
  assign N3416 = ~N3415;
  assign N3417 = N961 & N3126;
  assign N3418 = N3417 | N3131;
  assign N3419 = ~N3418;
  assign N3420 = N960 & N3126;
  assign N3421 = N3420 | N3128;
  assign N3422 = ~N3421;
  assign N3423 = ~N3128;
  assign N3424 = N959 & N3126;
  assign N3425 = N3424 | N3128;
  assign N3426 = ~N3425;
  assign N3427 = N958 & N3126;
  assign N3428 = N3427 | N3128;
  assign N3429 = ~N3428;
  assign N3430 = N957 & N3126;
  assign N3431 = N3430 | N3128;
  assign N3432 = ~N3431;
  assign N3433 = N956 & N3126;
  assign N3434 = N3433 | N3128;
  assign N3435 = ~N3434;
  assign N3436 = N955 & N3126;
  assign N3437 = N3436 | N3128;
  assign N3438 = ~N3437;
  assign N3439 = N954 & N3126;
  assign N3440 = N3439 | N3128;
  assign N3441 = ~N3440;
  assign N3442 = N953 & N3126;
  assign N3443 = N3442 | N3128;
  assign N3444 = ~N3443;
  assign N3445 = N952 & N3126;
  assign N3446 = N3445 | N3128;
  assign N3447 = ~N3446;
  assign N3448 = N951 & N3126;
  assign N3449 = N3448 | N3128;
  assign N3450 = ~N3449;
  assign N3451 = N950 & N3126;
  assign N3452 = N3451 | N3128;
  assign N3453 = ~N3452;
  assign N3454 = N949 & N3126;
  assign N3455 = N3454 | N3128;
  assign N3456 = ~N3455;
  assign N3457 = N948 & N3126;
  assign N3458 = N3457 | N3128;
  assign N3459 = ~N3458;
  assign N3460 = N947 & N3126;
  assign N3461 = N3460 | N3128;
  assign N3462 = ~N3461;
  assign N3463 = N946 & N3126;
  assign N3464 = N3463 | N3128;
  assign N3465 = ~N3464;
  assign N3466 = N945 & N3126;
  assign N3467 = N3466 | N3128;
  assign N3468 = ~N3467;
  assign N3469 = N944 & N3126;
  assign N3470 = N3469 | N3128;
  assign N3471 = ~N3470;
  assign N3472 = N943 & N3126;
  assign N3473 = N3472 | N3128;
  assign N3474 = ~N3473;
  assign N3475 = N942 & N3126;
  assign N3476 = N3475 | N3128;
  assign N3477 = ~N3476;
  assign N3478 = N941 & N3126;
  assign N3479 = N3478 | N3128;
  assign N3480 = ~N3479;
  assign N3481 = N940 & N3126;
  assign N3482 = N3481 | N3128;
  assign N3483 = ~N3482;
  assign N3484 = N939 & N3126;
  assign N3485 = N3484 | N3128;
  assign N3486 = ~N3485;
  assign N3487 = N938 & N3126;
  assign N3488 = N3487 | N3128;
  assign N3489 = ~N3488;
  assign N3490 = N937 & N3126;
  assign N3491 = N3490 | N3128;
  assign N3492 = ~N3491;
  assign N3493 = N936 & N3126;
  assign N3494 = N3493 | N3128;
  assign N3495 = ~N3494;
  assign N3496 = N935 & N3126;
  assign N3497 = N3496 | N3128;
  assign N3498 = ~N3497;
  assign N3499 = N934 & N3126;
  assign N3500 = N3499 | N3128;
  assign N3501 = ~N3500;
  assign N3502 = N933 & N3126;
  assign N3503 = N3502 | N3128;
  assign N3504 = ~N3503;
  assign N3505 = N932 & N3126;
  assign N3506 = N3505 | N3128;
  assign N3507 = ~N3506;
  assign N3508 = N931 & N3126;
  assign N3509 = N3508 | N3128;
  assign N3510 = ~N3509;
  assign N3511 = N930 & N3126;
  assign N3512 = N3511 | N3128;
  assign N3513 = ~N3512;
  assign N3514 = N929 & N3126;
  assign N3515 = N3514 | N3128;
  assign N3516 = ~N3515;
  assign N3517 = N928 & N3126;
  assign N3518 = N3517 | N3128;
  assign N3519 = ~N3518;

endmodule