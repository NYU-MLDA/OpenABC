module Queue_19
(
  clk,
  reset,
  io_enq_ready,
  io_enq_valid,
  io_enq_bits_addr,
  io_enq_bits_tag,
  io_enq_bits_cmd,
  io_enq_bits_typ,
  io_enq_bits_kill,
  io_enq_bits_phys,
  io_enq_bits_sdq_id,
  io_deq_ready,
  io_deq_valid,
  io_deq_bits_addr,
  io_deq_bits_tag,
  io_deq_bits_cmd,
  io_deq_bits_typ,
  io_deq_bits_kill,
  io_deq_bits_phys,
  io_deq_bits_sdq_id,
  io_count
);

  input [39:0] io_enq_bits_addr;
  input [9:0] io_enq_bits_tag;
  input [4:0] io_enq_bits_cmd;
  input [2:0] io_enq_bits_typ;
  input [4:0] io_enq_bits_sdq_id;
  output [39:0] io_deq_bits_addr;
  output [9:0] io_deq_bits_tag;
  output [4:0] io_deq_bits_cmd;
  output [2:0] io_deq_bits_typ;
  output [4:0] io_deq_bits_sdq_id;
  output [4:0] io_count;
  input clk;
  input reset;
  input io_enq_valid;
  input io_enq_bits_kill;
  input io_enq_bits_phys;
  input io_deq_ready;
  output io_enq_ready;
  output io_deq_valid;
  output io_deq_bits_kill;
  output io_deq_bits_phys;
  wire [39:0] io_deq_bits_addr;
  wire [9:0] io_deq_bits_tag;
  wire [4:0] io_deq_bits_cmd,io_deq_bits_sdq_id,io_count;
  wire [2:0] io_deq_bits_typ;
  wire io_enq_ready,io_deq_valid,io_deq_bits_kill,io_deq_bits_phys,N0,N1,N2,N3,N4,N5,
  N6,N7,N8,N9,N10,do_deq,do_enq,ptr_match,T9,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,empty,T27,full,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105;
  wire [3:0] T3,T6;
  reg [3:0] R1,R4;
  reg maybe_full;
  reg [1039:0] ram;
  assign ptr_match = R4 == R1;
  assign T9 = do_enq ^ do_deq;
  assign io_deq_bits_addr[39] = (N27)? ram[64] : 
                                (N29)? ram[129] : 
                                (N31)? ram[194] : 
                                (N33)? ram[259] : 
                                (N35)? ram[324] : 
                                (N37)? ram[389] : 
                                (N39)? ram[454] : 
                                (N41)? ram[519] : 
                                (N28)? ram[584] : 
                                (N30)? ram[649] : 
                                (N32)? ram[714] : 
                                (N34)? ram[779] : 
                                (N36)? ram[844] : 
                                (N38)? ram[909] : 
                                (N40)? ram[974] : 
                                (N42)? ram[1039] : 1'b0;
  assign io_deq_bits_addr[38] = (N27)? ram[63] : 
                                (N29)? ram[128] : 
                                (N31)? ram[193] : 
                                (N33)? ram[258] : 
                                (N35)? ram[323] : 
                                (N37)? ram[388] : 
                                (N39)? ram[453] : 
                                (N41)? ram[518] : 
                                (N28)? ram[583] : 
                                (N30)? ram[648] : 
                                (N32)? ram[713] : 
                                (N34)? ram[778] : 
                                (N36)? ram[843] : 
                                (N38)? ram[908] : 
                                (N40)? ram[973] : 
                                (N42)? ram[1038] : 1'b0;
  assign io_deq_bits_addr[37] = (N27)? ram[62] : 
                                (N29)? ram[127] : 
                                (N31)? ram[192] : 
                                (N33)? ram[257] : 
                                (N35)? ram[322] : 
                                (N37)? ram[387] : 
                                (N39)? ram[452] : 
                                (N41)? ram[517] : 
                                (N28)? ram[582] : 
                                (N30)? ram[647] : 
                                (N32)? ram[712] : 
                                (N34)? ram[777] : 
                                (N36)? ram[842] : 
                                (N38)? ram[907] : 
                                (N40)? ram[972] : 
                                (N42)? ram[1037] : 1'b0;
  assign io_deq_bits_addr[36] = (N27)? ram[61] : 
                                (N29)? ram[126] : 
                                (N31)? ram[191] : 
                                (N33)? ram[256] : 
                                (N35)? ram[321] : 
                                (N37)? ram[386] : 
                                (N39)? ram[451] : 
                                (N41)? ram[516] : 
                                (N28)? ram[581] : 
                                (N30)? ram[646] : 
                                (N32)? ram[711] : 
                                (N34)? ram[776] : 
                                (N36)? ram[841] : 
                                (N38)? ram[906] : 
                                (N40)? ram[971] : 
                                (N42)? ram[1036] : 1'b0;
  assign io_deq_bits_addr[35] = (N27)? ram[60] : 
                                (N29)? ram[125] : 
                                (N31)? ram[190] : 
                                (N33)? ram[255] : 
                                (N35)? ram[320] : 
                                (N37)? ram[385] : 
                                (N39)? ram[450] : 
                                (N41)? ram[515] : 
                                (N28)? ram[580] : 
                                (N30)? ram[645] : 
                                (N32)? ram[710] : 
                                (N34)? ram[775] : 
                                (N36)? ram[840] : 
                                (N38)? ram[905] : 
                                (N40)? ram[970] : 
                                (N42)? ram[1035] : 1'b0;
  assign io_deq_bits_addr[34] = (N27)? ram[59] : 
                                (N29)? ram[124] : 
                                (N31)? ram[189] : 
                                (N33)? ram[254] : 
                                (N35)? ram[319] : 
                                (N37)? ram[384] : 
                                (N39)? ram[449] : 
                                (N41)? ram[514] : 
                                (N28)? ram[579] : 
                                (N30)? ram[644] : 
                                (N32)? ram[709] : 
                                (N34)? ram[774] : 
                                (N36)? ram[839] : 
                                (N38)? ram[904] : 
                                (N40)? ram[969] : 
                                (N42)? ram[1034] : 1'b0;
  assign io_deq_bits_addr[33] = (N27)? ram[58] : 
                                (N29)? ram[123] : 
                                (N31)? ram[188] : 
                                (N33)? ram[253] : 
                                (N35)? ram[318] : 
                                (N37)? ram[383] : 
                                (N39)? ram[448] : 
                                (N41)? ram[513] : 
                                (N28)? ram[578] : 
                                (N30)? ram[643] : 
                                (N32)? ram[708] : 
                                (N34)? ram[773] : 
                                (N36)? ram[838] : 
                                (N38)? ram[903] : 
                                (N40)? ram[968] : 
                                (N42)? ram[1033] : 1'b0;
  assign io_deq_bits_addr[32] = (N27)? ram[57] : 
                                (N29)? ram[122] : 
                                (N31)? ram[187] : 
                                (N33)? ram[252] : 
                                (N35)? ram[317] : 
                                (N37)? ram[382] : 
                                (N39)? ram[447] : 
                                (N41)? ram[512] : 
                                (N28)? ram[577] : 
                                (N30)? ram[642] : 
                                (N32)? ram[707] : 
                                (N34)? ram[772] : 
                                (N36)? ram[837] : 
                                (N38)? ram[902] : 
                                (N40)? ram[967] : 
                                (N42)? ram[1032] : 1'b0;
  assign io_deq_bits_addr[31] = (N27)? ram[56] : 
                                (N29)? ram[121] : 
                                (N31)? ram[186] : 
                                (N33)? ram[251] : 
                                (N35)? ram[316] : 
                                (N37)? ram[381] : 
                                (N39)? ram[446] : 
                                (N41)? ram[511] : 
                                (N28)? ram[576] : 
                                (N30)? ram[641] : 
                                (N32)? ram[706] : 
                                (N34)? ram[771] : 
                                (N36)? ram[836] : 
                                (N38)? ram[901] : 
                                (N40)? ram[966] : 
                                (N42)? ram[1031] : 1'b0;
  assign io_deq_bits_addr[30] = (N27)? ram[55] : 
                                (N29)? ram[120] : 
                                (N31)? ram[185] : 
                                (N33)? ram[250] : 
                                (N35)? ram[315] : 
                                (N37)? ram[380] : 
                                (N39)? ram[445] : 
                                (N41)? ram[510] : 
                                (N28)? ram[575] : 
                                (N30)? ram[640] : 
                                (N32)? ram[705] : 
                                (N34)? ram[770] : 
                                (N36)? ram[835] : 
                                (N38)? ram[900] : 
                                (N40)? ram[965] : 
                                (N42)? ram[1030] : 1'b0;
  assign io_deq_bits_addr[29] = (N27)? ram[54] : 
                                (N29)? ram[119] : 
                                (N31)? ram[184] : 
                                (N33)? ram[249] : 
                                (N35)? ram[314] : 
                                (N37)? ram[379] : 
                                (N39)? ram[444] : 
                                (N41)? ram[509] : 
                                (N28)? ram[574] : 
                                (N30)? ram[639] : 
                                (N32)? ram[704] : 
                                (N34)? ram[769] : 
                                (N36)? ram[834] : 
                                (N38)? ram[899] : 
                                (N40)? ram[964] : 
                                (N42)? ram[1029] : 1'b0;
  assign io_deq_bits_addr[28] = (N27)? ram[53] : 
                                (N29)? ram[118] : 
                                (N31)? ram[183] : 
                                (N33)? ram[248] : 
                                (N35)? ram[313] : 
                                (N37)? ram[378] : 
                                (N39)? ram[443] : 
                                (N41)? ram[508] : 
                                (N28)? ram[573] : 
                                (N30)? ram[638] : 
                                (N32)? ram[703] : 
                                (N34)? ram[768] : 
                                (N36)? ram[833] : 
                                (N38)? ram[898] : 
                                (N40)? ram[963] : 
                                (N42)? ram[1028] : 1'b0;
  assign io_deq_bits_addr[27] = (N27)? ram[52] : 
                                (N29)? ram[117] : 
                                (N31)? ram[182] : 
                                (N33)? ram[247] : 
                                (N35)? ram[312] : 
                                (N37)? ram[377] : 
                                (N39)? ram[442] : 
                                (N41)? ram[507] : 
                                (N28)? ram[572] : 
                                (N30)? ram[637] : 
                                (N32)? ram[702] : 
                                (N34)? ram[767] : 
                                (N36)? ram[832] : 
                                (N38)? ram[897] : 
                                (N40)? ram[962] : 
                                (N42)? ram[1027] : 1'b0;
  assign io_deq_bits_addr[26] = (N27)? ram[51] : 
                                (N29)? ram[116] : 
                                (N31)? ram[181] : 
                                (N33)? ram[246] : 
                                (N35)? ram[311] : 
                                (N37)? ram[376] : 
                                (N39)? ram[441] : 
                                (N41)? ram[506] : 
                                (N28)? ram[571] : 
                                (N30)? ram[636] : 
                                (N32)? ram[701] : 
                                (N34)? ram[766] : 
                                (N36)? ram[831] : 
                                (N38)? ram[896] : 
                                (N40)? ram[961] : 
                                (N42)? ram[1026] : 1'b0;
  assign io_deq_bits_addr[25] = (N27)? ram[50] : 
                                (N29)? ram[115] : 
                                (N31)? ram[180] : 
                                (N33)? ram[245] : 
                                (N35)? ram[310] : 
                                (N37)? ram[375] : 
                                (N39)? ram[440] : 
                                (N41)? ram[505] : 
                                (N28)? ram[570] : 
                                (N30)? ram[635] : 
                                (N32)? ram[700] : 
                                (N34)? ram[765] : 
                                (N36)? ram[830] : 
                                (N38)? ram[895] : 
                                (N40)? ram[960] : 
                                (N42)? ram[1025] : 1'b0;
  assign io_deq_bits_addr[24] = (N27)? ram[49] : 
                                (N29)? ram[114] : 
                                (N31)? ram[179] : 
                                (N33)? ram[244] : 
                                (N35)? ram[309] : 
                                (N37)? ram[374] : 
                                (N39)? ram[439] : 
                                (N41)? ram[504] : 
                                (N28)? ram[569] : 
                                (N30)? ram[634] : 
                                (N32)? ram[699] : 
                                (N34)? ram[764] : 
                                (N36)? ram[829] : 
                                (N38)? ram[894] : 
                                (N40)? ram[959] : 
                                (N42)? ram[1024] : 1'b0;
  assign io_deq_bits_addr[23] = (N27)? ram[48] : 
                                (N29)? ram[113] : 
                                (N31)? ram[178] : 
                                (N33)? ram[243] : 
                                (N35)? ram[308] : 
                                (N37)? ram[373] : 
                                (N39)? ram[438] : 
                                (N41)? ram[503] : 
                                (N28)? ram[568] : 
                                (N30)? ram[633] : 
                                (N32)? ram[698] : 
                                (N34)? ram[763] : 
                                (N36)? ram[828] : 
                                (N38)? ram[893] : 
                                (N40)? ram[958] : 
                                (N42)? ram[1023] : 1'b0;
  assign io_deq_bits_addr[22] = (N27)? ram[47] : 
                                (N29)? ram[112] : 
                                (N31)? ram[177] : 
                                (N33)? ram[242] : 
                                (N35)? ram[307] : 
                                (N37)? ram[372] : 
                                (N39)? ram[437] : 
                                (N41)? ram[502] : 
                                (N28)? ram[567] : 
                                (N30)? ram[632] : 
                                (N32)? ram[697] : 
                                (N34)? ram[762] : 
                                (N36)? ram[827] : 
                                (N38)? ram[892] : 
                                (N40)? ram[957] : 
                                (N42)? ram[1022] : 1'b0;
  assign io_deq_bits_addr[21] = (N27)? ram[46] : 
                                (N29)? ram[111] : 
                                (N31)? ram[176] : 
                                (N33)? ram[241] : 
                                (N35)? ram[306] : 
                                (N37)? ram[371] : 
                                (N39)? ram[436] : 
                                (N41)? ram[501] : 
                                (N28)? ram[566] : 
                                (N30)? ram[631] : 
                                (N32)? ram[696] : 
                                (N34)? ram[761] : 
                                (N36)? ram[826] : 
                                (N38)? ram[891] : 
                                (N40)? ram[956] : 
                                (N42)? ram[1021] : 1'b0;
  assign io_deq_bits_addr[20] = (N27)? ram[45] : 
                                (N29)? ram[110] : 
                                (N31)? ram[175] : 
                                (N33)? ram[240] : 
                                (N35)? ram[305] : 
                                (N37)? ram[370] : 
                                (N39)? ram[435] : 
                                (N41)? ram[500] : 
                                (N28)? ram[565] : 
                                (N30)? ram[630] : 
                                (N32)? ram[695] : 
                                (N34)? ram[760] : 
                                (N36)? ram[825] : 
                                (N38)? ram[890] : 
                                (N40)? ram[955] : 
                                (N42)? ram[1020] : 1'b0;
  assign io_deq_bits_addr[19] = (N27)? ram[44] : 
                                (N29)? ram[109] : 
                                (N31)? ram[174] : 
                                (N33)? ram[239] : 
                                (N35)? ram[304] : 
                                (N37)? ram[369] : 
                                (N39)? ram[434] : 
                                (N41)? ram[499] : 
                                (N28)? ram[564] : 
                                (N30)? ram[629] : 
                                (N32)? ram[694] : 
                                (N34)? ram[759] : 
                                (N36)? ram[824] : 
                                (N38)? ram[889] : 
                                (N40)? ram[954] : 
                                (N42)? ram[1019] : 1'b0;
  assign io_deq_bits_addr[18] = (N27)? ram[43] : 
                                (N29)? ram[108] : 
                                (N31)? ram[173] : 
                                (N33)? ram[238] : 
                                (N35)? ram[303] : 
                                (N37)? ram[368] : 
                                (N39)? ram[433] : 
                                (N41)? ram[498] : 
                                (N28)? ram[563] : 
                                (N30)? ram[628] : 
                                (N32)? ram[693] : 
                                (N34)? ram[758] : 
                                (N36)? ram[823] : 
                                (N38)? ram[888] : 
                                (N40)? ram[953] : 
                                (N42)? ram[1018] : 1'b0;
  assign io_deq_bits_addr[17] = (N27)? ram[42] : 
                                (N29)? ram[107] : 
                                (N31)? ram[172] : 
                                (N33)? ram[237] : 
                                (N35)? ram[302] : 
                                (N37)? ram[367] : 
                                (N39)? ram[432] : 
                                (N41)? ram[497] : 
                                (N28)? ram[562] : 
                                (N30)? ram[627] : 
                                (N32)? ram[692] : 
                                (N34)? ram[757] : 
                                (N36)? ram[822] : 
                                (N38)? ram[887] : 
                                (N40)? ram[952] : 
                                (N42)? ram[1017] : 1'b0;
  assign io_deq_bits_addr[16] = (N27)? ram[41] : 
                                (N29)? ram[106] : 
                                (N31)? ram[171] : 
                                (N33)? ram[236] : 
                                (N35)? ram[301] : 
                                (N37)? ram[366] : 
                                (N39)? ram[431] : 
                                (N41)? ram[496] : 
                                (N28)? ram[561] : 
                                (N30)? ram[626] : 
                                (N32)? ram[691] : 
                                (N34)? ram[756] : 
                                (N36)? ram[821] : 
                                (N38)? ram[886] : 
                                (N40)? ram[951] : 
                                (N42)? ram[1016] : 1'b0;
  assign io_deq_bits_addr[15] = (N27)? ram[40] : 
                                (N29)? ram[105] : 
                                (N31)? ram[170] : 
                                (N33)? ram[235] : 
                                (N35)? ram[300] : 
                                (N37)? ram[365] : 
                                (N39)? ram[430] : 
                                (N41)? ram[495] : 
                                (N28)? ram[560] : 
                                (N30)? ram[625] : 
                                (N32)? ram[690] : 
                                (N34)? ram[755] : 
                                (N36)? ram[820] : 
                                (N38)? ram[885] : 
                                (N40)? ram[950] : 
                                (N42)? ram[1015] : 1'b0;
  assign io_deq_bits_addr[14] = (N27)? ram[39] : 
                                (N29)? ram[104] : 
                                (N31)? ram[169] : 
                                (N33)? ram[234] : 
                                (N35)? ram[299] : 
                                (N37)? ram[364] : 
                                (N39)? ram[429] : 
                                (N41)? ram[494] : 
                                (N28)? ram[559] : 
                                (N30)? ram[624] : 
                                (N32)? ram[689] : 
                                (N34)? ram[754] : 
                                (N36)? ram[819] : 
                                (N38)? ram[884] : 
                                (N40)? ram[949] : 
                                (N42)? ram[1014] : 1'b0;
  assign io_deq_bits_addr[13] = (N27)? ram[38] : 
                                (N29)? ram[103] : 
                                (N31)? ram[168] : 
                                (N33)? ram[233] : 
                                (N35)? ram[298] : 
                                (N37)? ram[363] : 
                                (N39)? ram[428] : 
                                (N41)? ram[493] : 
                                (N28)? ram[558] : 
                                (N30)? ram[623] : 
                                (N32)? ram[688] : 
                                (N34)? ram[753] : 
                                (N36)? ram[818] : 
                                (N38)? ram[883] : 
                                (N40)? ram[948] : 
                                (N42)? ram[1013] : 1'b0;
  assign io_deq_bits_addr[12] = (N27)? ram[37] : 
                                (N29)? ram[102] : 
                                (N31)? ram[167] : 
                                (N33)? ram[232] : 
                                (N35)? ram[297] : 
                                (N37)? ram[362] : 
                                (N39)? ram[427] : 
                                (N41)? ram[492] : 
                                (N28)? ram[557] : 
                                (N30)? ram[622] : 
                                (N32)? ram[687] : 
                                (N34)? ram[752] : 
                                (N36)? ram[817] : 
                                (N38)? ram[882] : 
                                (N40)? ram[947] : 
                                (N42)? ram[1012] : 1'b0;
  assign io_deq_bits_addr[11] = (N27)? ram[36] : 
                                (N29)? ram[101] : 
                                (N31)? ram[166] : 
                                (N33)? ram[231] : 
                                (N35)? ram[296] : 
                                (N37)? ram[361] : 
                                (N39)? ram[426] : 
                                (N41)? ram[491] : 
                                (N28)? ram[556] : 
                                (N30)? ram[621] : 
                                (N32)? ram[686] : 
                                (N34)? ram[751] : 
                                (N36)? ram[816] : 
                                (N38)? ram[881] : 
                                (N40)? ram[946] : 
                                (N42)? ram[1011] : 1'b0;
  assign io_deq_bits_addr[10] = (N27)? ram[35] : 
                                (N29)? ram[100] : 
                                (N31)? ram[165] : 
                                (N33)? ram[230] : 
                                (N35)? ram[295] : 
                                (N37)? ram[360] : 
                                (N39)? ram[425] : 
                                (N41)? ram[490] : 
                                (N28)? ram[555] : 
                                (N30)? ram[620] : 
                                (N32)? ram[685] : 
                                (N34)? ram[750] : 
                                (N36)? ram[815] : 
                                (N38)? ram[880] : 
                                (N40)? ram[945] : 
                                (N42)? ram[1010] : 1'b0;
  assign io_deq_bits_addr[9] = (N27)? ram[34] : 
                               (N29)? ram[99] : 
                               (N31)? ram[164] : 
                               (N33)? ram[229] : 
                               (N35)? ram[294] : 
                               (N37)? ram[359] : 
                               (N39)? ram[424] : 
                               (N41)? ram[489] : 
                               (N28)? ram[554] : 
                               (N30)? ram[619] : 
                               (N32)? ram[684] : 
                               (N34)? ram[749] : 
                               (N36)? ram[814] : 
                               (N38)? ram[879] : 
                               (N40)? ram[944] : 
                               (N42)? ram[1009] : 1'b0;
  assign io_deq_bits_addr[8] = (N27)? ram[33] : 
                               (N29)? ram[98] : 
                               (N31)? ram[163] : 
                               (N33)? ram[228] : 
                               (N35)? ram[293] : 
                               (N37)? ram[358] : 
                               (N39)? ram[423] : 
                               (N41)? ram[488] : 
                               (N28)? ram[553] : 
                               (N30)? ram[618] : 
                               (N32)? ram[683] : 
                               (N34)? ram[748] : 
                               (N36)? ram[813] : 
                               (N38)? ram[878] : 
                               (N40)? ram[943] : 
                               (N42)? ram[1008] : 1'b0;
  assign io_deq_bits_addr[7] = (N27)? ram[32] : 
                               (N29)? ram[97] : 
                               (N31)? ram[162] : 
                               (N33)? ram[227] : 
                               (N35)? ram[292] : 
                               (N37)? ram[357] : 
                               (N39)? ram[422] : 
                               (N41)? ram[487] : 
                               (N28)? ram[552] : 
                               (N30)? ram[617] : 
                               (N32)? ram[682] : 
                               (N34)? ram[747] : 
                               (N36)? ram[812] : 
                               (N38)? ram[877] : 
                               (N40)? ram[942] : 
                               (N42)? ram[1007] : 1'b0;
  assign io_deq_bits_addr[6] = (N27)? ram[31] : 
                               (N29)? ram[96] : 
                               (N31)? ram[161] : 
                               (N33)? ram[226] : 
                               (N35)? ram[291] : 
                               (N37)? ram[356] : 
                               (N39)? ram[421] : 
                               (N41)? ram[486] : 
                               (N28)? ram[551] : 
                               (N30)? ram[616] : 
                               (N32)? ram[681] : 
                               (N34)? ram[746] : 
                               (N36)? ram[811] : 
                               (N38)? ram[876] : 
                               (N40)? ram[941] : 
                               (N42)? ram[1006] : 1'b0;
  assign io_deq_bits_addr[5] = (N27)? ram[30] : 
                               (N29)? ram[95] : 
                               (N31)? ram[160] : 
                               (N33)? ram[225] : 
                               (N35)? ram[290] : 
                               (N37)? ram[355] : 
                               (N39)? ram[420] : 
                               (N41)? ram[485] : 
                               (N28)? ram[550] : 
                               (N30)? ram[615] : 
                               (N32)? ram[680] : 
                               (N34)? ram[745] : 
                               (N36)? ram[810] : 
                               (N38)? ram[875] : 
                               (N40)? ram[940] : 
                               (N42)? ram[1005] : 1'b0;
  assign io_deq_bits_addr[4] = (N27)? ram[29] : 
                               (N29)? ram[94] : 
                               (N31)? ram[159] : 
                               (N33)? ram[224] : 
                               (N35)? ram[289] : 
                               (N37)? ram[354] : 
                               (N39)? ram[419] : 
                               (N41)? ram[484] : 
                               (N28)? ram[549] : 
                               (N30)? ram[614] : 
                               (N32)? ram[679] : 
                               (N34)? ram[744] : 
                               (N36)? ram[809] : 
                               (N38)? ram[874] : 
                               (N40)? ram[939] : 
                               (N42)? ram[1004] : 1'b0;
  assign io_deq_bits_addr[3] = (N27)? ram[28] : 
                               (N29)? ram[93] : 
                               (N31)? ram[158] : 
                               (N33)? ram[223] : 
                               (N35)? ram[288] : 
                               (N37)? ram[353] : 
                               (N39)? ram[418] : 
                               (N41)? ram[483] : 
                               (N28)? ram[548] : 
                               (N30)? ram[613] : 
                               (N32)? ram[678] : 
                               (N34)? ram[743] : 
                               (N36)? ram[808] : 
                               (N38)? ram[873] : 
                               (N40)? ram[938] : 
                               (N42)? ram[1003] : 1'b0;
  assign io_deq_bits_addr[2] = (N27)? ram[27] : 
                               (N29)? ram[92] : 
                               (N31)? ram[157] : 
                               (N33)? ram[222] : 
                               (N35)? ram[287] : 
                               (N37)? ram[352] : 
                               (N39)? ram[417] : 
                               (N41)? ram[482] : 
                               (N28)? ram[547] : 
                               (N30)? ram[612] : 
                               (N32)? ram[677] : 
                               (N34)? ram[742] : 
                               (N36)? ram[807] : 
                               (N38)? ram[872] : 
                               (N40)? ram[937] : 
                               (N42)? ram[1002] : 1'b0;
  assign io_deq_bits_addr[1] = (N27)? ram[26] : 
                               (N29)? ram[91] : 
                               (N31)? ram[156] : 
                               (N33)? ram[221] : 
                               (N35)? ram[286] : 
                               (N37)? ram[351] : 
                               (N39)? ram[416] : 
                               (N41)? ram[481] : 
                               (N28)? ram[546] : 
                               (N30)? ram[611] : 
                               (N32)? ram[676] : 
                               (N34)? ram[741] : 
                               (N36)? ram[806] : 
                               (N38)? ram[871] : 
                               (N40)? ram[936] : 
                               (N42)? ram[1001] : 1'b0;
  assign io_deq_bits_addr[0] = (N27)? ram[25] : 
                               (N29)? ram[90] : 
                               (N31)? ram[155] : 
                               (N33)? ram[220] : 
                               (N35)? ram[285] : 
                               (N37)? ram[350] : 
                               (N39)? ram[415] : 
                               (N41)? ram[480] : 
                               (N28)? ram[545] : 
                               (N30)? ram[610] : 
                               (N32)? ram[675] : 
                               (N34)? ram[740] : 
                               (N36)? ram[805] : 
                               (N38)? ram[870] : 
                               (N40)? ram[935] : 
                               (N42)? ram[1000] : 1'b0;
  assign io_deq_bits_tag[9] = (N27)? ram[24] : 
                              (N29)? ram[89] : 
                              (N31)? ram[154] : 
                              (N33)? ram[219] : 
                              (N35)? ram[284] : 
                              (N37)? ram[349] : 
                              (N39)? ram[414] : 
                              (N41)? ram[479] : 
                              (N28)? ram[544] : 
                              (N30)? ram[609] : 
                              (N32)? ram[674] : 
                              (N34)? ram[739] : 
                              (N36)? ram[804] : 
                              (N38)? ram[869] : 
                              (N40)? ram[934] : 
                              (N42)? ram[999] : 1'b0;
  assign io_deq_bits_tag[8] = (N27)? ram[23] : 
                              (N29)? ram[88] : 
                              (N31)? ram[153] : 
                              (N33)? ram[218] : 
                              (N35)? ram[283] : 
                              (N37)? ram[348] : 
                              (N39)? ram[413] : 
                              (N41)? ram[478] : 
                              (N28)? ram[543] : 
                              (N30)? ram[608] : 
                              (N32)? ram[673] : 
                              (N34)? ram[738] : 
                              (N36)? ram[803] : 
                              (N38)? ram[868] : 
                              (N40)? ram[933] : 
                              (N42)? ram[998] : 1'b0;
  assign io_deq_bits_tag[7] = (N27)? ram[22] : 
                              (N29)? ram[87] : 
                              (N31)? ram[152] : 
                              (N33)? ram[217] : 
                              (N35)? ram[282] : 
                              (N37)? ram[347] : 
                              (N39)? ram[412] : 
                              (N41)? ram[477] : 
                              (N28)? ram[542] : 
                              (N30)? ram[607] : 
                              (N32)? ram[672] : 
                              (N34)? ram[737] : 
                              (N36)? ram[802] : 
                              (N38)? ram[867] : 
                              (N40)? ram[932] : 
                              (N42)? ram[997] : 1'b0;
  assign io_deq_bits_tag[6] = (N27)? ram[21] : 
                              (N29)? ram[86] : 
                              (N31)? ram[151] : 
                              (N33)? ram[216] : 
                              (N35)? ram[281] : 
                              (N37)? ram[346] : 
                              (N39)? ram[411] : 
                              (N41)? ram[476] : 
                              (N28)? ram[541] : 
                              (N30)? ram[606] : 
                              (N32)? ram[671] : 
                              (N34)? ram[736] : 
                              (N36)? ram[801] : 
                              (N38)? ram[866] : 
                              (N40)? ram[931] : 
                              (N42)? ram[996] : 1'b0;
  assign io_deq_bits_tag[5] = (N27)? ram[20] : 
                              (N29)? ram[85] : 
                              (N31)? ram[150] : 
                              (N33)? ram[215] : 
                              (N35)? ram[280] : 
                              (N37)? ram[345] : 
                              (N39)? ram[410] : 
                              (N41)? ram[475] : 
                              (N28)? ram[540] : 
                              (N30)? ram[605] : 
                              (N32)? ram[670] : 
                              (N34)? ram[735] : 
                              (N36)? ram[800] : 
                              (N38)? ram[865] : 
                              (N40)? ram[930] : 
                              (N42)? ram[995] : 1'b0;
  assign io_deq_bits_tag[4] = (N27)? ram[19] : 
                              (N29)? ram[84] : 
                              (N31)? ram[149] : 
                              (N33)? ram[214] : 
                              (N35)? ram[279] : 
                              (N37)? ram[344] : 
                              (N39)? ram[409] : 
                              (N41)? ram[474] : 
                              (N28)? ram[539] : 
                              (N30)? ram[604] : 
                              (N32)? ram[669] : 
                              (N34)? ram[734] : 
                              (N36)? ram[799] : 
                              (N38)? ram[864] : 
                              (N40)? ram[929] : 
                              (N42)? ram[994] : 1'b0;
  assign io_deq_bits_tag[3] = (N27)? ram[18] : 
                              (N29)? ram[83] : 
                              (N31)? ram[148] : 
                              (N33)? ram[213] : 
                              (N35)? ram[278] : 
                              (N37)? ram[343] : 
                              (N39)? ram[408] : 
                              (N41)? ram[473] : 
                              (N28)? ram[538] : 
                              (N30)? ram[603] : 
                              (N32)? ram[668] : 
                              (N34)? ram[733] : 
                              (N36)? ram[798] : 
                              (N38)? ram[863] : 
                              (N40)? ram[928] : 
                              (N42)? ram[993] : 1'b0;
  assign io_deq_bits_tag[2] = (N27)? ram[17] : 
                              (N29)? ram[82] : 
                              (N31)? ram[147] : 
                              (N33)? ram[212] : 
                              (N35)? ram[277] : 
                              (N37)? ram[342] : 
                              (N39)? ram[407] : 
                              (N41)? ram[472] : 
                              (N28)? ram[537] : 
                              (N30)? ram[602] : 
                              (N32)? ram[667] : 
                              (N34)? ram[732] : 
                              (N36)? ram[797] : 
                              (N38)? ram[862] : 
                              (N40)? ram[927] : 
                              (N42)? ram[992] : 1'b0;
  assign io_deq_bits_tag[1] = (N27)? ram[16] : 
                              (N29)? ram[81] : 
                              (N31)? ram[146] : 
                              (N33)? ram[211] : 
                              (N35)? ram[276] : 
                              (N37)? ram[341] : 
                              (N39)? ram[406] : 
                              (N41)? ram[471] : 
                              (N28)? ram[536] : 
                              (N30)? ram[601] : 
                              (N32)? ram[666] : 
                              (N34)? ram[731] : 
                              (N36)? ram[796] : 
                              (N38)? ram[861] : 
                              (N40)? ram[926] : 
                              (N42)? ram[991] : 1'b0;
  assign io_deq_bits_tag[0] = (N27)? ram[15] : 
                              (N29)? ram[80] : 
                              (N31)? ram[145] : 
                              (N33)? ram[210] : 
                              (N35)? ram[275] : 
                              (N37)? ram[340] : 
                              (N39)? ram[405] : 
                              (N41)? ram[470] : 
                              (N28)? ram[535] : 
                              (N30)? ram[600] : 
                              (N32)? ram[665] : 
                              (N34)? ram[730] : 
                              (N36)? ram[795] : 
                              (N38)? ram[860] : 
                              (N40)? ram[925] : 
                              (N42)? ram[990] : 1'b0;
  assign io_deq_bits_cmd[4] = (N27)? ram[14] : 
                              (N29)? ram[79] : 
                              (N31)? ram[144] : 
                              (N33)? ram[209] : 
                              (N35)? ram[274] : 
                              (N37)? ram[339] : 
                              (N39)? ram[404] : 
                              (N41)? ram[469] : 
                              (N28)? ram[534] : 
                              (N30)? ram[599] : 
                              (N32)? ram[664] : 
                              (N34)? ram[729] : 
                              (N36)? ram[794] : 
                              (N38)? ram[859] : 
                              (N40)? ram[924] : 
                              (N42)? ram[989] : 1'b0;
  assign io_deq_bits_cmd[3] = (N27)? ram[13] : 
                              (N29)? ram[78] : 
                              (N31)? ram[143] : 
                              (N33)? ram[208] : 
                              (N35)? ram[273] : 
                              (N37)? ram[338] : 
                              (N39)? ram[403] : 
                              (N41)? ram[468] : 
                              (N28)? ram[533] : 
                              (N30)? ram[598] : 
                              (N32)? ram[663] : 
                              (N34)? ram[728] : 
                              (N36)? ram[793] : 
                              (N38)? ram[858] : 
                              (N40)? ram[923] : 
                              (N42)? ram[988] : 1'b0;
  assign io_deq_bits_cmd[2] = (N27)? ram[12] : 
                              (N29)? ram[77] : 
                              (N31)? ram[142] : 
                              (N33)? ram[207] : 
                              (N35)? ram[272] : 
                              (N37)? ram[337] : 
                              (N39)? ram[402] : 
                              (N41)? ram[467] : 
                              (N28)? ram[532] : 
                              (N30)? ram[597] : 
                              (N32)? ram[662] : 
                              (N34)? ram[727] : 
                              (N36)? ram[792] : 
                              (N38)? ram[857] : 
                              (N40)? ram[922] : 
                              (N42)? ram[987] : 1'b0;
  assign io_deq_bits_cmd[1] = (N27)? ram[11] : 
                              (N29)? ram[76] : 
                              (N31)? ram[141] : 
                              (N33)? ram[206] : 
                              (N35)? ram[271] : 
                              (N37)? ram[336] : 
                              (N39)? ram[401] : 
                              (N41)? ram[466] : 
                              (N28)? ram[531] : 
                              (N30)? ram[596] : 
                              (N32)? ram[661] : 
                              (N34)? ram[726] : 
                              (N36)? ram[791] : 
                              (N38)? ram[856] : 
                              (N40)? ram[921] : 
                              (N42)? ram[986] : 1'b0;
  assign io_deq_bits_cmd[0] = (N27)? ram[10] : 
                              (N29)? ram[75] : 
                              (N31)? ram[140] : 
                              (N33)? ram[205] : 
                              (N35)? ram[270] : 
                              (N37)? ram[335] : 
                              (N39)? ram[400] : 
                              (N41)? ram[465] : 
                              (N28)? ram[530] : 
                              (N30)? ram[595] : 
                              (N32)? ram[660] : 
                              (N34)? ram[725] : 
                              (N36)? ram[790] : 
                              (N38)? ram[855] : 
                              (N40)? ram[920] : 
                              (N42)? ram[985] : 1'b0;
  assign io_deq_bits_typ[2] = (N27)? ram[9] : 
                              (N29)? ram[74] : 
                              (N31)? ram[139] : 
                              (N33)? ram[204] : 
                              (N35)? ram[269] : 
                              (N37)? ram[334] : 
                              (N39)? ram[399] : 
                              (N41)? ram[464] : 
                              (N28)? ram[529] : 
                              (N30)? ram[594] : 
                              (N32)? ram[659] : 
                              (N34)? ram[724] : 
                              (N36)? ram[789] : 
                              (N38)? ram[854] : 
                              (N40)? ram[919] : 
                              (N42)? ram[984] : 1'b0;
  assign io_deq_bits_typ[1] = (N27)? ram[8] : 
                              (N29)? ram[73] : 
                              (N31)? ram[138] : 
                              (N33)? ram[203] : 
                              (N35)? ram[268] : 
                              (N37)? ram[333] : 
                              (N39)? ram[398] : 
                              (N41)? ram[463] : 
                              (N28)? ram[528] : 
                              (N30)? ram[593] : 
                              (N32)? ram[658] : 
                              (N34)? ram[723] : 
                              (N36)? ram[788] : 
                              (N38)? ram[853] : 
                              (N40)? ram[918] : 
                              (N42)? ram[983] : 1'b0;
  assign io_deq_bits_typ[0] = (N27)? ram[7] : 
                              (N29)? ram[72] : 
                              (N31)? ram[137] : 
                              (N33)? ram[202] : 
                              (N35)? ram[267] : 
                              (N37)? ram[332] : 
                              (N39)? ram[397] : 
                              (N41)? ram[462] : 
                              (N28)? ram[527] : 
                              (N30)? ram[592] : 
                              (N32)? ram[657] : 
                              (N34)? ram[722] : 
                              (N36)? ram[787] : 
                              (N38)? ram[852] : 
                              (N40)? ram[917] : 
                              (N42)? ram[982] : 1'b0;
  assign io_deq_bits_kill = (N27)? ram[6] : 
                            (N29)? ram[71] : 
                            (N31)? ram[136] : 
                            (N33)? ram[201] : 
                            (N35)? ram[266] : 
                            (N37)? ram[331] : 
                            (N39)? ram[396] : 
                            (N41)? ram[461] : 
                            (N28)? ram[526] : 
                            (N30)? ram[591] : 
                            (N32)? ram[656] : 
                            (N34)? ram[721] : 
                            (N36)? ram[786] : 
                            (N38)? ram[851] : 
                            (N40)? ram[916] : 
                            (N42)? ram[981] : 1'b0;
  assign io_deq_bits_phys = (N27)? ram[5] : 
                            (N29)? ram[70] : 
                            (N31)? ram[135] : 
                            (N33)? ram[200] : 
                            (N35)? ram[265] : 
                            (N37)? ram[330] : 
                            (N39)? ram[395] : 
                            (N41)? ram[460] : 
                            (N28)? ram[525] : 
                            (N30)? ram[590] : 
                            (N32)? ram[655] : 
                            (N34)? ram[720] : 
                            (N36)? ram[785] : 
                            (N38)? ram[850] : 
                            (N40)? ram[915] : 
                            (N42)? ram[980] : 1'b0;
  assign io_deq_bits_sdq_id[4] = (N27)? ram[4] : 
                                 (N29)? ram[69] : 
                                 (N31)? ram[134] : 
                                 (N33)? ram[199] : 
                                 (N35)? ram[264] : 
                                 (N37)? ram[329] : 
                                 (N39)? ram[394] : 
                                 (N41)? ram[459] : 
                                 (N28)? ram[524] : 
                                 (N30)? ram[589] : 
                                 (N32)? ram[654] : 
                                 (N34)? ram[719] : 
                                 (N36)? ram[784] : 
                                 (N38)? ram[849] : 
                                 (N40)? ram[914] : 
                                 (N42)? ram[979] : 1'b0;
  assign io_deq_bits_sdq_id[3] = (N27)? ram[3] : 
                                 (N29)? ram[68] : 
                                 (N31)? ram[133] : 
                                 (N33)? ram[198] : 
                                 (N35)? ram[263] : 
                                 (N37)? ram[328] : 
                                 (N39)? ram[393] : 
                                 (N41)? ram[458] : 
                                 (N28)? ram[523] : 
                                 (N30)? ram[588] : 
                                 (N32)? ram[653] : 
                                 (N34)? ram[718] : 
                                 (N36)? ram[783] : 
                                 (N38)? ram[848] : 
                                 (N40)? ram[913] : 
                                 (N42)? ram[978] : 1'b0;
  assign io_deq_bits_sdq_id[2] = (N27)? ram[2] : 
                                 (N29)? ram[67] : 
                                 (N31)? ram[132] : 
                                 (N33)? ram[197] : 
                                 (N35)? ram[262] : 
                                 (N37)? ram[327] : 
                                 (N39)? ram[392] : 
                                 (N41)? ram[457] : 
                                 (N28)? ram[522] : 
                                 (N30)? ram[587] : 
                                 (N32)? ram[652] : 
                                 (N34)? ram[717] : 
                                 (N36)? ram[782] : 
                                 (N38)? ram[847] : 
                                 (N40)? ram[912] : 
                                 (N42)? ram[977] : 1'b0;
  assign io_deq_bits_sdq_id[1] = (N27)? ram[1] : 
                                 (N29)? ram[66] : 
                                 (N31)? ram[131] : 
                                 (N33)? ram[196] : 
                                 (N35)? ram[261] : 
                                 (N37)? ram[326] : 
                                 (N39)? ram[391] : 
                                 (N41)? ram[456] : 
                                 (N28)? ram[521] : 
                                 (N30)? ram[586] : 
                                 (N32)? ram[651] : 
                                 (N34)? ram[716] : 
                                 (N36)? ram[781] : 
                                 (N38)? ram[846] : 
                                 (N40)? ram[911] : 
                                 (N42)? ram[976] : 1'b0;
  assign io_deq_bits_sdq_id[0] = (N27)? ram[0] : 
                                 (N29)? ram[65] : 
                                 (N31)? ram[130] : 
                                 (N33)? ram[195] : 
                                 (N35)? ram[260] : 
                                 (N37)? ram[325] : 
                                 (N39)? ram[390] : 
                                 (N41)? ram[455] : 
                                 (N28)? ram[520] : 
                                 (N30)? ram[585] : 
                                 (N32)? ram[650] : 
                                 (N34)? ram[715] : 
                                 (N36)? ram[780] : 
                                 (N38)? ram[845] : 
                                 (N40)? ram[910] : 
                                 (N42)? ram[975] : 1'b0;

  always @(posedge clk) begin
    if(N45) begin
      R1[3] <= N49;
    end 
  end


  always @(posedge clk) begin
    if(N45) begin
      R1[2] <= N48;
    end 
  end


  always @(posedge clk) begin
    if(N45) begin
      R1[1] <= N47;
    end 
  end


  always @(posedge clk) begin
    if(N45) begin
      R1[0] <= N46;
    end 
  end


  always @(posedge clk) begin
    if(N52) begin
      R4[3] <= N56;
    end 
  end


  always @(posedge clk) begin
    if(N52) begin
      R4[2] <= N55;
    end 
  end


  always @(posedge clk) begin
    if(N52) begin
      R4[1] <= N54;
    end 
  end


  always @(posedge clk) begin
    if(N52) begin
      R4[0] <= N53;
    end 
  end


  always @(posedge clk) begin
    if(N59) begin
      maybe_full <= N60;
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1039] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1038] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1037] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1036] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1035] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1034] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1033] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1032] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1031] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1030] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1029] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1028] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1027] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1026] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1025] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1024] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1023] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1022] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1021] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1020] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1019] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1018] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1017] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1016] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1015] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1014] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1013] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1012] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1011] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1010] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1009] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1008] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1007] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1006] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1005] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1004] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1003] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1002] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1001] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[1000] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[999] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[998] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[997] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[996] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[995] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[994] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[993] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[992] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[991] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[990] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[989] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[988] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[987] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[986] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[985] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[984] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[983] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[982] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[981] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[980] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[979] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[978] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[977] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[976] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N93) begin
      ram[975] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[974] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[973] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[972] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[971] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[970] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[969] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[968] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[967] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[966] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[965] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[964] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[963] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[962] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[961] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[960] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[959] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[958] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[957] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[956] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[955] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[954] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[953] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[952] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[951] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[950] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[949] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[948] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[947] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[946] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[945] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[944] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[943] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[942] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[941] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[940] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[939] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[938] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[937] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[936] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[935] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[934] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[933] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[932] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[931] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[930] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[929] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[928] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[927] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[926] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[925] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[924] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[923] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[922] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[921] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[920] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[919] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[918] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[917] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[916] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[915] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[914] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[913] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[912] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[911] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N92) begin
      ram[910] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[909] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[908] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[907] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[906] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[905] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[904] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[903] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[902] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[901] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[900] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[899] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[898] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[897] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[896] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[895] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[894] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[893] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[892] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[891] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[890] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[889] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[888] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[887] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[886] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[885] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[884] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[883] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[882] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[881] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[880] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[879] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[878] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[877] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[876] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[875] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[874] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[873] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[872] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[871] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[870] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[869] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[868] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[867] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[866] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[865] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[864] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[863] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[862] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[861] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[860] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[859] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[858] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[857] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[856] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[855] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[854] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[853] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[852] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[851] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[850] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[849] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[848] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[847] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[846] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N91) begin
      ram[845] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[844] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[843] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[842] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[841] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[840] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[839] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[838] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[837] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[836] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[835] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[834] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[833] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[832] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[831] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[830] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[829] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[828] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[827] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[826] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[825] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[824] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[823] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[822] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[821] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[820] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[819] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[818] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[817] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[816] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[815] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[814] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[813] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[812] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[811] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[810] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[809] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[808] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[807] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[806] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[805] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[804] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[803] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[802] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[801] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[800] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[799] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[798] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[797] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[796] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[795] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[794] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[793] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[792] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[791] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[790] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[789] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[788] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[787] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[786] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[785] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[784] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[783] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[782] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[781] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N90) begin
      ram[780] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[779] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[778] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[777] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[776] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[775] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[774] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[773] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[772] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[771] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[770] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[769] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[768] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[767] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[766] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[765] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[764] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[763] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[762] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[761] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[760] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[759] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[758] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[757] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[756] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[755] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[754] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[753] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[752] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[751] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[750] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[749] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[748] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[747] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[746] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[745] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[744] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[743] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[742] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[741] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[740] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[739] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[738] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[737] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[736] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[735] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[734] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[733] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[732] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[731] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[730] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[729] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[728] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[727] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[726] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[725] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[724] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[723] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[722] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[721] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[720] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[719] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[718] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[717] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[716] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N89) begin
      ram[715] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[714] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[713] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[712] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[711] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[710] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[709] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[708] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[707] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[706] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[705] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[704] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[703] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[702] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[701] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[700] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[699] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[698] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[697] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[696] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[695] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[694] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[693] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[692] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[691] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[690] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[689] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[688] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[687] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[686] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[685] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[684] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[683] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[682] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[681] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[680] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[679] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[678] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[677] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[676] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[675] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[674] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[673] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[672] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[671] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[670] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[669] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[668] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[667] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[666] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[665] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[664] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[663] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[662] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[661] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[660] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[659] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[658] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[657] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[656] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[655] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[654] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[653] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[652] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[651] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N88) begin
      ram[650] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[649] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[648] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[647] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[646] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[645] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[644] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[643] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[642] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[641] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[640] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[639] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[638] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[637] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[636] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[635] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[634] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[633] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[632] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[631] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[630] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[629] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[628] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[627] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[626] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[625] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[624] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[623] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[622] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[621] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[620] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[619] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[618] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[617] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[616] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[615] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[614] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[613] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[612] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[611] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[610] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[609] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[608] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[607] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[606] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[605] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[604] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[603] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[602] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[601] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[600] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[599] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[598] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[597] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[596] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[595] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[594] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[593] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[592] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[591] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[590] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[589] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[588] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[587] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[586] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N87) begin
      ram[585] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[584] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[583] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[582] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[581] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[580] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[579] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[578] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[577] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[576] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[575] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[574] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[573] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[572] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[571] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[570] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[569] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[568] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[567] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[566] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[565] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[564] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[563] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[562] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[561] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[560] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[559] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[558] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[557] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[556] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[555] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[554] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[553] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[552] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[551] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[550] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[549] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[548] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[547] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[546] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[545] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[544] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[543] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[542] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[541] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[540] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[539] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[538] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[537] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[536] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[535] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[534] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[533] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[532] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[531] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[530] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[529] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[528] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[527] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[526] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[525] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[524] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[523] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[522] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[521] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N86) begin
      ram[520] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[519] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[518] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[517] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[516] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[515] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[514] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[513] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[512] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[511] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[510] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[509] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[508] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[507] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[506] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[505] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[504] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[503] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[502] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[501] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[500] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[499] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[498] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[497] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[496] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[495] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[494] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[493] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[492] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[491] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[490] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[489] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[488] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[487] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[486] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[485] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[484] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[483] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[482] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[481] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[480] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[479] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[478] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[477] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[476] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[475] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[474] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[473] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[472] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[471] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[470] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[469] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[468] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[467] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[466] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[465] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[464] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[463] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[462] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[461] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[460] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[459] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[458] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[457] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[456] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N85) begin
      ram[455] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[454] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[453] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[452] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[451] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[450] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[449] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[448] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[447] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[446] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[445] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[444] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[443] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[442] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[441] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[440] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[439] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[438] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[437] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[436] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[435] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[434] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[433] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[432] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[431] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[430] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[429] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[428] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[427] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[426] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[425] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[424] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[423] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[422] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[421] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[420] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[419] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[418] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[417] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[416] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[415] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[414] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[413] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[412] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[411] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[410] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[409] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[408] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[407] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[406] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[405] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[404] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[403] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[402] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[401] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[400] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[399] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[398] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[397] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[396] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[395] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[394] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[393] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[392] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[391] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N84) begin
      ram[390] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[389] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[388] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[387] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[386] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[385] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[384] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[383] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[382] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[381] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[380] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[379] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[378] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[377] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[376] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[375] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[374] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[373] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[372] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[371] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[370] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[369] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[368] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[367] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[366] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[365] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[364] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[363] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[362] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[361] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[360] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[359] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[358] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[357] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[356] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[355] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[354] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[353] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[352] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[351] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[350] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[349] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[348] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[347] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[346] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[345] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[344] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[343] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[342] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[341] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[340] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[339] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[338] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[337] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[336] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[335] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[334] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[333] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[332] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[331] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[330] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[329] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[328] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[327] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[326] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N83) begin
      ram[325] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[324] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[323] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[322] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[321] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[320] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[319] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[318] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[317] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[316] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[315] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[314] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[313] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[312] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[311] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[310] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[309] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[308] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[307] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[306] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[305] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[304] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[303] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[302] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[301] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[300] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[299] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[298] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[297] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[296] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[295] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[294] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[293] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[292] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[291] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[290] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[289] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[288] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[287] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[286] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[285] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[284] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[283] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[282] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[281] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[280] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[279] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[278] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[277] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[276] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[275] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[274] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[273] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[272] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[271] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[270] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[269] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[268] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[267] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[266] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[265] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[264] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[263] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[262] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[261] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N82) begin
      ram[260] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[259] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[258] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[257] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[256] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[255] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[254] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[253] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[252] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[251] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[250] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[249] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[248] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[247] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[246] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[245] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[244] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[243] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[242] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[241] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[240] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[239] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[238] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[237] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[236] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[235] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[234] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[233] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[232] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[231] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[230] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[229] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[228] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[227] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[226] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[225] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[224] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[223] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[222] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[221] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[220] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[219] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[218] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[217] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[216] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[215] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[214] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[213] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[212] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[211] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[210] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[209] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[208] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[207] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[206] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[205] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[204] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[203] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[202] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[201] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[200] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[199] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[198] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[197] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[196] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N81) begin
      ram[195] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[194] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[193] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[192] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[191] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[190] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[189] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[188] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[187] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[186] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[185] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[184] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[183] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[182] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[181] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[180] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[179] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[178] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[177] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[176] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[175] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[174] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[173] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[172] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[171] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[170] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[169] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[168] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[167] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[166] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[165] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[164] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[163] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[162] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[161] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[160] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[159] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[158] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[157] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[156] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[155] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[154] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[153] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[152] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[151] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[150] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[149] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[148] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[147] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[146] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[145] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[144] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[143] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[142] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[141] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[140] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[139] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[138] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[137] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[136] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[135] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[134] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[133] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[132] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[131] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N80) begin
      ram[130] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[129] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[128] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[127] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[126] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[125] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[124] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[123] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[122] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[121] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[120] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[119] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[118] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[117] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[116] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[115] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[114] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[113] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[112] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[111] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[110] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[109] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[108] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[107] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[106] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[105] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[104] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[103] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[102] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[101] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[100] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[99] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[98] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[97] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[96] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[95] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[94] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[93] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[92] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[91] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[90] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[89] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[88] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[87] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[86] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[85] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[84] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[83] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[82] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[81] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[80] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[79] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[78] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[77] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[76] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[75] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[74] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[73] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[72] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[71] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[70] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[69] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[68] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[67] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[66] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N79) begin
      ram[65] <= io_enq_bits_sdq_id[0];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[64] <= io_enq_bits_addr[39];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[63] <= io_enq_bits_addr[38];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[62] <= io_enq_bits_addr[37];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[61] <= io_enq_bits_addr[36];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[60] <= io_enq_bits_addr[35];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[59] <= io_enq_bits_addr[34];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[58] <= io_enq_bits_addr[33];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[57] <= io_enq_bits_addr[32];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[56] <= io_enq_bits_addr[31];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[55] <= io_enq_bits_addr[30];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[54] <= io_enq_bits_addr[29];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[53] <= io_enq_bits_addr[28];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[52] <= io_enq_bits_addr[27];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[51] <= io_enq_bits_addr[26];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[50] <= io_enq_bits_addr[25];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[49] <= io_enq_bits_addr[24];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[48] <= io_enq_bits_addr[23];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[47] <= io_enq_bits_addr[22];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[46] <= io_enq_bits_addr[21];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[45] <= io_enq_bits_addr[20];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[44] <= io_enq_bits_addr[19];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[43] <= io_enq_bits_addr[18];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[42] <= io_enq_bits_addr[17];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[41] <= io_enq_bits_addr[16];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[40] <= io_enq_bits_addr[15];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[39] <= io_enq_bits_addr[14];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[38] <= io_enq_bits_addr[13];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[37] <= io_enq_bits_addr[12];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[36] <= io_enq_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[35] <= io_enq_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[34] <= io_enq_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[33] <= io_enq_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[32] <= io_enq_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[31] <= io_enq_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[30] <= io_enq_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[29] <= io_enq_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[28] <= io_enq_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[27] <= io_enq_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[26] <= io_enq_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[25] <= io_enq_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[24] <= io_enq_bits_tag[9];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[23] <= io_enq_bits_tag[8];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[22] <= io_enq_bits_tag[7];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[21] <= io_enq_bits_tag[6];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[20] <= io_enq_bits_tag[5];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[19] <= io_enq_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[18] <= io_enq_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[17] <= io_enq_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[16] <= io_enq_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[15] <= io_enq_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[14] <= io_enq_bits_cmd[4];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[13] <= io_enq_bits_cmd[3];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[12] <= io_enq_bits_cmd[2];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[11] <= io_enq_bits_cmd[1];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[10] <= io_enq_bits_cmd[0];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[9] <= io_enq_bits_typ[2];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[8] <= io_enq_bits_typ[1];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[7] <= io_enq_bits_typ[0];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[6] <= io_enq_bits_kill;
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[5] <= io_enq_bits_phys;
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[4] <= io_enq_bits_sdq_id[4];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[3] <= io_enq_bits_sdq_id[3];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[2] <= io_enq_bits_sdq_id[2];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[1] <= io_enq_bits_sdq_id[1];
    end 
  end


  always @(posedge clk) begin
    if(N78) begin
      ram[0] <= io_enq_bits_sdq_id[0];
    end 
  end

  assign io_count[3:0] = R4 - R1;
  assign T3 = R1 + 1'b1;
  assign T6 = R4 + 1'b1;
  assign N98 = R4[2] & R4[3];
  assign N99 = N0 & R4[3];
  assign N0 = ~R4[2];
  assign N100 = R4[2] & N1;
  assign N1 = ~R4[3];
  assign N101 = N2 & N3;
  assign N2 = ~R4[2];
  assign N3 = ~R4[3];
  assign N102 = R4[0] & R4[1];
  assign N103 = N4 & R4[1];
  assign N4 = ~R4[0];
  assign N104 = R4[0] & N5;
  assign N5 = ~R4[1];
  assign N105 = N6 & N7;
  assign N6 = ~R4[0];
  assign N7 = ~R4[1];
  assign N77 = N98 & N102;
  assign N76 = N98 & N103;
  assign N75 = N98 & N104;
  assign N74 = N98 & N105;
  assign N73 = N99 & N102;
  assign N72 = N99 & N103;
  assign N71 = N99 & N104;
  assign N70 = N99 & N105;
  assign N69 = N100 & N102;
  assign N68 = N100 & N103;
  assign N67 = N100 & N104;
  assign N66 = N100 & N105;
  assign N65 = N101 & N102;
  assign N64 = N101 & N103;
  assign N63 = N101 & N104;
  assign N62 = N101 & N105;
  assign N45 = (N8)? 1'b1 : 
               (N95)? 1'b1 : 
               (N44)? 1'b0 : 1'b0;
  assign N8 = reset;
  assign { N49, N48, N47, N46 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N95)? T3 : 1'b0;
  assign N52 = (N8)? 1'b1 : 
               (N96)? 1'b1 : 
               (N51)? 1'b0 : 1'b0;
  assign { N56, N55, N54, N53 } = (N8)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                  (N96)? T6 : 1'b0;
  assign N59 = (N8)? 1'b1 : 
               (N97)? 1'b1 : 
               (N58)? 1'b0 : 1'b0;
  assign N60 = (N8)? 1'b0 : 
               (N97)? do_enq : 1'b0;
  assign { N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78 } = (N9)? { N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62 } : 
                                                                                              (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N9 = do_enq;
  assign N10 = N61;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign io_count[4] = maybe_full & ptr_match;
  assign N11 = ~R1[0];
  assign N12 = ~R1[1];
  assign N13 = N11 & N12;
  assign N14 = N11 & R1[1];
  assign N15 = R1[0] & N12;
  assign N16 = R1[0] & R1[1];
  assign N17 = ~R1[2];
  assign N18 = N13 & N17;
  assign N19 = N13 & R1[2];
  assign N20 = N15 & N17;
  assign N21 = N15 & R1[2];
  assign N22 = N14 & N17;
  assign N23 = N14 & R1[2];
  assign N24 = N16 & N17;
  assign N25 = N16 & R1[2];
  assign N26 = ~R1[3];
  assign N27 = N18 & N26;
  assign N28 = N18 & R1[3];
  assign N29 = N20 & N26;
  assign N30 = N20 & R1[3];
  assign N31 = N22 & N26;
  assign N32 = N22 & R1[3];
  assign N33 = N24 & N26;
  assign N34 = N24 & R1[3];
  assign N35 = N19 & N26;
  assign N36 = N19 & R1[3];
  assign N37 = N21 & N26;
  assign N38 = N21 & R1[3];
  assign N39 = N23 & N26;
  assign N40 = N23 & R1[3];
  assign N41 = N25 & N26;
  assign N42 = N25 & R1[3];
  assign io_deq_valid = ~empty;
  assign empty = ptr_match & T27;
  assign T27 = ~maybe_full;
  assign io_enq_ready = ~full;
  assign full = ptr_match & maybe_full;
  assign N43 = do_deq | reset;
  assign N44 = ~N43;
  assign N50 = do_enq | reset;
  assign N51 = ~N50;
  assign N57 = T9 | reset;
  assign N58 = ~N57;
  assign N61 = ~do_enq;
  assign N94 = ~reset;
  assign N95 = do_deq & N94;
  assign N96 = do_enq & N94;
  assign N97 = T9 & N94;

endmodule