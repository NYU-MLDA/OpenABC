module RoundRawFNToRecFN
(
  io_invalidExc,
  io_infiniteExc,
  io_in_sign,
  io_in_isNaN,
  io_in_isInf,
  io_in_isZero,
  io_in_sExp,
  io_in_sig,
  io_roundingMode,
  io_out,
  io_exceptionFlags
);

  input [9:0] io_in_sExp;
  input [26:0] io_in_sig;
  input [1:0] io_roundingMode;
  output [32:0] io_out;
  output [4:0] io_exceptionFlags;
  input io_invalidExc;
  input io_infiniteExc;
  input io_in_sign;
  input io_in_isNaN;
  input io_in_isInf;
  input io_in_isZero;
  wire [32:0] io_out;
  wire [4:0] io_exceptionFlags;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,io_invalidExc,io_infiniteExc,T3,commonCase,
  anyRound,T60_0,T17_5,T17_3,T17_1,T18_4,T18_2,T21_3,T21_2,T36_13,T36_11,T36_9,T36_7,
  T36_5,T36_3,T36_1,T37_12,T37_10,T37_8,T37_6,T37_4,T37_2,T40_11,T40_10,T40_7,T40_6,
  T40_3,T40_2,T41_9,T41_8,T41_5,T41_4,T44_7,T44_6,T44_5,T44_4,T66,T65,T68,T67,
  notNaN_isSpecialInfOut,common_underflow,T69,common_overflow,T140_9,T88,N10,T82,N11,
  T84,T83,T93,T89,roundMagUp,T92,T90,T91,T99_0,T101,T100,overflow_roundMagUp,T105,
  N12,N13,T106,common_totalUnderflow,notNaN_isInfOut,T110,pegMinNonzeroMagOut,T115,
  T128,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,SV2V_UNCONNECTED_3,
  SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,
  SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,SV2V_UNCONNECTED_10,
  SV2V_UNCONNECTED_11,SV2V_UNCONNECTED_12,SV2V_UNCONNECTED_13,
  SV2V_UNCONNECTED_14,SV2V_UNCONNECTED_15,SV2V_UNCONNECTED_16,SV2V_UNCONNECTED_17,
  SV2V_UNCONNECTED_18,SV2V_UNCONNECTED_19,SV2V_UNCONNECTED_20,
  SV2V_UNCONNECTED_21,SV2V_UNCONNECTED_22,SV2V_UNCONNECTED_23,
  SV2V_UNCONNECTED_24,SV2V_UNCONNECTED_25,SV2V_UNCONNECTED_26,SV2V_UNCONNECTED_27,
  SV2V_UNCONNECTED_28,SV2V_UNCONNECTED_29,SV2V_UNCONNECTED_30,
  SV2V_UNCONNECTED_31,SV2V_UNCONNECTED_32,SV2V_UNCONNECTED_33,
  SV2V_UNCONNECTED_34,SV2V_UNCONNECTED_35,SV2V_UNCONNECTED_36,SV2V_UNCONNECTED_37,
  SV2V_UNCONNECTED_38,SV2V_UNCONNECTED_39,SV2V_UNCONNECTED_40,
  SV2V_UNCONNECTED_41,SV2V_UNCONNECTED_42,SV2V_UNCONNECTED_43,
  SV2V_UNCONNECTED_44,SV2V_UNCONNECTED_45,SV2V_UNCONNECTED_46,SV2V_UNCONNECTED_47,
  SV2V_UNCONNECTED_48,SV2V_UNCONNECTED_49,SV2V_UNCONNECTED_50,
  SV2V_UNCONNECTED_51,SV2V_UNCONNECTED_52,SV2V_UNCONNECTED_53,
  SV2V_UNCONNECTED_54,SV2V_UNCONNECTED_55,SV2V_UNCONNECTED_56,SV2V_UNCONNECTED_57,
  SV2V_UNCONNECTED_58,SV2V_UNCONNECTED_59,SV2V_UNCONNECTED_60,
  SV2V_UNCONNECTED_61,SV2V_UNCONNECTED_62,SV2V_UNCONNECTED_63,
  SV2V_UNCONNECTED_64,SV2V_UNCONNECTED_65,SV2V_UNCONNECTED_66,SV2V_UNCONNECTED_67,
  SV2V_UNCONNECTED_68,SV2V_UNCONNECTED_69,SV2V_UNCONNECTED_70,
  SV2V_UNCONNECTED_71,SV2V_UNCONNECTED_72,SV2V_UNCONNECTED_73,
  SV2V_UNCONNECTED_74,SV2V_UNCONNECTED_75,SV2V_UNCONNECTED_76,SV2V_UNCONNECTED_77,
  SV2V_UNCONNECTED_78,SV2V_UNCONNECTED_79,SV2V_UNCONNECTED_80,
  SV2V_UNCONNECTED_81,SV2V_UNCONNECTED_82,SV2V_UNCONNECTED_83,
  SV2V_UNCONNECTED_84,SV2V_UNCONNECTED_85,SV2V_UNCONNECTED_86,SV2V_UNCONNECTED_87,
  SV2V_UNCONNECTED_88,SV2V_UNCONNECTED_89,SV2V_UNCONNECTED_90,
  SV2V_UNCONNECTED_91,SV2V_UNCONNECTED_92,SV2V_UNCONNECTED_93,
  SV2V_UNCONNECTED_94,SV2V_UNCONNECTED_95,SV2V_UNCONNECTED_96,SV2V_UNCONNECTED_97,
  SV2V_UNCONNECTED_98,SV2V_UNCONNECTED_99,SV2V_UNCONNECTED_100,
  SV2V_UNCONNECTED_101,SV2V_UNCONNECTED_102,SV2V_UNCONNECTED_103,
  SV2V_UNCONNECTED_104,SV2V_UNCONNECTED_105,SV2V_UNCONNECTED_106,
  SV2V_UNCONNECTED_107,SV2V_UNCONNECTED_108,SV2V_UNCONNECTED_109,
  SV2V_UNCONNECTED_110,SV2V_UNCONNECTED_111,SV2V_UNCONNECTED_112,SV2V_UNCONNECTED_113,
  SV2V_UNCONNECTED_114,SV2V_UNCONNECTED_115,SV2V_UNCONNECTED_116,
  SV2V_UNCONNECTED_117,SV2V_UNCONNECTED_118,SV2V_UNCONNECTED_119,
  SV2V_UNCONNECTED_120,SV2V_UNCONNECTED_121,SV2V_UNCONNECTED_122,
  SV2V_UNCONNECTED_123,SV2V_UNCONNECTED_124,SV2V_UNCONNECTED_125,
  SV2V_UNCONNECTED_126,SV2V_UNCONNECTED_127,SV2V_UNCONNECTED_128,SV2V_UNCONNECTED_129,
  SV2V_UNCONNECTED_130,SV2V_UNCONNECTED_131,SV2V_UNCONNECTED_132,
  SV2V_UNCONNECTED_133,SV2V_UNCONNECTED_134,SV2V_UNCONNECTED_135,
  SV2V_UNCONNECTED_136,SV2V_UNCONNECTED_137,SV2V_UNCONNECTED_138,
  SV2V_UNCONNECTED_139,SV2V_UNCONNECTED_140,SV2V_UNCONNECTED_141,
  SV2V_UNCONNECTED_142,SV2V_UNCONNECTED_143,SV2V_UNCONNECTED_144,SV2V_UNCONNECTED_145,
  SV2V_UNCONNECTED_146,SV2V_UNCONNECTED_147,SV2V_UNCONNECTED_148,
  SV2V_UNCONNECTED_149,SV2V_UNCONNECTED_150,SV2V_UNCONNECTED_151,
  SV2V_UNCONNECTED_152,SV2V_UNCONNECTED_153,SV2V_UNCONNECTED_154,
  SV2V_UNCONNECTED_155,SV2V_UNCONNECTED_156,SV2V_UNCONNECTED_157,
  SV2V_UNCONNECTED_158,SV2V_UNCONNECTED_159,SV2V_UNCONNECTED_160,SV2V_UNCONNECTED_161,
  SV2V_UNCONNECTED_162,SV2V_UNCONNECTED_163,SV2V_UNCONNECTED_164,
  SV2V_UNCONNECTED_165,SV2V_UNCONNECTED_166,SV2V_UNCONNECTED_167,
  SV2V_UNCONNECTED_168,SV2V_UNCONNECTED_169,SV2V_UNCONNECTED_170,
  SV2V_UNCONNECTED_171,SV2V_UNCONNECTED_172,SV2V_UNCONNECTED_173,
  SV2V_UNCONNECTED_174,SV2V_UNCONNECTED_175,SV2V_UNCONNECTED_176,SV2V_UNCONNECTED_177,
  SV2V_UNCONNECTED_178,SV2V_UNCONNECTED_179,SV2V_UNCONNECTED_180,
  SV2V_UNCONNECTED_181,SV2V_UNCONNECTED_182,SV2V_UNCONNECTED_183,
  SV2V_UNCONNECTED_184,SV2V_UNCONNECTED_185,SV2V_UNCONNECTED_186,
  SV2V_UNCONNECTED_187,SV2V_UNCONNECTED_188,SV2V_UNCONNECTED_189,
  SV2V_UNCONNECTED_190,SV2V_UNCONNECTED_191,SV2V_UNCONNECTED_192,SV2V_UNCONNECTED_193,
  SV2V_UNCONNECTED_194,SV2V_UNCONNECTED_195,SV2V_UNCONNECTED_196,
  SV2V_UNCONNECTED_197,SV2V_UNCONNECTED_198,SV2V_UNCONNECTED_199,
  SV2V_UNCONNECTED_200,SV2V_UNCONNECTED_201,SV2V_UNCONNECTED_202,
  SV2V_UNCONNECTED_203,SV2V_UNCONNECTED_204,SV2V_UNCONNECTED_205,
  SV2V_UNCONNECTED_206,SV2V_UNCONNECTED_207,SV2V_UNCONNECTED_208,SV2V_UNCONNECTED_209,
  SV2V_UNCONNECTED_210,SV2V_UNCONNECTED_211,SV2V_UNCONNECTED_212,
  SV2V_UNCONNECTED_213,SV2V_UNCONNECTED_214,SV2V_UNCONNECTED_215,
  SV2V_UNCONNECTED_216,SV2V_UNCONNECTED_217,SV2V_UNCONNECTED_218,
  SV2V_UNCONNECTED_219,SV2V_UNCONNECTED_220,SV2V_UNCONNECTED_221,
  SV2V_UNCONNECTED_222,SV2V_UNCONNECTED_223,SV2V_UNCONNECTED_224,SV2V_UNCONNECTED_225,
  SV2V_UNCONNECTED_226,SV2V_UNCONNECTED_227,SV2V_UNCONNECTED_228,
  SV2V_UNCONNECTED_229,SV2V_UNCONNECTED_230,SV2V_UNCONNECTED_231,
  SV2V_UNCONNECTED_232,SV2V_UNCONNECTED_233,SV2V_UNCONNECTED_234,
  SV2V_UNCONNECTED_235,SV2V_UNCONNECTED_236,SV2V_UNCONNECTED_237,
  SV2V_UNCONNECTED_238,SV2V_UNCONNECTED_239,SV2V_UNCONNECTED_240,SV2V_UNCONNECTED_241,
  SV2V_UNCONNECTED_242,SV2V_UNCONNECTED_243,SV2V_UNCONNECTED_244,
  SV2V_UNCONNECTED_245,SV2V_UNCONNECTED_246,SV2V_UNCONNECTED_247,
  SV2V_UNCONNECTED_248,SV2V_UNCONNECTED_249,SV2V_UNCONNECTED_250,
  SV2V_UNCONNECTED_251,SV2V_UNCONNECTED_252,SV2V_UNCONNECTED_253,
  SV2V_UNCONNECTED_254,SV2V_UNCONNECTED_255,SV2V_UNCONNECTED_256,SV2V_UNCONNECTED_257,
  SV2V_UNCONNECTED_258,SV2V_UNCONNECTED_259,SV2V_UNCONNECTED_260,
  SV2V_UNCONNECTED_261,SV2V_UNCONNECTED_262,SV2V_UNCONNECTED_263,
  SV2V_UNCONNECTED_264,SV2V_UNCONNECTED_265,SV2V_UNCONNECTED_266,
  SV2V_UNCONNECTED_267,SV2V_UNCONNECTED_268,SV2V_UNCONNECTED_269,
  SV2V_UNCONNECTED_270,SV2V_UNCONNECTED_271,SV2V_UNCONNECTED_272,SV2V_UNCONNECTED_273,
  SV2V_UNCONNECTED_274,SV2V_UNCONNECTED_275,SV2V_UNCONNECTED_276,
  SV2V_UNCONNECTED_277,SV2V_UNCONNECTED_278,SV2V_UNCONNECTED_279,
  SV2V_UNCONNECTED_280,SV2V_UNCONNECTED_281,SV2V_UNCONNECTED_282,
  SV2V_UNCONNECTED_283,SV2V_UNCONNECTED_284,SV2V_UNCONNECTED_285,
  SV2V_UNCONNECTED_286,SV2V_UNCONNECTED_287,SV2V_UNCONNECTED_288,SV2V_UNCONNECTED_289,
  SV2V_UNCONNECTED_290,SV2V_UNCONNECTED_291,SV2V_UNCONNECTED_292,
  SV2V_UNCONNECTED_293,SV2V_UNCONNECTED_294,SV2V_UNCONNECTED_295,
  SV2V_UNCONNECTED_296,SV2V_UNCONNECTED_297,SV2V_UNCONNECTED_298,
  SV2V_UNCONNECTED_299,SV2V_UNCONNECTED_300,SV2V_UNCONNECTED_301,
  SV2V_UNCONNECTED_302,SV2V_UNCONNECTED_303,SV2V_UNCONNECTED_304,SV2V_UNCONNECTED_305,
  SV2V_UNCONNECTED_306,SV2V_UNCONNECTED_307,SV2V_UNCONNECTED_308,
  SV2V_UNCONNECTED_309,SV2V_UNCONNECTED_310,SV2V_UNCONNECTED_311,
  SV2V_UNCONNECTED_312,SV2V_UNCONNECTED_313,SV2V_UNCONNECTED_314,
  SV2V_UNCONNECTED_315,SV2V_UNCONNECTED_316,SV2V_UNCONNECTED_317,
  SV2V_UNCONNECTED_318,SV2V_UNCONNECTED_319,SV2V_UNCONNECTED_320,SV2V_UNCONNECTED_321,
  SV2V_UNCONNECTED_322,SV2V_UNCONNECTED_323,SV2V_UNCONNECTED_324,
  SV2V_UNCONNECTED_325,SV2V_UNCONNECTED_326,SV2V_UNCONNECTED_327,
  SV2V_UNCONNECTED_328,SV2V_UNCONNECTED_329,SV2V_UNCONNECTED_330,
  SV2V_UNCONNECTED_331,SV2V_UNCONNECTED_332,SV2V_UNCONNECTED_333,
  SV2V_UNCONNECTED_334,SV2V_UNCONNECTED_335,SV2V_UNCONNECTED_336,SV2V_UNCONNECTED_337,
  SV2V_UNCONNECTED_338,SV2V_UNCONNECTED_339,SV2V_UNCONNECTED_340,
  SV2V_UNCONNECTED_341,SV2V_UNCONNECTED_342,SV2V_UNCONNECTED_343,
  SV2V_UNCONNECTED_344,SV2V_UNCONNECTED_345,SV2V_UNCONNECTED_346,
  SV2V_UNCONNECTED_347,SV2V_UNCONNECTED_348,SV2V_UNCONNECTED_349,
  SV2V_UNCONNECTED_350,SV2V_UNCONNECTED_351,SV2V_UNCONNECTED_352,SV2V_UNCONNECTED_353,
  SV2V_UNCONNECTED_354,SV2V_UNCONNECTED_355,SV2V_UNCONNECTED_356,
  SV2V_UNCONNECTED_357,SV2V_UNCONNECTED_358,SV2V_UNCONNECTED_359,
  SV2V_UNCONNECTED_360,SV2V_UNCONNECTED_361,SV2V_UNCONNECTED_362,
  SV2V_UNCONNECTED_363,SV2V_UNCONNECTED_364,SV2V_UNCONNECTED_365,
  SV2V_UNCONNECTED_366,SV2V_UNCONNECTED_367,SV2V_UNCONNECTED_368,SV2V_UNCONNECTED_369,
  SV2V_UNCONNECTED_370,SV2V_UNCONNECTED_371,SV2V_UNCONNECTED_372,
  SV2V_UNCONNECTED_373,SV2V_UNCONNECTED_374,SV2V_UNCONNECTED_375,
  SV2V_UNCONNECTED_376,SV2V_UNCONNECTED_377,SV2V_UNCONNECTED_378,
  SV2V_UNCONNECTED_379,SV2V_UNCONNECTED_380,SV2V_UNCONNECTED_381,
  SV2V_UNCONNECTED_382;
  wire [26:0] T4,T62,roundPosMask;
  wire [25:1] T129;
  wire [24:0] T7,T8,T141,T142,T86;
  wire [24:24] T60;
  wire [7:0] T11;
  wire [15:0] T12;
  wire [8:0] T14,T108,T111,T113,T116,T119,T117,T122,T120,T125,T123,T126;
  wire [7:7] T17,T20,T121;
  wire [6:6] T18,T114,T118;
  wire [7:6] T21,T24;
  wire [5:4] T22;
  wire [15:15] T36,T39;
  wire [14:14] T37;
  wire [15:14] T40,T43;
  wire [13:12] T41;
  wire [15:12] T44,T47;
  wire [11:8] T45;
  wire [0:0] T138,T145;
  wire [25:0] T139,T78,T79,T80;
  wire [1:0] T70,T140;
  wire [2:0] T71;
  wire [6:0] sRoundedExp;
  wire [23:0] roundedSig;
  wire [26:2] T77;
  wire [22:0] T98,T102,common_fractOut;
  wire [22:22] T97,T99;
  wire [8:8] T107,T109,T112,T124,T127;
  assign io_exceptionFlags[4] = io_invalidExc;
  assign io_exceptionFlags[3] = io_infiniteExc;
  assign T138[0] = $signed(io_in_sExp) < $signed(1'b0);
  assign T69 = $signed(io_in_sExp) < $signed({ 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T70 });
  assign common_overflow = $signed({ 1'b0, 1'b1, 1'b1 }) <= $signed(T71);
  assign common_totalUnderflow = $signed({ T71, sRoundedExp }) < $signed({ 1'b0, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 });
  assign N15 = ~io_roundingMode[1];
  assign N16 = io_roundingMode[0] | N15;
  assign N17 = ~N16;
  assign N18 = io_roundingMode[0] & io_roundingMode[1];
  assign N19 = io_roundingMode[0] | io_roundingMode[1];
  assign N20 = ~N19;
  assign N21 = T62[25] | T62[26];
  assign N22 = T62[24] | N21;
  assign N23 = T62[23] | N22;
  assign N24 = T62[22] | N23;
  assign N25 = T62[21] | N24;
  assign N26 = T62[20] | N25;
  assign N27 = T62[19] | N26;
  assign N28 = T62[18] | N27;
  assign N29 = T62[17] | N28;
  assign N30 = T62[16] | N29;
  assign N31 = T62[15] | N30;
  assign N32 = T62[14] | N31;
  assign N33 = T62[13] | N32;
  assign N34 = T62[12] | N33;
  assign N35 = T62[11] | N34;
  assign N36 = T62[10] | N35;
  assign N37 = T62[9] | N36;
  assign N38 = T62[8] | N37;
  assign N39 = T62[7] | N38;
  assign N40 = T62[6] | N39;
  assign N41 = T62[5] | N40;
  assign N42 = T62[4] | N41;
  assign N43 = T62[3] | N42;
  assign N44 = T62[2] | N43;
  assign N45 = T62[1] | N44;
  assign N46 = T62[0] | N45;
  assign N47 = T4[25] | T4[26];
  assign N48 = T4[24] | N47;
  assign N49 = T4[23] | N48;
  assign N50 = T4[22] | N49;
  assign N51 = T4[21] | N50;
  assign N52 = T4[20] | N51;
  assign N53 = T4[19] | N52;
  assign N54 = T4[18] | N53;
  assign N55 = T4[17] | N54;
  assign N56 = T4[16] | N55;
  assign N57 = T4[15] | N56;
  assign N58 = T4[14] | N57;
  assign N59 = T4[13] | N58;
  assign N60 = T4[12] | N59;
  assign N61 = T4[11] | N60;
  assign N62 = T4[10] | N61;
  assign N63 = T4[9] | N62;
  assign N64 = T4[8] | N63;
  assign N65 = T4[7] | N64;
  assign N66 = T4[6] | N65;
  assign N67 = T4[5] | N66;
  assign N68 = T4[4] | N67;
  assign N69 = T4[3] | N68;
  assign N70 = T4[2] | N69;
  assign N71 = T4[1] | N70;
  assign N72 = T4[0] | N71;
  assign { SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, SV2V_UNCONNECTED_16, SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, SV2V_UNCONNECTED_32, SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, SV2V_UNCONNECTED_49, SV2V_UNCONNECTED_50, SV2V_UNCONNECTED_51, SV2V_UNCONNECTED_52, SV2V_UNCONNECTED_53, SV2V_UNCONNECTED_54, SV2V_UNCONNECTED_55, SV2V_UNCONNECTED_56, SV2V_UNCONNECTED_57, SV2V_UNCONNECTED_58, SV2V_UNCONNECTED_59, SV2V_UNCONNECTED_60, SV2V_UNCONNECTED_61, SV2V_UNCONNECTED_62, SV2V_UNCONNECTED_63, SV2V_UNCONNECTED_64, SV2V_UNCONNECTED_65, SV2V_UNCONNECTED_66, SV2V_UNCONNECTED_67, SV2V_UNCONNECTED_68, SV2V_UNCONNECTED_69, SV2V_UNCONNECTED_70, SV2V_UNCONNECTED_71, SV2V_UNCONNECTED_72, SV2V_UNCONNECTED_73, SV2V_UNCONNECTED_74, SV2V_UNCONNECTED_75, SV2V_UNCONNECTED_76, SV2V_UNCONNECTED_77, SV2V_UNCONNECTED_78, SV2V_UNCONNECTED_79, SV2V_UNCONNECTED_80, SV2V_UNCONNECTED_81, SV2V_UNCONNECTED_82, SV2V_UNCONNECTED_83, SV2V_UNCONNECTED_84, SV2V_UNCONNECTED_85, SV2V_UNCONNECTED_86, SV2V_UNCONNECTED_87, SV2V_UNCONNECTED_88, SV2V_UNCONNECTED_89, SV2V_UNCONNECTED_90, SV2V_UNCONNECTED_91, SV2V_UNCONNECTED_92, SV2V_UNCONNECTED_93, SV2V_UNCONNECTED_94, SV2V_UNCONNECTED_95, SV2V_UNCONNECTED_96, SV2V_UNCONNECTED_97, SV2V_UNCONNECTED_98, SV2V_UNCONNECTED_99, SV2V_UNCONNECTED_100, SV2V_UNCONNECTED_101, SV2V_UNCONNECTED_102, SV2V_UNCONNECTED_103, SV2V_UNCONNECTED_104, SV2V_UNCONNECTED_105, SV2V_UNCONNECTED_106, SV2V_UNCONNECTED_107, SV2V_UNCONNECTED_108, SV2V_UNCONNECTED_109, SV2V_UNCONNECTED_110, SV2V_UNCONNECTED_111, SV2V_UNCONNECTED_112, SV2V_UNCONNECTED_113, SV2V_UNCONNECTED_114, SV2V_UNCONNECTED_115, SV2V_UNCONNECTED_116, SV2V_UNCONNECTED_117, SV2V_UNCONNECTED_118, SV2V_UNCONNECTED_119, SV2V_UNCONNECTED_120, SV2V_UNCONNECTED_121, SV2V_UNCONNECTED_122, SV2V_UNCONNECTED_123, SV2V_UNCONNECTED_124, SV2V_UNCONNECTED_125, SV2V_UNCONNECTED_126, SV2V_UNCONNECTED_127, SV2V_UNCONNECTED_128, SV2V_UNCONNECTED_129, SV2V_UNCONNECTED_130, SV2V_UNCONNECTED_131, SV2V_UNCONNECTED_132, SV2V_UNCONNECTED_133, SV2V_UNCONNECTED_134, SV2V_UNCONNECTED_135, SV2V_UNCONNECTED_136, SV2V_UNCONNECTED_137, SV2V_UNCONNECTED_138, SV2V_UNCONNECTED_139, SV2V_UNCONNECTED_140, SV2V_UNCONNECTED_141, SV2V_UNCONNECTED_142, SV2V_UNCONNECTED_143, SV2V_UNCONNECTED_144, SV2V_UNCONNECTED_145, SV2V_UNCONNECTED_146, SV2V_UNCONNECTED_147, SV2V_UNCONNECTED_148, SV2V_UNCONNECTED_149, SV2V_UNCONNECTED_150, SV2V_UNCONNECTED_151, SV2V_UNCONNECTED_152, SV2V_UNCONNECTED_153, SV2V_UNCONNECTED_154, SV2V_UNCONNECTED_155, SV2V_UNCONNECTED_156, SV2V_UNCONNECTED_157, SV2V_UNCONNECTED_158, SV2V_UNCONNECTED_159, SV2V_UNCONNECTED_160, SV2V_UNCONNECTED_161, SV2V_UNCONNECTED_162, SV2V_UNCONNECTED_163, SV2V_UNCONNECTED_164, SV2V_UNCONNECTED_165, SV2V_UNCONNECTED_166, SV2V_UNCONNECTED_167, SV2V_UNCONNECTED_168, SV2V_UNCONNECTED_169, SV2V_UNCONNECTED_170, SV2V_UNCONNECTED_171, SV2V_UNCONNECTED_172, SV2V_UNCONNECTED_173, SV2V_UNCONNECTED_174, SV2V_UNCONNECTED_175, SV2V_UNCONNECTED_176, SV2V_UNCONNECTED_177, SV2V_UNCONNECTED_178, SV2V_UNCONNECTED_179, SV2V_UNCONNECTED_180, SV2V_UNCONNECTED_181, SV2V_UNCONNECTED_182, SV2V_UNCONNECTED_183, SV2V_UNCONNECTED_184, SV2V_UNCONNECTED_185, SV2V_UNCONNECTED_186, SV2V_UNCONNECTED_187, SV2V_UNCONNECTED_188, SV2V_UNCONNECTED_189, SV2V_UNCONNECTED_190, SV2V_UNCONNECTED_191, SV2V_UNCONNECTED_192, SV2V_UNCONNECTED_193, SV2V_UNCONNECTED_194, SV2V_UNCONNECTED_195, SV2V_UNCONNECTED_196, SV2V_UNCONNECTED_197, SV2V_UNCONNECTED_198, SV2V_UNCONNECTED_199, SV2V_UNCONNECTED_200, SV2V_UNCONNECTED_201, SV2V_UNCONNECTED_202, SV2V_UNCONNECTED_203, SV2V_UNCONNECTED_204, SV2V_UNCONNECTED_205, SV2V_UNCONNECTED_206, SV2V_UNCONNECTED_207, SV2V_UNCONNECTED_208, SV2V_UNCONNECTED_209, SV2V_UNCONNECTED_210, SV2V_UNCONNECTED_211, SV2V_UNCONNECTED_212, SV2V_UNCONNECTED_213, SV2V_UNCONNECTED_214, SV2V_UNCONNECTED_215, SV2V_UNCONNECTED_216, SV2V_UNCONNECTED_217, SV2V_UNCONNECTED_218, SV2V_UNCONNECTED_219, SV2V_UNCONNECTED_220, SV2V_UNCONNECTED_221, SV2V_UNCONNECTED_222, SV2V_UNCONNECTED_223, SV2V_UNCONNECTED_224, SV2V_UNCONNECTED_225, SV2V_UNCONNECTED_226, SV2V_UNCONNECTED_227, SV2V_UNCONNECTED_228, SV2V_UNCONNECTED_229, SV2V_UNCONNECTED_230, SV2V_UNCONNECTED_231, SV2V_UNCONNECTED_232, SV2V_UNCONNECTED_233, SV2V_UNCONNECTED_234, SV2V_UNCONNECTED_235, SV2V_UNCONNECTED_236, SV2V_UNCONNECTED_237, SV2V_UNCONNECTED_238, SV2V_UNCONNECTED_239, SV2V_UNCONNECTED_240, SV2V_UNCONNECTED_241, SV2V_UNCONNECTED_242, SV2V_UNCONNECTED_243, SV2V_UNCONNECTED_244, SV2V_UNCONNECTED_245, SV2V_UNCONNECTED_246, SV2V_UNCONNECTED_247, SV2V_UNCONNECTED_248, SV2V_UNCONNECTED_249, SV2V_UNCONNECTED_250, SV2V_UNCONNECTED_251, SV2V_UNCONNECTED_252, SV2V_UNCONNECTED_253, SV2V_UNCONNECTED_254, SV2V_UNCONNECTED_255, SV2V_UNCONNECTED_256, SV2V_UNCONNECTED_257, SV2V_UNCONNECTED_258, SV2V_UNCONNECTED_259, SV2V_UNCONNECTED_260, SV2V_UNCONNECTED_261, SV2V_UNCONNECTED_262, SV2V_UNCONNECTED_263, SV2V_UNCONNECTED_264, SV2V_UNCONNECTED_265, SV2V_UNCONNECTED_266, SV2V_UNCONNECTED_267, SV2V_UNCONNECTED_268, SV2V_UNCONNECTED_269, SV2V_UNCONNECTED_270, SV2V_UNCONNECTED_271, SV2V_UNCONNECTED_272, SV2V_UNCONNECTED_273, SV2V_UNCONNECTED_274, SV2V_UNCONNECTED_275, SV2V_UNCONNECTED_276, SV2V_UNCONNECTED_277, SV2V_UNCONNECTED_278, SV2V_UNCONNECTED_279, SV2V_UNCONNECTED_280, SV2V_UNCONNECTED_281, SV2V_UNCONNECTED_282, SV2V_UNCONNECTED_283, SV2V_UNCONNECTED_284, SV2V_UNCONNECTED_285, SV2V_UNCONNECTED_286, SV2V_UNCONNECTED_287, SV2V_UNCONNECTED_288, SV2V_UNCONNECTED_289, SV2V_UNCONNECTED_290, SV2V_UNCONNECTED_291, SV2V_UNCONNECTED_292, SV2V_UNCONNECTED_293, SV2V_UNCONNECTED_294, SV2V_UNCONNECTED_295, SV2V_UNCONNECTED_296, SV2V_UNCONNECTED_297, SV2V_UNCONNECTED_298, SV2V_UNCONNECTED_299, SV2V_UNCONNECTED_300, SV2V_UNCONNECTED_301, SV2V_UNCONNECTED_302, SV2V_UNCONNECTED_303, SV2V_UNCONNECTED_304, SV2V_UNCONNECTED_305, SV2V_UNCONNECTED_306, SV2V_UNCONNECTED_307, SV2V_UNCONNECTED_308, SV2V_UNCONNECTED_309, SV2V_UNCONNECTED_310, SV2V_UNCONNECTED_311, SV2V_UNCONNECTED_312, SV2V_UNCONNECTED_313, SV2V_UNCONNECTED_314, SV2V_UNCONNECTED_315, SV2V_UNCONNECTED_316, SV2V_UNCONNECTED_317, SV2V_UNCONNECTED_318, SV2V_UNCONNECTED_319, SV2V_UNCONNECTED_320, SV2V_UNCONNECTED_321, SV2V_UNCONNECTED_322, SV2V_UNCONNECTED_323, SV2V_UNCONNECTED_324, SV2V_UNCONNECTED_325, SV2V_UNCONNECTED_326, SV2V_UNCONNECTED_327, SV2V_UNCONNECTED_328, SV2V_UNCONNECTED_329, SV2V_UNCONNECTED_330, SV2V_UNCONNECTED_331, SV2V_UNCONNECTED_332, SV2V_UNCONNECTED_333, SV2V_UNCONNECTED_334, SV2V_UNCONNECTED_335, SV2V_UNCONNECTED_336, SV2V_UNCONNECTED_337, SV2V_UNCONNECTED_338, SV2V_UNCONNECTED_339, SV2V_UNCONNECTED_340, SV2V_UNCONNECTED_341, SV2V_UNCONNECTED_342, SV2V_UNCONNECTED_343, SV2V_UNCONNECTED_344, SV2V_UNCONNECTED_345, SV2V_UNCONNECTED_346, SV2V_UNCONNECTED_347, SV2V_UNCONNECTED_348, SV2V_UNCONNECTED_349, SV2V_UNCONNECTED_350, SV2V_UNCONNECTED_351, SV2V_UNCONNECTED_352, SV2V_UNCONNECTED_353, SV2V_UNCONNECTED_354, SV2V_UNCONNECTED_355, SV2V_UNCONNECTED_356, SV2V_UNCONNECTED_357, SV2V_UNCONNECTED_358, SV2V_UNCONNECTED_359, SV2V_UNCONNECTED_360, SV2V_UNCONNECTED_361, SV2V_UNCONNECTED_362, SV2V_UNCONNECTED_363, SV2V_UNCONNECTED_364, SV2V_UNCONNECTED_365, SV2V_UNCONNECTED_366, SV2V_UNCONNECTED_367, SV2V_UNCONNECTED_368, SV2V_UNCONNECTED_369, SV2V_UNCONNECTED_370, SV2V_UNCONNECTED_371, SV2V_UNCONNECTED_372, SV2V_UNCONNECTED_373, SV2V_UNCONNECTED_374, SV2V_UNCONNECTED_375, SV2V_UNCONNECTED_376, SV2V_UNCONNECTED_377, SV2V_UNCONNECTED_378, SV2V_UNCONNECTED_379, SV2V_UNCONNECTED_380, SV2V_UNCONNECTED_381, SV2V_UNCONNECTED_382, T8[0:0], T11, T12 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> T14;
  assign { T60[24:24], T60_0 } = 1'b0 - T138[0];
  assign T142 = T86 + 1'b1;
  assign { T71, sRoundedExp } = io_in_sExp + { T140_9, T140_9, T140_9, T140_9, T140_9, T140_9, T140_9, 1'b0, T140 };
  assign { T99[22:22], T99_0 } = 1'b0 - T145[0];
  assign { T140, roundedSig } = (N0)? T78 : 
                                (N1)? { 1'b0, T141 } : 1'b0;
  assign N0 = T88;
  assign N1 = N10;
  assign T80[25:1] = (N2)? T129 : 
                     (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = T80[0];
  assign N3 = N11;
  assign T102 = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N5)? common_fractOut : 1'b0;
  assign N4 = T105;
  assign N5 = N12;
  assign common_fractOut = (N6)? roundedSig[23:1] : 
                           (N7)? roundedSig[22:0] : 1'b0;
  assign N6 = T70[0];
  assign N7 = T70[1];
  assign io_out[32] = (N8)? 1'b0 : 
                      (N9)? io_in_sign : 1'b0;
  assign N8 = T97[22];
  assign N9 = N14;
  assign io_exceptionFlags[0] = io_exceptionFlags[2] | T3;
  assign T3 = commonCase & anyRound;
  assign anyRound = N46 | N72;
  assign T4[26] = io_in_sig[26] & 1'b0;
  assign T4[25] = io_in_sig[25] & T129[25];
  assign T4[24] = io_in_sig[24] & T129[24];
  assign T4[23] = io_in_sig[23] & T129[23];
  assign T4[22] = io_in_sig[22] & T129[22];
  assign T4[21] = io_in_sig[21] & T129[21];
  assign T4[20] = io_in_sig[20] & T129[20];
  assign T4[19] = io_in_sig[19] & T129[19];
  assign T4[18] = io_in_sig[18] & T129[18];
  assign T4[17] = io_in_sig[17] & T129[17];
  assign T4[16] = io_in_sig[16] & T129[16];
  assign T4[15] = io_in_sig[15] & T129[15];
  assign T4[14] = io_in_sig[14] & T129[14];
  assign T4[13] = io_in_sig[13] & T129[13];
  assign T4[12] = io_in_sig[12] & T129[12];
  assign T4[11] = io_in_sig[11] & T129[11];
  assign T4[10] = io_in_sig[10] & T129[10];
  assign T4[9] = io_in_sig[9] & T129[9];
  assign T4[8] = io_in_sig[8] & T129[8];
  assign T4[7] = io_in_sig[7] & T129[7];
  assign T4[6] = io_in_sig[6] & T129[6];
  assign T4[5] = io_in_sig[5] & T129[5];
  assign T4[4] = io_in_sig[4] & T129[4];
  assign T4[3] = io_in_sig[3] & T129[3];
  assign T4[2] = io_in_sig[2] & T129[2];
  assign T4[1] = io_in_sig[1] & T129[1];
  assign T4[0] = io_in_sig[0] & 1'b1;
  assign T129[25] = T7[24] | 1'b0;
  assign T129[24] = T7[23] | 1'b0;
  assign T129[23] = T7[22] | 1'b0;
  assign T129[22] = T7[21] | 1'b0;
  assign T129[21] = T7[20] | 1'b0;
  assign T129[20] = T7[19] | 1'b0;
  assign T129[19] = T7[18] | 1'b0;
  assign T129[18] = T7[17] | 1'b0;
  assign T129[17] = T7[16] | 1'b0;
  assign T129[16] = T7[15] | 1'b0;
  assign T129[15] = T7[14] | 1'b0;
  assign T129[14] = T7[13] | 1'b0;
  assign T129[13] = T7[12] | 1'b0;
  assign T129[12] = T7[11] | 1'b0;
  assign T129[11] = T7[10] | 1'b0;
  assign T129[10] = T7[9] | 1'b0;
  assign T129[9] = T7[8] | 1'b0;
  assign T129[8] = T7[7] | 1'b0;
  assign T129[7] = T7[6] | 1'b0;
  assign T129[6] = T7[5] | 1'b0;
  assign T129[5] = T7[4] | 1'b0;
  assign T129[4] = T7[3] | 1'b0;
  assign T129[3] = T7[2] | 1'b0;
  assign T129[2] = T7[1] | 1'b0;
  assign T129[1] = T7[0] | io_in_sig[26];
  assign T7[24] = T60[24] | T8[24];
  assign T7[23] = T60[24] | T8[23];
  assign T7[22] = T60[24] | T8[22];
  assign T7[21] = T60[24] | T8[21];
  assign T7[20] = T60[24] | T8[20];
  assign T7[19] = T60[24] | T8[19];
  assign T7[18] = T60[24] | T8[18];
  assign T7[17] = T60[24] | T8[17];
  assign T7[16] = T60[24] | T8[16];
  assign T7[15] = T60[24] | T8[15];
  assign T7[14] = T60[24] | T8[14];
  assign T7[13] = T60[24] | T8[13];
  assign T7[12] = T60[24] | T8[12];
  assign T7[11] = T60[24] | T8[11];
  assign T7[10] = T60[24] | T8[10];
  assign T7[9] = T60[24] | T8[9];
  assign T7[8] = T60[24] | T8[8];
  assign T7[7] = T60[24] | T8[7];
  assign T7[6] = T60[24] | T8[6];
  assign T7[5] = T60[24] | T8[5];
  assign T7[4] = T60[24] | T8[4];
  assign T7[3] = T60[24] | T8[3];
  assign T7[2] = T60[24] | T8[2];
  assign T7[1] = T60[24] | T8[1];
  assign T7[0] = T60_0 | T8[0];
  assign T14[8] = ~io_in_sExp[8];
  assign T14[7] = ~io_in_sExp[7];
  assign T14[6] = ~io_in_sExp[6];
  assign T14[5] = ~io_in_sExp[5];
  assign T14[4] = ~io_in_sExp[4];
  assign T14[3] = ~io_in_sExp[3];
  assign T14[2] = ~io_in_sExp[2];
  assign T14[1] = ~io_in_sExp[1];
  assign T14[0] = ~io_in_sExp[0];
  assign T8[8] = 1'b0 | T17[7];
  assign T8[7] = T20[7] | 1'b0;
  assign T8[6] = 1'b0 | T17_5;
  assign T8[5] = T18[6] | 1'b0;
  assign T8[4] = 1'b0 | T17_3;
  assign T8[3] = T18_4 | 1'b0;
  assign T8[2] = 1'b0 | T17_1;
  assign T8[1] = T18_2 | 1'b0;
  assign T20[7] = 1'b0 | T21[7];
  assign T17[7] = 1'b0 | T21[6];
  assign T18[6] = T24[7] | 1'b0;
  assign T17_5 = T24[6] | 1'b0;
  assign T18_4 = 1'b0 | T21_3;
  assign T17_3 = 1'b0 | T21_2;
  assign T18_2 = T22[5] | 1'b0;
  assign T17_1 = T22[4] | 1'b0;
  assign T24[7] = 1'b0 | T11[3];
  assign T24[6] = 1'b0 | T11[2];
  assign T21[7] = 1'b0 | T11[1];
  assign T21[6] = 1'b0 | T11[0];
  assign T22[5] = T11[7] | 1'b0;
  assign T22[4] = T11[6] | 1'b0;
  assign T21_3 = T11[5] | 1'b0;
  assign T21_2 = T11[4] | 1'b0;
  assign T8[24] = 1'b0 | T36[15];
  assign T8[23] = T39[15] | 1'b0;
  assign T8[22] = 1'b0 | T36_13;
  assign T8[21] = T37[14] | 1'b0;
  assign T8[20] = 1'b0 | T36_11;
  assign T8[19] = T37_12 | 1'b0;
  assign T8[18] = 1'b0 | T36_9;
  assign T8[17] = T37_10 | 1'b0;
  assign T8[16] = 1'b0 | T36_7;
  assign T8[15] = T37_8 | 1'b0;
  assign T8[14] = 1'b0 | T36_5;
  assign T8[13] = T37_6 | 1'b0;
  assign T8[12] = 1'b0 | T36_3;
  assign T8[11] = T37_4 | 1'b0;
  assign T8[10] = 1'b0 | T36_1;
  assign T8[9] = T37_2 | 1'b0;
  assign T39[15] = 1'b0 | T40[15];
  assign T36[15] = 1'b0 | T40[14];
  assign T37[14] = T43[15] | 1'b0;
  assign T36_13 = T43[14] | 1'b0;
  assign T37_12 = 1'b0 | T40_11;
  assign T36_11 = 1'b0 | T40_10;
  assign T37_10 = T41[13] | 1'b0;
  assign T36_9 = T41[12] | 1'b0;
  assign T37_8 = 1'b0 | T40_7;
  assign T36_7 = 1'b0 | T40_6;
  assign T37_6 = T41_9 | 1'b0;
  assign T36_5 = T41_8 | 1'b0;
  assign T37_4 = 1'b0 | T40_3;
  assign T36_3 = 1'b0 | T40_2;
  assign T37_2 = T41_5 | 1'b0;
  assign T36_1 = T41_4 | 1'b0;
  assign T43[15] = 1'b0 | T44[15];
  assign T43[14] = 1'b0 | T44[14];
  assign T40[15] = 1'b0 | T44[13];
  assign T40[14] = 1'b0 | T44[12];
  assign T41[13] = T47[15] | 1'b0;
  assign T41[12] = T47[14] | 1'b0;
  assign T40_11 = T47[13] | 1'b0;
  assign T40_10 = T47[12] | 1'b0;
  assign T41_9 = 1'b0 | T44_7;
  assign T41_8 = 1'b0 | T44_6;
  assign T40_7 = 1'b0 | T44_5;
  assign T40_6 = 1'b0 | T44_4;
  assign T41_5 = T45[11] | 1'b0;
  assign T41_4 = T45[10] | 1'b0;
  assign T40_3 = T45[9] | 1'b0;
  assign T40_2 = T45[8] | 1'b0;
  assign T47[15] = 1'b0 | T12[7];
  assign T47[14] = 1'b0 | T12[6];
  assign T47[13] = 1'b0 | T12[5];
  assign T47[12] = 1'b0 | T12[4];
  assign T44[15] = 1'b0 | T12[3];
  assign T44[14] = 1'b0 | T12[2];
  assign T44[13] = 1'b0 | T12[1];
  assign T44[12] = 1'b0 | T12[0];
  assign T45[11] = T12[15] | 1'b0;
  assign T45[10] = T12[14] | 1'b0;
  assign T45[9] = T12[13] | 1'b0;
  assign T45[8] = T12[12] | 1'b0;
  assign T44_7 = T12[11] | 1'b0;
  assign T44_6 = T12[10] | 1'b0;
  assign T44_5 = T12[9] | 1'b0;
  assign T44_4 = T12[8] | 1'b0;
  assign T62[26] = io_in_sig[26] & roundPosMask[26];
  assign T62[25] = io_in_sig[25] & roundPosMask[25];
  assign T62[24] = io_in_sig[24] & roundPosMask[24];
  assign T62[23] = io_in_sig[23] & roundPosMask[23];
  assign T62[22] = io_in_sig[22] & roundPosMask[22];
  assign T62[21] = io_in_sig[21] & roundPosMask[21];
  assign T62[20] = io_in_sig[20] & roundPosMask[20];
  assign T62[19] = io_in_sig[19] & roundPosMask[19];
  assign T62[18] = io_in_sig[18] & roundPosMask[18];
  assign T62[17] = io_in_sig[17] & roundPosMask[17];
  assign T62[16] = io_in_sig[16] & roundPosMask[16];
  assign T62[15] = io_in_sig[15] & roundPosMask[15];
  assign T62[14] = io_in_sig[14] & roundPosMask[14];
  assign T62[13] = io_in_sig[13] & roundPosMask[13];
  assign T62[12] = io_in_sig[12] & roundPosMask[12];
  assign T62[11] = io_in_sig[11] & roundPosMask[11];
  assign T62[10] = io_in_sig[10] & roundPosMask[10];
  assign T62[9] = io_in_sig[9] & roundPosMask[9];
  assign T62[8] = io_in_sig[8] & roundPosMask[8];
  assign T62[7] = io_in_sig[7] & roundPosMask[7];
  assign T62[6] = io_in_sig[6] & roundPosMask[6];
  assign T62[5] = io_in_sig[5] & roundPosMask[5];
  assign T62[4] = io_in_sig[4] & roundPosMask[4];
  assign T62[3] = io_in_sig[3] & roundPosMask[3];
  assign T62[2] = io_in_sig[2] & roundPosMask[2];
  assign T62[1] = io_in_sig[1] & roundPosMask[1];
  assign T62[0] = io_in_sig[0] & roundPosMask[0];
  assign roundPosMask[26] = 1'b0 & T129[25];
  assign roundPosMask[25] = T139[25] & T129[24];
  assign roundPosMask[24] = T139[24] & T129[23];
  assign roundPosMask[23] = T139[23] & T129[22];
  assign roundPosMask[22] = T139[22] & T129[21];
  assign roundPosMask[21] = T139[21] & T129[20];
  assign roundPosMask[20] = T139[20] & T129[19];
  assign roundPosMask[19] = T139[19] & T129[18];
  assign roundPosMask[18] = T139[18] & T129[17];
  assign roundPosMask[17] = T139[17] & T129[16];
  assign roundPosMask[16] = T139[16] & T129[15];
  assign roundPosMask[15] = T139[15] & T129[14];
  assign roundPosMask[14] = T139[14] & T129[13];
  assign roundPosMask[13] = T139[13] & T129[12];
  assign roundPosMask[12] = T139[12] & T129[11];
  assign roundPosMask[11] = T139[11] & T129[10];
  assign roundPosMask[10] = T139[10] & T129[9];
  assign roundPosMask[9] = T139[9] & T129[8];
  assign roundPosMask[8] = T139[8] & T129[7];
  assign roundPosMask[7] = T139[7] & T129[6];
  assign roundPosMask[6] = T139[6] & T129[5];
  assign roundPosMask[5] = T139[5] & T129[4];
  assign roundPosMask[4] = T139[4] & T129[3];
  assign roundPosMask[3] = T139[3] & T129[2];
  assign roundPosMask[2] = T139[2] & T129[1];
  assign roundPosMask[1] = T139[1] & 1'b1;
  assign roundPosMask[0] = T139[0] & 1'b1;
  assign T139[25] = ~T129[25];
  assign T139[24] = ~T129[24];
  assign T139[23] = ~T129[23];
  assign T139[22] = ~T129[22];
  assign T139[21] = ~T129[21];
  assign T139[20] = ~T129[20];
  assign T139[19] = ~T129[19];
  assign T139[18] = ~T129[18];
  assign T139[17] = ~T129[17];
  assign T139[16] = ~T129[16];
  assign T139[15] = ~T129[15];
  assign T139[14] = ~T129[14];
  assign T139[13] = ~T129[13];
  assign T139[12] = ~T129[12];
  assign T139[11] = ~T129[11];
  assign T139[10] = ~T129[10];
  assign T139[9] = ~T129[9];
  assign T139[8] = ~T129[8];
  assign T139[7] = ~T129[7];
  assign T139[6] = ~T129[6];
  assign T139[5] = ~T129[5];
  assign T139[4] = ~T129[4];
  assign T139[3] = ~T129[3];
  assign T139[2] = ~T129[2];
  assign T139[1] = ~T129[1];
  assign T139[0] = ~1'b1;
  assign commonCase = T66 & T65;
  assign T65 = ~io_in_isZero;
  assign T66 = T68 & T67;
  assign T67 = ~notNaN_isSpecialInfOut;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T68 = ~T97[22];
  assign T97[22] = io_invalidExc | io_in_isNaN;
  assign io_exceptionFlags[1] = commonCase & common_underflow;
  assign common_underflow = anyRound & T69;
  assign io_exceptionFlags[2] = commonCase & common_overflow;
  assign N10 = ~T88;
  assign T141[24] = io_in_sig[26] & T77[26];
  assign T141[23] = io_in_sig[25] & T77[25];
  assign T141[22] = io_in_sig[24] & T77[24];
  assign T141[21] = io_in_sig[23] & T77[23];
  assign T141[20] = io_in_sig[22] & T77[22];
  assign T141[19] = io_in_sig[21] & T77[21];
  assign T141[18] = io_in_sig[20] & T77[20];
  assign T141[17] = io_in_sig[19] & T77[19];
  assign T141[16] = io_in_sig[18] & T77[18];
  assign T141[15] = io_in_sig[17] & T77[17];
  assign T141[14] = io_in_sig[16] & T77[16];
  assign T141[13] = io_in_sig[15] & T77[15];
  assign T141[12] = io_in_sig[14] & T77[14];
  assign T141[11] = io_in_sig[13] & T77[13];
  assign T141[10] = io_in_sig[12] & T77[12];
  assign T141[9] = io_in_sig[11] & T77[11];
  assign T141[8] = io_in_sig[10] & T77[10];
  assign T141[7] = io_in_sig[9] & T77[9];
  assign T141[6] = io_in_sig[8] & T77[8];
  assign T141[5] = io_in_sig[7] & T77[7];
  assign T141[4] = io_in_sig[6] & T77[6];
  assign T141[3] = io_in_sig[5] & T77[5];
  assign T141[2] = io_in_sig[4] & T77[4];
  assign T141[1] = io_in_sig[3] & T77[3];
  assign T141[0] = io_in_sig[2] & T77[2];
  assign T77[26] = ~T129[25];
  assign T77[25] = ~T129[24];
  assign T77[24] = ~T129[23];
  assign T77[23] = ~T129[22];
  assign T77[22] = ~T129[21];
  assign T77[21] = ~T129[20];
  assign T77[20] = ~T129[19];
  assign T77[19] = ~T129[18];
  assign T77[18] = ~T129[17];
  assign T77[17] = ~T129[16];
  assign T77[16] = ~T129[15];
  assign T77[15] = ~T129[14];
  assign T77[14] = ~T129[13];
  assign T77[13] = ~T129[12];
  assign T77[12] = ~T129[11];
  assign T77[11] = ~T129[10];
  assign T77[10] = ~T129[9];
  assign T77[9] = ~T129[8];
  assign T77[8] = ~T129[7];
  assign T77[7] = ~T129[6];
  assign T77[6] = ~T129[5];
  assign T77[5] = ~T129[4];
  assign T77[4] = ~T129[3];
  assign T77[3] = ~T129[2];
  assign T77[2] = ~T129[1];
  assign T78[25] = 1'b0 & T79[25];
  assign T78[24] = T142[24] & T79[24];
  assign T78[23] = T142[23] & T79[23];
  assign T78[22] = T142[22] & T79[22];
  assign T78[21] = T142[21] & T79[21];
  assign T78[20] = T142[20] & T79[20];
  assign T78[19] = T142[19] & T79[19];
  assign T78[18] = T142[18] & T79[18];
  assign T78[17] = T142[17] & T79[17];
  assign T78[16] = T142[16] & T79[16];
  assign T78[15] = T142[15] & T79[15];
  assign T78[14] = T142[14] & T79[14];
  assign T78[13] = T142[13] & T79[13];
  assign T78[12] = T142[12] & T79[12];
  assign T78[11] = T142[11] & T79[11];
  assign T78[10] = T142[10] & T79[10];
  assign T78[9] = T142[9] & T79[9];
  assign T78[8] = T142[8] & T79[8];
  assign T78[7] = T142[7] & T79[7];
  assign T78[6] = T142[6] & T79[6];
  assign T78[5] = T142[5] & T79[5];
  assign T78[4] = T142[4] & T79[4];
  assign T78[3] = T142[3] & T79[3];
  assign T78[2] = T142[2] & T79[2];
  assign T78[1] = T142[1] & T79[1];
  assign T78[0] = T142[0] & T79[0];
  assign T79[25] = ~T80[25];
  assign T79[24] = ~T80[24];
  assign T79[23] = ~T80[23];
  assign T79[22] = ~T80[22];
  assign T79[21] = ~T80[21];
  assign T79[20] = ~T80[20];
  assign T79[19] = ~T80[19];
  assign T79[18] = ~T80[18];
  assign T79[17] = ~T80[17];
  assign T79[16] = ~T80[16];
  assign T79[15] = ~T80[15];
  assign T79[14] = ~T80[14];
  assign T79[13] = ~T80[13];
  assign T79[12] = ~T80[12];
  assign T79[11] = ~T80[11];
  assign T79[10] = ~T80[10];
  assign T79[9] = ~T80[9];
  assign T79[8] = ~T80[8];
  assign T79[7] = ~T80[7];
  assign T79[6] = ~T80[6];
  assign T79[5] = ~T80[5];
  assign T79[4] = ~T80[4];
  assign T79[3] = ~T80[3];
  assign T79[2] = ~T80[2];
  assign T79[1] = ~T80[1];
  assign T79[0] = ~T80[0];
  assign N11 = ~T82;
  assign T80[0] = T82;
  assign T82 = T84 & T83;
  assign T83 = ~N72;
  assign T84 = N20 & N46;
  assign T86[24] = io_in_sig[26] | T129[25];
  assign T86[23] = io_in_sig[25] | T129[24];
  assign T86[22] = io_in_sig[24] | T129[23];
  assign T86[21] = io_in_sig[23] | T129[22];
  assign T86[20] = io_in_sig[22] | T129[21];
  assign T86[19] = io_in_sig[21] | T129[20];
  assign T86[18] = io_in_sig[20] | T129[19];
  assign T86[17] = io_in_sig[19] | T129[18];
  assign T86[16] = io_in_sig[18] | T129[17];
  assign T86[15] = io_in_sig[17] | T129[16];
  assign T86[14] = io_in_sig[16] | T129[15];
  assign T86[13] = io_in_sig[15] | T129[14];
  assign T86[12] = io_in_sig[14] | T129[13];
  assign T86[11] = io_in_sig[13] | T129[12];
  assign T86[10] = io_in_sig[12] | T129[11];
  assign T86[9] = io_in_sig[11] | T129[10];
  assign T86[8] = io_in_sig[10] | T129[9];
  assign T86[7] = io_in_sig[9] | T129[8];
  assign T86[6] = io_in_sig[8] | T129[7];
  assign T86[5] = io_in_sig[7] | T129[6];
  assign T86[4] = io_in_sig[6] | T129[5];
  assign T86[3] = io_in_sig[5] | T129[4];
  assign T86[2] = io_in_sig[4] | T129[3];
  assign T86[1] = io_in_sig[3] | T129[2];
  assign T86[0] = io_in_sig[2] | T129[1];
  assign T88 = T93 | T89;
  assign T89 = roundMagUp & anyRound;
  assign roundMagUp = T92 | T90;
  assign T90 = N18 & T91;
  assign T91 = ~io_in_sign;
  assign T92 = N17 & io_in_sign;
  assign T93 = N20 & N46;
  assign T140_9 = 1'b0;
  assign io_out[22] = T98[22] | T97[22];
  assign io_out[21] = T98[21] | 1'b0;
  assign io_out[20] = T98[20] | 1'b0;
  assign io_out[19] = T98[19] | 1'b0;
  assign io_out[18] = T98[18] | 1'b0;
  assign io_out[17] = T98[17] | 1'b0;
  assign io_out[16] = T98[16] | 1'b0;
  assign io_out[15] = T98[15] | 1'b0;
  assign io_out[14] = T98[14] | 1'b0;
  assign io_out[13] = T98[13] | 1'b0;
  assign io_out[12] = T98[12] | 1'b0;
  assign io_out[11] = T98[11] | 1'b0;
  assign io_out[10] = T98[10] | 1'b0;
  assign io_out[9] = T98[9] | 1'b0;
  assign io_out[8] = T98[8] | 1'b0;
  assign io_out[7] = T98[7] | 1'b0;
  assign io_out[6] = T98[6] | 1'b0;
  assign io_out[5] = T98[5] | 1'b0;
  assign io_out[4] = T98[4] | 1'b0;
  assign io_out[3] = T98[3] | 1'b0;
  assign io_out[2] = T98[2] | 1'b0;
  assign io_out[1] = T98[1] | 1'b0;
  assign io_out[0] = T98[0] | 1'b0;
  assign T98[22] = T102[22] | T99[22];
  assign T98[21] = T102[21] | T99[22];
  assign T98[20] = T102[20] | T99[22];
  assign T98[19] = T102[19] | T99[22];
  assign T98[18] = T102[18] | T99[22];
  assign T98[17] = T102[17] | T99[22];
  assign T98[16] = T102[16] | T99[22];
  assign T98[15] = T102[15] | T99[22];
  assign T98[14] = T102[14] | T99[22];
  assign T98[13] = T102[13] | T99[22];
  assign T98[12] = T102[12] | T99[22];
  assign T98[11] = T102[11] | T99[22];
  assign T98[10] = T102[10] | T99[22];
  assign T98[9] = T102[9] | T99[22];
  assign T98[8] = T102[8] | T99[22];
  assign T98[7] = T102[7] | T99[22];
  assign T98[6] = T102[6] | T99[22];
  assign T98[5] = T102[5] | T99[22];
  assign T98[4] = T102[4] | T99[22];
  assign T98[3] = T102[3] | T99[22];
  assign T98[2] = T102[2] | T99[22];
  assign T98[1] = T102[1] | T99[22];
  assign T98[0] = T102[0] | T99_0;
  assign T145[0] = T101 & T100;
  assign T100 = ~overflow_roundMagUp;
  assign overflow_roundMagUp = N20 | roundMagUp;
  assign T101 = commonCase & io_exceptionFlags[2];
  assign N12 = ~T105;
  assign N13 = ~io_in_sig[26];
  assign T70[0] = io_in_sig[26];
  assign T70[1] = N13;
  assign T105 = T106 | T97[22];
  assign T106 = common_totalUnderflow & roundMagUp;
  assign io_out[31] = T108[8] | T107[8];
  assign io_out[30] = T108[7] | T107[8];
  assign io_out[29] = T108[6] | T107[8];
  assign io_out[28] = T108[5] | 1'b0;
  assign io_out[27] = T108[4] | 1'b0;
  assign io_out[26] = T108[3] | 1'b0;
  assign io_out[25] = T108[2] | 1'b0;
  assign io_out[24] = T108[1] | 1'b0;
  assign io_out[23] = T108[0] | 1'b0;
  assign T107[8] = T97[22];
  assign T108[8] = T111[8] | T109[8];
  assign T108[7] = T111[7] | T109[8];
  assign T108[6] = T111[6] | 1'b0;
  assign T108[5] = T111[5] | 1'b0;
  assign T108[4] = T111[4] | 1'b0;
  assign T108[3] = T111[3] | 1'b0;
  assign T108[2] = T111[2] | 1'b0;
  assign T108[1] = T111[1] | 1'b0;
  assign T108[0] = T111[0] | 1'b0;
  assign T109[8] = notNaN_isInfOut;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T110;
  assign T110 = io_exceptionFlags[2] & overflow_roundMagUp;
  assign T111[8] = T113[8] | T112[8];
  assign T111[7] = T113[7] | 1'b0;
  assign T111[6] = T113[6] | T112[8];
  assign T111[5] = T113[5] | T112[8];
  assign T111[4] = T113[4] | T112[8];
  assign T111[3] = T113[3] | T112[8];
  assign T111[2] = T113[2] | T112[8];
  assign T111[1] = T113[1] | T112[8];
  assign T111[0] = T113[0] | T112[8];
  assign T112[8] = T145[0];
  assign T113[8] = T116[8] | 1'b0;
  assign T113[7] = T116[7] | 1'b0;
  assign T113[6] = T116[6] | T114[6];
  assign T113[5] = T116[5] | T114[6];
  assign T113[4] = T116[4] | 1'b0;
  assign T113[3] = T116[3] | T114[6];
  assign T113[2] = T116[2] | 1'b0;
  assign T113[1] = T116[1] | T114[6];
  assign T113[0] = T116[0] | T114[6];
  assign T114[6] = pegMinNonzeroMagOut;
  assign pegMinNonzeroMagOut = T115 & roundMagUp;
  assign T115 = commonCase & common_totalUnderflow;
  assign T116[8] = T119[8] & T117[8];
  assign T116[7] = T119[7] & T117[7];
  assign T116[6] = T119[6] & T117[6];
  assign T116[5] = T119[5] & T117[5];
  assign T116[4] = T119[4] & T117[4];
  assign T116[3] = T119[3] & T117[3];
  assign T116[2] = T119[2] & T117[2];
  assign T116[1] = T119[1] & T117[1];
  assign T116[0] = T119[0] & T117[0];
  assign T117[8] = ~1'b0;
  assign T117[7] = ~1'b0;
  assign T117[6] = ~T118[6];
  assign T117[5] = ~1'b0;
  assign T117[4] = ~1'b0;
  assign T117[3] = ~1'b0;
  assign T117[2] = ~1'b0;
  assign T117[1] = ~1'b0;
  assign T117[0] = ~1'b0;
  assign T118[6] = notNaN_isInfOut;
  assign T119[8] = T122[8] & T120[8];
  assign T119[7] = T122[7] & T120[7];
  assign T119[6] = T122[6] & T120[6];
  assign T119[5] = T122[5] & T120[5];
  assign T119[4] = T122[4] & T120[4];
  assign T119[3] = T122[3] & T120[3];
  assign T119[2] = T122[2] & T120[2];
  assign T119[1] = T122[1] & T120[1];
  assign T119[0] = T122[0] & T120[0];
  assign T120[8] = ~1'b0;
  assign T120[7] = ~T121[7];
  assign T120[6] = ~1'b0;
  assign T120[5] = ~1'b0;
  assign T120[4] = ~1'b0;
  assign T120[3] = ~1'b0;
  assign T120[2] = ~1'b0;
  assign T120[1] = ~1'b0;
  assign T120[0] = ~1'b0;
  assign T121[7] = T145[0];
  assign T122[8] = T125[8] & T123[8];
  assign T122[7] = T125[7] & T123[7];
  assign T122[6] = T125[6] & T123[6];
  assign T122[5] = T125[5] & T123[5];
  assign T122[4] = T125[4] & T123[4];
  assign T122[3] = T125[3] & T123[3];
  assign T122[2] = T125[2] & T123[2];
  assign T122[1] = T125[1] & T123[1];
  assign T122[0] = T125[0] & T123[0];
  assign T123[8] = ~T124[8];
  assign T123[7] = ~T124[8];
  assign T123[6] = ~1'b0;
  assign T123[5] = ~1'b0;
  assign T123[4] = ~T124[8];
  assign T123[3] = ~1'b0;
  assign T123[2] = ~T124[8];
  assign T123[1] = ~1'b0;
  assign T123[0] = ~1'b0;
  assign T124[8] = pegMinNonzeroMagOut;
  assign T125[8] = T71[1] & T126[8];
  assign T125[7] = T71[0] & T126[7];
  assign T125[6] = sRoundedExp[6] & T126[6];
  assign T125[5] = sRoundedExp[5] & T126[5];
  assign T125[4] = sRoundedExp[4] & T126[4];
  assign T125[3] = sRoundedExp[3] & T126[3];
  assign T125[2] = sRoundedExp[2] & T126[2];
  assign T125[1] = sRoundedExp[1] & T126[1];
  assign T125[0] = sRoundedExp[0] & T126[0];
  assign T126[8] = ~T127[8];
  assign T126[7] = ~T127[8];
  assign T126[6] = ~T127[8];
  assign T126[5] = ~1'b0;
  assign T126[4] = ~1'b0;
  assign T126[3] = ~1'b0;
  assign T126[2] = ~1'b0;
  assign T126[1] = ~1'b0;
  assign T126[0] = ~1'b0;
  assign T127[8] = T128;
  assign T128 = io_in_isZero | common_totalUnderflow;
  assign N14 = ~T97[22];

endmodule