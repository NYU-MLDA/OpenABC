module Mul54
(
  clk,
  io_val_s0,
  io_latch_a_s0,
  io_a_s0,
  io_latch_b_s0,
  io_b_s0,
  io_c_s2,
  io_result_s3
);

  input [53:0] io_a_s0;
  input [53:0] io_b_s0;
  input [104:0] io_c_s2;
  output [104:0] io_result_s3;
  input clk;
  input io_val_s0;
  input io_latch_a_s0;
  input io_latch_b_s0;
  wire T6,T9;
  wire [104:0] T1,T2;
  reg [104:0] io_result_s3;
  reg [53:0] reg_b_s2,reg_b_s1,reg_a_s2,reg_a_s1;
  reg val_s1,val_s2;

  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[104] <= T1[104];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[103] <= T1[103];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[102] <= T1[102];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[101] <= T1[101];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[100] <= T1[100];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[99] <= T1[99];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[98] <= T1[98];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[97] <= T1[97];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[96] <= T1[96];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[95] <= T1[95];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[94] <= T1[94];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[93] <= T1[93];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[92] <= T1[92];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[91] <= T1[91];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[90] <= T1[90];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[89] <= T1[89];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[88] <= T1[88];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[87] <= T1[87];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[86] <= T1[86];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[85] <= T1[85];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[84] <= T1[84];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[83] <= T1[83];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[82] <= T1[82];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[81] <= T1[81];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[80] <= T1[80];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[79] <= T1[79];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[78] <= T1[78];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[77] <= T1[77];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[76] <= T1[76];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[75] <= T1[75];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[74] <= T1[74];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[73] <= T1[73];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[72] <= T1[72];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[71] <= T1[71];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[70] <= T1[70];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[69] <= T1[69];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[68] <= T1[68];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[67] <= T1[67];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[66] <= T1[66];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[65] <= T1[65];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[64] <= T1[64];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[63] <= T1[63];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[62] <= T1[62];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[61] <= T1[61];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[60] <= T1[60];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[59] <= T1[59];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[58] <= T1[58];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[57] <= T1[57];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[56] <= T1[56];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[55] <= T1[55];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[54] <= T1[54];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[53] <= T1[53];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[52] <= T1[52];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[51] <= T1[51];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[50] <= T1[50];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[49] <= T1[49];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[48] <= T1[48];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[47] <= T1[47];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[46] <= T1[46];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[45] <= T1[45];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[44] <= T1[44];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[43] <= T1[43];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[42] <= T1[42];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[41] <= T1[41];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[40] <= T1[40];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[39] <= T1[39];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[38] <= T1[38];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[37] <= T1[37];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[36] <= T1[36];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[35] <= T1[35];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[34] <= T1[34];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[33] <= T1[33];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[32] <= T1[32];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[31] <= T1[31];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[30] <= T1[30];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[29] <= T1[29];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[28] <= T1[28];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[27] <= T1[27];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[26] <= T1[26];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[25] <= T1[25];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[24] <= T1[24];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[23] <= T1[23];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[22] <= T1[22];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[21] <= T1[21];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[20] <= T1[20];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[19] <= T1[19];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[18] <= T1[18];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[17] <= T1[17];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[16] <= T1[16];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[15] <= T1[15];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[14] <= T1[14];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[13] <= T1[13];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[12] <= T1[12];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[11] <= T1[11];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[10] <= T1[10];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[9] <= T1[9];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[8] <= T1[8];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[7] <= T1[7];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[6] <= T1[6];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[5] <= T1[5];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[4] <= T1[4];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[3] <= T1[3];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[2] <= T1[2];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[1] <= T1[1];
    end 
  end


  always @(posedge clk) begin
    if(val_s2) begin
      io_result_s3[0] <= T1[0];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[53] <= reg_b_s1[53];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[52] <= reg_b_s1[52];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[51] <= reg_b_s1[51];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[50] <= reg_b_s1[50];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[49] <= reg_b_s1[49];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[48] <= reg_b_s1[48];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[47] <= reg_b_s1[47];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[46] <= reg_b_s1[46];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[45] <= reg_b_s1[45];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[44] <= reg_b_s1[44];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[43] <= reg_b_s1[43];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[42] <= reg_b_s1[42];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[41] <= reg_b_s1[41];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[40] <= reg_b_s1[40];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[39] <= reg_b_s1[39];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[38] <= reg_b_s1[38];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[37] <= reg_b_s1[37];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[36] <= reg_b_s1[36];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[35] <= reg_b_s1[35];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[34] <= reg_b_s1[34];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[33] <= reg_b_s1[33];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[32] <= reg_b_s1[32];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[31] <= reg_b_s1[31];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[30] <= reg_b_s1[30];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[29] <= reg_b_s1[29];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[28] <= reg_b_s1[28];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[27] <= reg_b_s1[27];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[26] <= reg_b_s1[26];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[25] <= reg_b_s1[25];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[24] <= reg_b_s1[24];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[23] <= reg_b_s1[23];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[22] <= reg_b_s1[22];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[21] <= reg_b_s1[21];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[20] <= reg_b_s1[20];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[19] <= reg_b_s1[19];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[18] <= reg_b_s1[18];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[17] <= reg_b_s1[17];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[16] <= reg_b_s1[16];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[15] <= reg_b_s1[15];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[14] <= reg_b_s1[14];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[13] <= reg_b_s1[13];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[12] <= reg_b_s1[12];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[11] <= reg_b_s1[11];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[10] <= reg_b_s1[10];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[9] <= reg_b_s1[9];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[8] <= reg_b_s1[8];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[7] <= reg_b_s1[7];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[6] <= reg_b_s1[6];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[5] <= reg_b_s1[5];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[4] <= reg_b_s1[4];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[3] <= reg_b_s1[3];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[2] <= reg_b_s1[2];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[1] <= reg_b_s1[1];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_b_s2[0] <= reg_b_s1[0];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[53] <= io_b_s0[53];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[52] <= io_b_s0[52];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[51] <= io_b_s0[51];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[50] <= io_b_s0[50];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[49] <= io_b_s0[49];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[48] <= io_b_s0[48];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[47] <= io_b_s0[47];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[46] <= io_b_s0[46];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[45] <= io_b_s0[45];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[44] <= io_b_s0[44];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[43] <= io_b_s0[43];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[42] <= io_b_s0[42];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[41] <= io_b_s0[41];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[40] <= io_b_s0[40];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[39] <= io_b_s0[39];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[38] <= io_b_s0[38];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[37] <= io_b_s0[37];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[36] <= io_b_s0[36];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[35] <= io_b_s0[35];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[34] <= io_b_s0[34];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[33] <= io_b_s0[33];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[32] <= io_b_s0[32];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[31] <= io_b_s0[31];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[30] <= io_b_s0[30];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[29] <= io_b_s0[29];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[28] <= io_b_s0[28];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[27] <= io_b_s0[27];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[26] <= io_b_s0[26];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[25] <= io_b_s0[25];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[24] <= io_b_s0[24];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[23] <= io_b_s0[23];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[22] <= io_b_s0[22];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[21] <= io_b_s0[21];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[20] <= io_b_s0[20];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[19] <= io_b_s0[19];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[18] <= io_b_s0[18];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[17] <= io_b_s0[17];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[16] <= io_b_s0[16];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[15] <= io_b_s0[15];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[14] <= io_b_s0[14];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[13] <= io_b_s0[13];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[12] <= io_b_s0[12];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[11] <= io_b_s0[11];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[10] <= io_b_s0[10];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[9] <= io_b_s0[9];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[8] <= io_b_s0[8];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[7] <= io_b_s0[7];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[6] <= io_b_s0[6];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[5] <= io_b_s0[5];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[4] <= io_b_s0[4];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[3] <= io_b_s0[3];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[2] <= io_b_s0[2];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[1] <= io_b_s0[1];
    end 
  end


  always @(posedge clk) begin
    if(T6) begin
      reg_b_s1[0] <= io_b_s0[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      val_s1 <= io_val_s0;
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[53] <= reg_a_s1[53];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[52] <= reg_a_s1[52];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[51] <= reg_a_s1[51];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[50] <= reg_a_s1[50];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[49] <= reg_a_s1[49];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[48] <= reg_a_s1[48];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[47] <= reg_a_s1[47];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[46] <= reg_a_s1[46];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[45] <= reg_a_s1[45];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[44] <= reg_a_s1[44];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[43] <= reg_a_s1[43];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[42] <= reg_a_s1[42];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[41] <= reg_a_s1[41];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[40] <= reg_a_s1[40];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[39] <= reg_a_s1[39];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[38] <= reg_a_s1[38];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[37] <= reg_a_s1[37];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[36] <= reg_a_s1[36];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[35] <= reg_a_s1[35];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[34] <= reg_a_s1[34];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[33] <= reg_a_s1[33];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[32] <= reg_a_s1[32];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[31] <= reg_a_s1[31];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[30] <= reg_a_s1[30];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[29] <= reg_a_s1[29];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[28] <= reg_a_s1[28];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[27] <= reg_a_s1[27];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[26] <= reg_a_s1[26];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[25] <= reg_a_s1[25];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[24] <= reg_a_s1[24];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[23] <= reg_a_s1[23];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[22] <= reg_a_s1[22];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[21] <= reg_a_s1[21];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[20] <= reg_a_s1[20];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[19] <= reg_a_s1[19];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[18] <= reg_a_s1[18];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[17] <= reg_a_s1[17];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[16] <= reg_a_s1[16];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[15] <= reg_a_s1[15];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[14] <= reg_a_s1[14];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[13] <= reg_a_s1[13];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[12] <= reg_a_s1[12];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[11] <= reg_a_s1[11];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[10] <= reg_a_s1[10];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[9] <= reg_a_s1[9];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[8] <= reg_a_s1[8];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[7] <= reg_a_s1[7];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[6] <= reg_a_s1[6];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[5] <= reg_a_s1[5];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[4] <= reg_a_s1[4];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[3] <= reg_a_s1[3];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[2] <= reg_a_s1[2];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[1] <= reg_a_s1[1];
    end 
  end


  always @(posedge clk) begin
    if(val_s1) begin
      reg_a_s2[0] <= reg_a_s1[0];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[53] <= io_a_s0[53];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[52] <= io_a_s0[52];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[51] <= io_a_s0[51];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[50] <= io_a_s0[50];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[49] <= io_a_s0[49];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[48] <= io_a_s0[48];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[47] <= io_a_s0[47];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[46] <= io_a_s0[46];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[45] <= io_a_s0[45];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[44] <= io_a_s0[44];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[43] <= io_a_s0[43];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[42] <= io_a_s0[42];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[41] <= io_a_s0[41];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[40] <= io_a_s0[40];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[39] <= io_a_s0[39];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[38] <= io_a_s0[38];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[37] <= io_a_s0[37];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[36] <= io_a_s0[36];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[35] <= io_a_s0[35];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[34] <= io_a_s0[34];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[33] <= io_a_s0[33];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[32] <= io_a_s0[32];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[31] <= io_a_s0[31];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[30] <= io_a_s0[30];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[29] <= io_a_s0[29];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[28] <= io_a_s0[28];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[27] <= io_a_s0[27];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[26] <= io_a_s0[26];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[25] <= io_a_s0[25];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[24] <= io_a_s0[24];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[23] <= io_a_s0[23];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[22] <= io_a_s0[22];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[21] <= io_a_s0[21];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[20] <= io_a_s0[20];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[19] <= io_a_s0[19];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[18] <= io_a_s0[18];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[17] <= io_a_s0[17];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[16] <= io_a_s0[16];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[15] <= io_a_s0[15];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[14] <= io_a_s0[14];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[13] <= io_a_s0[13];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[12] <= io_a_s0[12];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[11] <= io_a_s0[11];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[10] <= io_a_s0[10];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[9] <= io_a_s0[9];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[8] <= io_a_s0[8];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[7] <= io_a_s0[7];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[6] <= io_a_s0[6];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[5] <= io_a_s0[5];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[4] <= io_a_s0[4];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[3] <= io_a_s0[3];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[2] <= io_a_s0[2];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[1] <= io_a_s0[1];
    end 
  end


  always @(posedge clk) begin
    if(T9) begin
      reg_a_s1[0] <= io_a_s0[0];
    end 
  end


  always @(posedge clk) begin
    if(1'b1) begin
      val_s2 <= val_s1;
    end 
  end

  assign T2 = reg_a_s2 * reg_b_s2;
  assign T1 = T2 + io_c_s2;
  assign T6 = io_val_s0 & io_latch_b_s0;
  assign T9 = io_val_s0 & io_latch_a_s0;

endmodule