module arbiter_00000003_64
(
  clk_i,
  rst_ni,
  data_req_i,
  address_i,
  data_wdata_i,
  data_we_i,
  data_be_i,
  data_size_i,
  data_gnt_o,
  data_rvalid_o,
  data_rdata_o,
  id_i,
  id_o,
  gnt_id_i,
  data_req_o,
  address_o,
  data_wdata_o,
  data_we_o,
  data_be_o,
  data_size_o,
  data_gnt_i,
  data_rvalid_i,
  data_rdata_i
);

  input [2:0] data_req_i;
  input [191:0] address_i;
  input [191:0] data_wdata_i;
  input [2:0] data_we_i;
  input [23:0] data_be_i;
  input [5:0] data_size_i;
  output [2:0] data_gnt_o;
  output [2:0] data_rvalid_o;
  output [191:0] data_rdata_o;
  input [1:0] id_i;
  output [1:0] id_o;
  input [1:0] gnt_id_i;
  output [63:0] address_o;
  output [63:0] data_wdata_o;
  output [7:0] data_be_o;
  output [1:0] data_size_o;
  input [63:0] data_rdata_i;
  input clk_i;
  input rst_ni;
  input data_gnt_i;
  input data_rvalid_i;
  output data_req_o;
  output data_we_o;
  wire [2:0] data_gnt_o,data_rvalid_o;
  wire [191:0] data_rdata_o;
  wire [1:0] id_o,data_size_o,state_d;
  wire [63:0] address_o,data_wdata_o;
  wire [7:0] data_be_o;
  wire data_req_o,data_we_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,
  N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,
  N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,
  N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,
  N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,
  N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,
  N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,
  N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,
  N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,
  N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,
  N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,
  N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,
  N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,
  N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,
  N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,
  N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,
  N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,
  N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,
  N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,
  N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,
  N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,
  N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,
  N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,
  N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,
  N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,
  N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,
  N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,
  N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,
  N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,
  N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,
  N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,
  N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,
  N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,
  N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,
  N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,
  N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,
  N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,
  N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,
  N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,
  N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,
  N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,
  N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,
  N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,
  N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,
  N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
  N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,
  N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,
  N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,
  N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,
  N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,
  N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,
  N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,
  N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,
  N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,
  N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,
  N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,
  N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,
  N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,
  N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,
  N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,
  N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,
  N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,
  N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,
  N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,
  N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,
  N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,
  N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,
  N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,
  N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,
  N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,
  N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,
  N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,
  N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,
  N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,
  N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,
  N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,
  N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,
  N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230;
  reg [140:0] req_q;
  reg [1:0] state_q;
  assign N39 = N37 & N38;
  assign N40 = N37 | state_q[0];

  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[140] <= 1'b0;
    end else if(N1225) begin
      req_q[140] <= N1072;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[139] <= 1'b0;
    end else if(N1227) begin
      req_q[139] <= N1071;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[138] <= 1'b0;
    end else if(N1227) begin
      req_q[138] <= N1070;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[137] <= 1'b0;
    end else if(N1227) begin
      req_q[137] <= N1069;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[136] <= 1'b0;
    end else if(N1227) begin
      req_q[136] <= N1068;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[135] <= 1'b0;
    end else if(N1227) begin
      req_q[135] <= N1067;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[134] <= 1'b0;
    end else if(N1227) begin
      req_q[134] <= N1066;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[133] <= 1'b0;
    end else if(N1227) begin
      req_q[133] <= N1065;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[132] <= 1'b0;
    end else if(N1227) begin
      req_q[132] <= N1064;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[131] <= 1'b0;
    end else if(N1227) begin
      req_q[131] <= N1063;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[130] <= 1'b0;
    end else if(N1227) begin
      req_q[130] <= N1062;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[129] <= 1'b0;
    end else if(N1227) begin
      req_q[129] <= N1061;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[128] <= 1'b0;
    end else if(N1227) begin
      req_q[128] <= N1060;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[127] <= 1'b0;
    end else if(N1227) begin
      req_q[127] <= N1059;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[126] <= 1'b0;
    end else if(N1227) begin
      req_q[126] <= N1058;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[125] <= 1'b0;
    end else if(N1227) begin
      req_q[125] <= N1057;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[124] <= 1'b0;
    end else if(N1227) begin
      req_q[124] <= N1056;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[123] <= 1'b0;
    end else if(N1227) begin
      req_q[123] <= N1055;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[122] <= 1'b0;
    end else if(N1227) begin
      req_q[122] <= N1054;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[121] <= 1'b0;
    end else if(N1227) begin
      req_q[121] <= N1053;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[120] <= 1'b0;
    end else if(N1227) begin
      req_q[120] <= N1052;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[119] <= 1'b0;
    end else if(N1227) begin
      req_q[119] <= N1051;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[118] <= 1'b0;
    end else if(N1227) begin
      req_q[118] <= N1050;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[117] <= 1'b0;
    end else if(N1227) begin
      req_q[117] <= N1049;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[116] <= 1'b0;
    end else if(N1227) begin
      req_q[116] <= N1048;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[115] <= 1'b0;
    end else if(N1227) begin
      req_q[115] <= N1047;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[114] <= 1'b0;
    end else if(N1227) begin
      req_q[114] <= N1046;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[113] <= 1'b0;
    end else if(N1227) begin
      req_q[113] <= N1045;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[112] <= 1'b0;
    end else if(N1227) begin
      req_q[112] <= N1044;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[111] <= 1'b0;
    end else if(N1227) begin
      req_q[111] <= N1043;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[110] <= 1'b0;
    end else if(N1227) begin
      req_q[110] <= N1042;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[109] <= 1'b0;
    end else if(N1227) begin
      req_q[109] <= N1041;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[108] <= 1'b0;
    end else if(N1227) begin
      req_q[108] <= N1040;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[107] <= 1'b0;
    end else if(N1227) begin
      req_q[107] <= N1039;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[106] <= 1'b0;
    end else if(N1227) begin
      req_q[106] <= N1038;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[105] <= 1'b0;
    end else if(N1227) begin
      req_q[105] <= N1037;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[104] <= 1'b0;
    end else if(N1227) begin
      req_q[104] <= N1036;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[103] <= 1'b0;
    end else if(N1227) begin
      req_q[103] <= N1035;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[102] <= 1'b0;
    end else if(N1227) begin
      req_q[102] <= N1034;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[101] <= 1'b0;
    end else if(N1227) begin
      req_q[101] <= N1033;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[100] <= 1'b0;
    end else if(N1227) begin
      req_q[100] <= N1032;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[99] <= 1'b0;
    end else if(N1227) begin
      req_q[99] <= N1031;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[98] <= 1'b0;
    end else if(N1225) begin
      req_q[98] <= N1030;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[97] <= 1'b0;
    end else if(N1225) begin
      req_q[97] <= N1029;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[96] <= 1'b0;
    end else if(N1225) begin
      req_q[96] <= N1028;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[95] <= 1'b0;
    end else if(N1225) begin
      req_q[95] <= N1027;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[94] <= 1'b0;
    end else if(N1225) begin
      req_q[94] <= N1026;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[93] <= 1'b0;
    end else if(N1225) begin
      req_q[93] <= N1025;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[92] <= 1'b0;
    end else if(N1225) begin
      req_q[92] <= N1024;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[91] <= 1'b0;
    end else if(N1225) begin
      req_q[91] <= N1023;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[90] <= 1'b0;
    end else if(N1225) begin
      req_q[90] <= N1022;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[89] <= 1'b0;
    end else if(N1225) begin
      req_q[89] <= N1021;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[88] <= 1'b0;
    end else if(N1225) begin
      req_q[88] <= N1020;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[87] <= 1'b0;
    end else if(N1225) begin
      req_q[87] <= N1019;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[86] <= 1'b0;
    end else if(N1225) begin
      req_q[86] <= N1018;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[85] <= 1'b0;
    end else if(N1225) begin
      req_q[85] <= N1017;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[84] <= 1'b0;
    end else if(N1225) begin
      req_q[84] <= N1016;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[83] <= 1'b0;
    end else if(N1225) begin
      req_q[83] <= N1015;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[82] <= 1'b0;
    end else if(N1225) begin
      req_q[82] <= N1014;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[81] <= 1'b0;
    end else if(N1225) begin
      req_q[81] <= N1013;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[80] <= 1'b0;
    end else if(N1225) begin
      req_q[80] <= N1012;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[79] <= 1'b0;
    end else if(N1225) begin
      req_q[79] <= N1011;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[78] <= 1'b0;
    end else if(N1225) begin
      req_q[78] <= N1010;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[77] <= 1'b0;
    end else if(N1225) begin
      req_q[77] <= N1009;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[76] <= 1'b0;
    end else if(N1225) begin
      req_q[76] <= N1008;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[75] <= 1'b0;
    end else if(N1225) begin
      req_q[75] <= N1007;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[74] <= 1'b0;
    end else if(N1225) begin
      req_q[74] <= N1006;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[73] <= 1'b0;
    end else if(N1225) begin
      req_q[73] <= N1005;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[72] <= 1'b0;
    end else if(N1225) begin
      req_q[72] <= N1004;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[71] <= 1'b0;
    end else if(N1225) begin
      req_q[71] <= N1003;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[70] <= 1'b0;
    end else if(N1225) begin
      req_q[70] <= N1002;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[69] <= 1'b0;
    end else if(N1225) begin
      req_q[69] <= N1001;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[68] <= 1'b0;
    end else if(N1225) begin
      req_q[68] <= N1000;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[67] <= 1'b0;
    end else if(N1225) begin
      req_q[67] <= N999;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[66] <= 1'b0;
    end else if(N1225) begin
      req_q[66] <= N998;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[65] <= 1'b0;
    end else if(N1225) begin
      req_q[65] <= N997;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[64] <= 1'b0;
    end else if(N1225) begin
      req_q[64] <= N996;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[63] <= 1'b0;
    end else if(N1225) begin
      req_q[63] <= N995;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[62] <= 1'b0;
    end else if(N1225) begin
      req_q[62] <= N994;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[61] <= 1'b0;
    end else if(N1225) begin
      req_q[61] <= N993;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[60] <= 1'b0;
    end else if(N1225) begin
      req_q[60] <= N992;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[59] <= 1'b0;
    end else if(N1225) begin
      req_q[59] <= N991;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[58] <= 1'b0;
    end else if(N1225) begin
      req_q[58] <= N990;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[57] <= 1'b0;
    end else if(N1225) begin
      req_q[57] <= N989;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[56] <= 1'b0;
    end else if(N1225) begin
      req_q[56] <= N988;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[55] <= 1'b0;
    end else if(N1225) begin
      req_q[55] <= N987;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[54] <= 1'b0;
    end else if(N1225) begin
      req_q[54] <= N986;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[53] <= 1'b0;
    end else if(N1225) begin
      req_q[53] <= N985;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[52] <= 1'b0;
    end else if(N1225) begin
      req_q[52] <= N984;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[51] <= 1'b0;
    end else if(N1225) begin
      req_q[51] <= N983;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[50] <= 1'b0;
    end else if(N1225) begin
      req_q[50] <= N982;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[49] <= 1'b0;
    end else if(N1225) begin
      req_q[49] <= N981;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[48] <= 1'b0;
    end else if(N1225) begin
      req_q[48] <= N980;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[47] <= 1'b0;
    end else if(N1225) begin
      req_q[47] <= N979;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[46] <= 1'b0;
    end else if(N1225) begin
      req_q[46] <= N978;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[45] <= 1'b0;
    end else if(N1225) begin
      req_q[45] <= N977;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[44] <= 1'b0;
    end else if(N1225) begin
      req_q[44] <= N976;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[43] <= 1'b0;
    end else if(N1225) begin
      req_q[43] <= N975;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[42] <= 1'b0;
    end else if(N1225) begin
      req_q[42] <= N974;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[41] <= 1'b0;
    end else if(N1225) begin
      req_q[41] <= N973;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[40] <= 1'b0;
    end else if(N1225) begin
      req_q[40] <= N972;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[39] <= 1'b0;
    end else if(N1225) begin
      req_q[39] <= N971;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[38] <= 1'b0;
    end else if(N1225) begin
      req_q[38] <= N970;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[37] <= 1'b0;
    end else if(N1225) begin
      req_q[37] <= N969;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[36] <= 1'b0;
    end else if(N1225) begin
      req_q[36] <= N968;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[35] <= 1'b0;
    end else if(N1225) begin
      req_q[35] <= N967;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[34] <= 1'b0;
    end else if(N1225) begin
      req_q[34] <= N966;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[33] <= 1'b0;
    end else if(N1225) begin
      req_q[33] <= N965;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[32] <= 1'b0;
    end else if(N1225) begin
      req_q[32] <= N964;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[31] <= 1'b0;
    end else if(N1225) begin
      req_q[31] <= N963;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[30] <= 1'b0;
    end else if(N1225) begin
      req_q[30] <= N962;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[29] <= 1'b0;
    end else if(N1225) begin
      req_q[29] <= N961;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[28] <= 1'b0;
    end else if(N1225) begin
      req_q[28] <= N960;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[27] <= 1'b0;
    end else if(N1225) begin
      req_q[27] <= N959;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[26] <= 1'b0;
    end else if(N1225) begin
      req_q[26] <= N958;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[25] <= 1'b0;
    end else if(N1225) begin
      req_q[25] <= N957;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[24] <= 1'b0;
    end else if(N1225) begin
      req_q[24] <= N956;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[23] <= 1'b0;
    end else if(N1225) begin
      req_q[23] <= N955;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[22] <= 1'b0;
    end else if(N1225) begin
      req_q[22] <= N954;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[21] <= 1'b0;
    end else if(N1225) begin
      req_q[21] <= N953;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[20] <= 1'b0;
    end else if(N1225) begin
      req_q[20] <= N952;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[19] <= 1'b0;
    end else if(N1225) begin
      req_q[19] <= N951;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[18] <= 1'b0;
    end else if(N1225) begin
      req_q[18] <= N950;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[17] <= 1'b0;
    end else if(N1225) begin
      req_q[17] <= N949;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[16] <= 1'b0;
    end else if(N1225) begin
      req_q[16] <= N948;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[15] <= 1'b0;
    end else if(N1225) begin
      req_q[15] <= N947;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[14] <= 1'b0;
    end else if(N1225) begin
      req_q[14] <= N946;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[13] <= 1'b0;
    end else if(N1225) begin
      req_q[13] <= N945;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[12] <= 1'b0;
    end else if(N1225) begin
      req_q[12] <= N944;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[11] <= 1'b0;
    end else if(N1225) begin
      req_q[11] <= N943;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[10] <= 1'b0;
    end else if(N1225) begin
      req_q[10] <= N942;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[9] <= 1'b0;
    end else if(N1225) begin
      req_q[9] <= N941;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[8] <= 1'b0;
    end else if(N1225) begin
      req_q[8] <= N940;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[7] <= 1'b0;
    end else if(N1225) begin
      req_q[7] <= N939;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[6] <= 1'b0;
    end else if(N1225) begin
      req_q[6] <= N938;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[5] <= 1'b0;
    end else if(N1225) begin
      req_q[5] <= N937;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[4] <= 1'b0;
    end else if(N1225) begin
      req_q[4] <= N936;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[3] <= 1'b0;
    end else if(N1225) begin
      req_q[3] <= N935;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[2] <= 1'b0;
    end else if(N1225) begin
      req_q[2] <= N934;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[1] <= 1'b0;
    end else if(N1225) begin
      req_q[1] <= N933;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      req_q[0] <= 1'b0;
    end else if(N1225) begin
      req_q[0] <= N932;
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      state_q[1] <= 1'b0;
    end else if(N1230) begin
      state_q[1] <= state_d[1];
    end 
  end


  always @(posedge clk_i or posedge N1223) begin
    if(N1223) begin
      state_q[0] <= 1'b0;
    end else if(N1230) begin
      state_q[0] <= state_d[0];
    end 
  end

  assign N33 = N0 & req_q[140];
  assign N0 = ~req_q[139];
  assign N32 = req_q[139] & N1;
  assign N1 = ~req_q[140];
  assign N31 = N2 & N3;
  assign N2 = ~req_q[139];
  assign N3 = ~req_q[140];
  assign N1219 = N4 & req_q[140];
  assign N4 = ~req_q[139];
  assign N1218 = req_q[139] & N5;
  assign N5 = ~req_q[140];
  assign N1217 = N6 & N7;
  assign N6 = ~req_q[139];
  assign N7 = ~req_q[140];
  assign N1073 = N8 & N9;
  assign N8 = ~N1214;
  assign N9 = ~N1213;
  assign N1138 = N10 & N11;
  assign N10 = ~N1214;
  assign N11 = ~N1213;
  assign { data_rdata_o[0:0], data_rdata_o[1:1], data_rdata_o[2:2], data_rdata_o[3:3], data_rdata_o[4:4], data_rdata_o[5:5], data_rdata_o[6:6], data_rdata_o[7:7], data_rdata_o[8:8], data_rdata_o[9:9], data_rdata_o[10:10], data_rdata_o[11:11], data_rdata_o[12:12], data_rdata_o[13:13], data_rdata_o[14:14], data_rdata_o[15:15], data_rdata_o[16:16], data_rdata_o[17:17], data_rdata_o[18:18], data_rdata_o[19:19], data_rdata_o[20:20], data_rdata_o[21:21], data_rdata_o[22:22], data_rdata_o[23:23], data_rdata_o[24:24], data_rdata_o[25:25], data_rdata_o[26:26], data_rdata_o[27:27], data_rdata_o[28:28], data_rdata_o[29:29], data_rdata_o[30:30], data_rdata_o[31:31], data_rdata_o[32:32], data_rdata_o[33:33], data_rdata_o[34:34], data_rdata_o[35:35], data_rdata_o[36:36], data_rdata_o[37:37], data_rdata_o[38:38], data_rdata_o[39:39], data_rdata_o[40:40], data_rdata_o[41:41], data_rdata_o[42:42], data_rdata_o[43:43], data_rdata_o[44:44], data_rdata_o[45:45], data_rdata_o[46:46], data_rdata_o[47:47], data_rdata_o[48:48], data_rdata_o[49:49], data_rdata_o[50:50], data_rdata_o[51:51], data_rdata_o[52:52], data_rdata_o[53:53], data_rdata_o[54:54], data_rdata_o[55:55], data_rdata_o[56:56], data_rdata_o[57:57], data_rdata_o[58:58], data_rdata_o[59:59], data_rdata_o[60:60], data_rdata_o[61:61], data_rdata_o[62:62], data_rdata_o[63:63] } = (N12)? { data_rdata_i[0:0], data_rdata_i[1:1], data_rdata_i[2:2], data_rdata_i[3:3], data_rdata_i[4:4], data_rdata_i[5:5], data_rdata_i[6:6], data_rdata_i[7:7], data_rdata_i[8:8], data_rdata_i[9:9], data_rdata_i[10:10], data_rdata_i[11:11], data_rdata_i[12:12], data_rdata_i[13:13], data_rdata_i[14:14], data_rdata_i[15:15], data_rdata_i[16:16], data_rdata_i[17:17], data_rdata_i[18:18], data_rdata_i[19:19], data_rdata_i[20:20], data_rdata_i[21:21], data_rdata_i[22:22], data_rdata_i[23:23], data_rdata_i[24:24], data_rdata_i[25:25], data_rdata_i[26:26], data_rdata_i[27:27], data_rdata_i[28:28], data_rdata_i[29:29], data_rdata_i[30:30], data_rdata_i[31:31], data_rdata_i[32:32], data_rdata_i[33:33], data_rdata_i[34:34], data_rdata_i[35:35], data_rdata_i[36:36], data_rdata_i[37:37], data_rdata_i[38:38], data_rdata_i[39:39], data_rdata_i[40:40], data_rdata_i[41:41], data_rdata_i[42:42], data_rdata_i[43:43], data_rdata_i[44:44], data_rdata_i[45:45], data_rdata_i[46:46], data_rdata_i[47:47], data_rdata_i[48:48], data_rdata_i[49:49], data_rdata_i[50:50], data_rdata_i[51:51], data_rdata_i[52:52], data_rdata_i[53:53], data_rdata_i[54:54], data_rdata_i[55:55], data_rdata_i[56:56], data_rdata_i[57:57], data_rdata_i[58:58], data_rdata_i[59:59], data_rdata_i[60:60], data_rdata_i[61:61], data_rdata_i[62:62], data_rdata_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N31;
  assign { data_rdata_o[64:64], data_rdata_o[65:65], data_rdata_o[66:66], data_rdata_o[67:67], data_rdata_o[68:68], data_rdata_o[69:69], data_rdata_o[70:70], data_rdata_o[71:71], data_rdata_o[72:72], data_rdata_o[73:73], data_rdata_o[74:74], data_rdata_o[75:75], data_rdata_o[76:76], data_rdata_o[77:77], data_rdata_o[78:78], data_rdata_o[79:79], data_rdata_o[80:80], data_rdata_o[81:81], data_rdata_o[82:82], data_rdata_o[83:83], data_rdata_o[84:84], data_rdata_o[85:85], data_rdata_o[86:86], data_rdata_o[87:87], data_rdata_o[88:88], data_rdata_o[89:89], data_rdata_o[90:90], data_rdata_o[91:91], data_rdata_o[92:92], data_rdata_o[93:93], data_rdata_o[94:94], data_rdata_o[95:95], data_rdata_o[96:96], data_rdata_o[97:97], data_rdata_o[98:98], data_rdata_o[99:99], data_rdata_o[100:100], data_rdata_o[101:101], data_rdata_o[102:102], data_rdata_o[103:103], data_rdata_o[104:104], data_rdata_o[105:105], data_rdata_o[106:106], data_rdata_o[107:107], data_rdata_o[108:108], data_rdata_o[109:109], data_rdata_o[110:110], data_rdata_o[111:111], data_rdata_o[112:112], data_rdata_o[113:113], data_rdata_o[114:114], data_rdata_o[115:115], data_rdata_o[116:116], data_rdata_o[117:117], data_rdata_o[118:118], data_rdata_o[119:119], data_rdata_o[120:120], data_rdata_o[121:121], data_rdata_o[122:122], data_rdata_o[123:123], data_rdata_o[124:124], data_rdata_o[125:125], data_rdata_o[126:126], data_rdata_o[127:127] } = (N13)? { data_rdata_i[0:0], data_rdata_i[1:1], data_rdata_i[2:2], data_rdata_i[3:3], data_rdata_i[4:4], data_rdata_i[5:5], data_rdata_i[6:6], data_rdata_i[7:7], data_rdata_i[8:8], data_rdata_i[9:9], data_rdata_i[10:10], data_rdata_i[11:11], data_rdata_i[12:12], data_rdata_i[13:13], data_rdata_i[14:14], data_rdata_i[15:15], data_rdata_i[16:16], data_rdata_i[17:17], data_rdata_i[18:18], data_rdata_i[19:19], data_rdata_i[20:20], data_rdata_i[21:21], data_rdata_i[22:22], data_rdata_i[23:23], data_rdata_i[24:24], data_rdata_i[25:25], data_rdata_i[26:26], data_rdata_i[27:27], data_rdata_i[28:28], data_rdata_i[29:29], data_rdata_i[30:30], data_rdata_i[31:31], data_rdata_i[32:32], data_rdata_i[33:33], data_rdata_i[34:34], data_rdata_i[35:35], data_rdata_i[36:36], data_rdata_i[37:37], data_rdata_i[38:38], data_rdata_i[39:39], data_rdata_i[40:40], data_rdata_i[41:41], data_rdata_i[42:42], data_rdata_i[43:43], data_rdata_i[44:44], data_rdata_i[45:45], data_rdata_i[46:46], data_rdata_i[47:47], data_rdata_i[48:48], data_rdata_i[49:49], data_rdata_i[50:50], data_rdata_i[51:51], data_rdata_i[52:52], data_rdata_i[53:53], data_rdata_i[54:54], data_rdata_i[55:55], data_rdata_i[56:56], data_rdata_i[57:57], data_rdata_i[58:58], data_rdata_i[59:59], data_rdata_i[60:60], data_rdata_i[61:61], data_rdata_i[62:62], data_rdata_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      (N35)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N13 = N32;
  assign { data_rdata_o[128:128], data_rdata_o[129:129], data_rdata_o[130:130], data_rdata_o[131:131], data_rdata_o[132:132], data_rdata_o[133:133], data_rdata_o[134:134], data_rdata_o[135:135], data_rdata_o[136:136], data_rdata_o[137:137], data_rdata_o[138:138], data_rdata_o[139:139], data_rdata_o[140:140], data_rdata_o[141:141], data_rdata_o[142:142], data_rdata_o[143:143], data_rdata_o[144:144], data_rdata_o[145:145], data_rdata_o[146:146], data_rdata_o[147:147], data_rdata_o[148:148], data_rdata_o[149:149], data_rdata_o[150:150], data_rdata_o[151:151], data_rdata_o[152:152], data_rdata_o[153:153], data_rdata_o[154:154], data_rdata_o[155:155], data_rdata_o[156:156], data_rdata_o[157:157], data_rdata_o[158:158], data_rdata_o[159:159], data_rdata_o[160:160], data_rdata_o[161:161], data_rdata_o[162:162], data_rdata_o[163:163], data_rdata_o[164:164], data_rdata_o[165:165], data_rdata_o[166:166], data_rdata_o[167:167], data_rdata_o[168:168], data_rdata_o[169:169], data_rdata_o[170:170], data_rdata_o[171:171], data_rdata_o[172:172], data_rdata_o[173:173], data_rdata_o[174:174], data_rdata_o[175:175], data_rdata_o[176:176], data_rdata_o[177:177], data_rdata_o[178:178], data_rdata_o[179:179], data_rdata_o[180:180], data_rdata_o[181:181], data_rdata_o[182:182], data_rdata_o[183:183], data_rdata_o[184:184], data_rdata_o[185:185], data_rdata_o[186:186], data_rdata_o[187:187], data_rdata_o[188:188], data_rdata_o[189:189], data_rdata_o[190:190], data_rdata_o[191:191] } = (N14)? { data_rdata_i[0:0], data_rdata_i[1:1], data_rdata_i[2:2], data_rdata_i[3:3], data_rdata_i[4:4], data_rdata_i[5:5], data_rdata_i[6:6], data_rdata_i[7:7], data_rdata_i[8:8], data_rdata_i[9:9], data_rdata_i[10:10], data_rdata_i[11:11], data_rdata_i[12:12], data_rdata_i[13:13], data_rdata_i[14:14], data_rdata_i[15:15], data_rdata_i[16:16], data_rdata_i[17:17], data_rdata_i[18:18], data_rdata_i[19:19], data_rdata_i[20:20], data_rdata_i[21:21], data_rdata_i[22:22], data_rdata_i[23:23], data_rdata_i[24:24], data_rdata_i[25:25], data_rdata_i[26:26], data_rdata_i[27:27], data_rdata_i[28:28], data_rdata_i[29:29], data_rdata_i[30:30], data_rdata_i[31:31], data_rdata_i[32:32], data_rdata_i[33:33], data_rdata_i[34:34], data_rdata_i[35:35], data_rdata_i[36:36], data_rdata_i[37:37], data_rdata_i[38:38], data_rdata_i[39:39], data_rdata_i[40:40], data_rdata_i[41:41], data_rdata_i[42:42], data_rdata_i[43:43], data_rdata_i[44:44], data_rdata_i[45:45], data_rdata_i[46:46], data_rdata_i[47:47], data_rdata_i[48:48], data_rdata_i[49:49], data_rdata_i[50:50], data_rdata_i[51:51], data_rdata_i[52:52], data_rdata_i[53:53], data_rdata_i[54:54], data_rdata_i[55:55], data_rdata_i[56:56], data_rdata_i[57:57], data_rdata_i[58:58], data_rdata_i[59:59], data_rdata_i[60:60], data_rdata_i[61:61], data_rdata_i[62:62], data_rdata_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N36)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N14 = N33;
  assign N43 = (N15)? data_req_i[0] : 
               (N42)? 1'b0 : 1'b0;
  assign N15 = data_req_i[0];
  assign { N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44 } = (N15)? { 1'b0, 1'b0, address_i[63:0], data_wdata_i[63:0], data_size_i[1:0], data_be_i[7:0], data_we_i[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N42)? req_q : 1'b0;
  assign { N186, N185 } = (N15)? { 1'b1, 1'b0 } : 
                          (N42)? state_q : 1'b0;
  assign N187 = ~data_req_i[0];
  assign N190 = (N16)? data_req_i[1] : 
                (N189)? N43 : 1'b0;
  assign N16 = data_req_i[1];
  assign N191 = (N16)? data_req_i[1] : 
                (N189)? 1'b0 : 1'b0;
  assign { N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192 } = (N16)? { 1'b0, 1'b1, address_i[127:64], data_wdata_i[127:64], data_size_i[3:2], data_be_i[15:8], data_we_i[1:1] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N189)? { N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44 } : 1'b0;
  assign { N334, N333 } = (N16)? { 1'b1, 1'b0 } : 
                          (N189)? { N186, N185 } : 1'b0;
  assign N335 = (N16)? 1'b0 : 
                (N189)? N187 : 1'b0;
  assign N338 = (N17)? data_req_i[2] : 
                (N337)? N190 : 1'b0;
  assign N17 = data_req_i[2];
  assign N339 = (N17)? data_req_i[2] : 
                (N337)? 1'b0 : 1'b0;
  assign N340 = (N17)? 1'b0 : 
                (N337)? data_req_i[1] : 1'b0;
  assign { N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341 } = (N17)? { 1'b1, 1'b0, address_i[191:128], data_wdata_i[191:128], data_size_i[5:4], data_be_i[23:16], data_we_i[2:2] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N337)? { N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192 } : 1'b0;
  assign { N483, N482 } = (N17)? { 1'b1, 1'b0 } : 
                          (N337)? { N334, N333 } : 1'b0;
  assign { N486, N485 } = (N18)? { N483, N482 } : 
                          (N484)? { N334, N333 } : 1'b0;
  assign N18 = N335;
  assign N487 = (N18)? N338 : 
                (N484)? N190 : 1'b0;
  assign N488 = (N18)? N339 : 
                (N484)? 1'b0 : 1'b0;
  assign { N490, N489 } = (N18)? { data_req_i[2:2], N340 } : 
                          (N484)? { 1'b0, data_req_i[1:1] } : 1'b0;
  assign { N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491 } = (N18)? { N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N484)? { N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192 } : 1'b0;
  assign { N633, N632 } = (N18)? { N486, N485 } : 
                          (N19)? { N334, N333 } : 1'b0;
  assign N19 = N336;
  assign N634 = (N18)? N487 : 
                (N19)? N190 : 1'b0;
  assign N635 = (N18)? N488 : 
                (N19)? 1'b0 : 1'b0;
  assign { N637, N636 } = (N18)? { N490, N489 } : 
                          (N19)? { 1'b0, data_req_i[1:1] } : 1'b0;
  assign { N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } = (N18)? { N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N19)? { N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192 } : 1'b0;
  assign { N780, N779 } = (N20)? { N633, N632 } : 
                          (N15)? { N186, N185 } : 1'b0;
  assign N20 = N188;
  assign N781 = (N20)? N634 : 
                (N15)? N43 : 1'b0;
  assign { N783, N782 } = (N20)? { N635, N191 } : 
                          (N15)? { 1'b0, 1'b0 } : 1'b0;
  assign { N785, N784 } = (N20)? { N637, N636 } : 
                          (N15)? { 1'b0, 1'b0 } : 1'b0;
  assign { N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786 } = (N20)? { N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N15)? { N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44 } : 1'b0;
  assign { N928, N927 } = (N21)? { N780, N779 } : 
                          (N15)? { N186, N185 } : 1'b0;
  assign N21 = N187;
  assign N929 = (N21)? N781 : 
                (N15)? N43 : 1'b0;
  assign { N931, N930 } = (N21)? { N783, N782 } : 
                          (N15)? { 1'b0, 1'b0 } : 1'b0;
  assign { N1213, N1214 } = (N21)? { N785, N784 } : 
                            (N15)? { 1'b0, 1'b0 } : 1'b0;
  assign { N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932 } = (N21)? { N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N15)? { N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44 } : 1'b0;
  assign { N1222, N1221, N1220 } = (N22)? { N1219, N1218, N1217 } : 
                                   (N23)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = data_rvalid_i;
  assign N23 = N1216;
  assign state_d = (N24)? { N928, N927 } : 
                   (N25)? { 1'b0, 1'b0 } : 1'b0;
  assign N24 = N39;
  assign N25 = N41;
  assign data_gnt_o = (N24)? { N931, N930, N43 } : 
                      (N25)? { 1'b0, 1'b0, 1'b0 } : 
                      (N26)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = state_q[0];
  assign data_req_o = (N24)? N929 : 
                      (N25)? 1'b1 : 
                      (N26)? 1'b0 : 1'b0;
  assign id_o = (N24)? { N1213, N1214 } : 
                (N25)? req_q[140:139] : 
                (N26)? req_q[140:139] : 1'b0;
  assign address_o = (N24)? { N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137 } : 
                     (N25)? req_q[138:75] : 
                     (N26)? req_q[138:75] : 1'b0;
  assign data_wdata_o = (N24)? { N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202 } : 
                        (N25)? req_q[74:11] : 
                        (N26)? req_q[74:11] : 1'b0;
  assign data_be_o = (N24)? { N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210 } : 
                     (N25)? req_q[8:1] : 
                     (N26)? req_q[8:1] : 1'b0;
  assign data_size_o = (N24)? { N1211, N1212 } : 
                       (N25)? req_q[10:9] : 
                       (N26)? req_q[10:9] : 1'b0;
  assign data_we_o = (N24)? N1215 : 
                     (N25)? req_q[0] : 
                     (N26)? req_q[0] : 1'b0;
  assign data_rvalid_o = (N24)? { 1'b0, 1'b0, 1'b0 } : 
                         (N25)? { N1222, N1221, N1220 } : 
                         (N26)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1074 = (N27)? address_i[63] : 
                 (N28)? address_i[127] : 
                 (N29)? address_i[191] : 1'b0;
  assign N27 = N1073;
  assign N28 = N1214;
  assign N29 = N1213;
  assign N1075 = (N27)? address_i[62] : 
                 (N28)? address_i[126] : 
                 (N29)? address_i[190] : 1'b0;
  assign N1076 = (N27)? address_i[61] : 
                 (N28)? address_i[125] : 
                 (N29)? address_i[189] : 1'b0;
  assign N1077 = (N27)? address_i[60] : 
                 (N28)? address_i[124] : 
                 (N29)? address_i[188] : 1'b0;
  assign N1078 = (N27)? address_i[59] : 
                 (N28)? address_i[123] : 
                 (N29)? address_i[187] : 1'b0;
  assign N1079 = (N27)? address_i[58] : 
                 (N28)? address_i[122] : 
                 (N29)? address_i[186] : 1'b0;
  assign N1080 = (N27)? address_i[57] : 
                 (N28)? address_i[121] : 
                 (N29)? address_i[185] : 1'b0;
  assign N1081 = (N27)? address_i[56] : 
                 (N28)? address_i[120] : 
                 (N29)? address_i[184] : 1'b0;
  assign N1082 = (N27)? address_i[55] : 
                 (N28)? address_i[119] : 
                 (N29)? address_i[183] : 1'b0;
  assign N1083 = (N27)? address_i[54] : 
                 (N28)? address_i[118] : 
                 (N29)? address_i[182] : 1'b0;
  assign N1084 = (N27)? address_i[53] : 
                 (N28)? address_i[117] : 
                 (N29)? address_i[181] : 1'b0;
  assign N1085 = (N27)? address_i[52] : 
                 (N28)? address_i[116] : 
                 (N29)? address_i[180] : 1'b0;
  assign N1086 = (N27)? address_i[51] : 
                 (N28)? address_i[115] : 
                 (N29)? address_i[179] : 1'b0;
  assign N1087 = (N27)? address_i[50] : 
                 (N28)? address_i[114] : 
                 (N29)? address_i[178] : 1'b0;
  assign N1088 = (N27)? address_i[49] : 
                 (N28)? address_i[113] : 
                 (N29)? address_i[177] : 1'b0;
  assign N1089 = (N27)? address_i[48] : 
                 (N28)? address_i[112] : 
                 (N29)? address_i[176] : 1'b0;
  assign N1090 = (N27)? address_i[47] : 
                 (N28)? address_i[111] : 
                 (N29)? address_i[175] : 1'b0;
  assign N1091 = (N27)? address_i[46] : 
                 (N28)? address_i[110] : 
                 (N29)? address_i[174] : 1'b0;
  assign N1092 = (N27)? address_i[45] : 
                 (N28)? address_i[109] : 
                 (N29)? address_i[173] : 1'b0;
  assign N1093 = (N27)? address_i[44] : 
                 (N28)? address_i[108] : 
                 (N29)? address_i[172] : 1'b0;
  assign N1094 = (N27)? address_i[43] : 
                 (N28)? address_i[107] : 
                 (N29)? address_i[171] : 1'b0;
  assign N1095 = (N27)? address_i[42] : 
                 (N28)? address_i[106] : 
                 (N29)? address_i[170] : 1'b0;
  assign N1096 = (N27)? address_i[41] : 
                 (N28)? address_i[105] : 
                 (N29)? address_i[169] : 1'b0;
  assign N1097 = (N27)? address_i[40] : 
                 (N28)? address_i[104] : 
                 (N29)? address_i[168] : 1'b0;
  assign N1098 = (N27)? address_i[39] : 
                 (N28)? address_i[103] : 
                 (N29)? address_i[167] : 1'b0;
  assign N1099 = (N27)? address_i[38] : 
                 (N28)? address_i[102] : 
                 (N29)? address_i[166] : 1'b0;
  assign N1100 = (N27)? address_i[37] : 
                 (N28)? address_i[101] : 
                 (N29)? address_i[165] : 1'b0;
  assign N1101 = (N27)? address_i[36] : 
                 (N28)? address_i[100] : 
                 (N29)? address_i[164] : 1'b0;
  assign N1102 = (N27)? address_i[35] : 
                 (N28)? address_i[99] : 
                 (N29)? address_i[163] : 1'b0;
  assign N1103 = (N27)? address_i[34] : 
                 (N28)? address_i[98] : 
                 (N29)? address_i[162] : 1'b0;
  assign N1104 = (N27)? address_i[33] : 
                 (N28)? address_i[97] : 
                 (N29)? address_i[161] : 1'b0;
  assign N1105 = (N27)? address_i[32] : 
                 (N28)? address_i[96] : 
                 (N29)? address_i[160] : 1'b0;
  assign N1106 = (N27)? address_i[31] : 
                 (N28)? address_i[95] : 
                 (N29)? address_i[159] : 1'b0;
  assign N1107 = (N27)? address_i[30] : 
                 (N28)? address_i[94] : 
                 (N29)? address_i[158] : 1'b0;
  assign N1108 = (N27)? address_i[29] : 
                 (N28)? address_i[93] : 
                 (N29)? address_i[157] : 1'b0;
  assign N1109 = (N27)? address_i[28] : 
                 (N28)? address_i[92] : 
                 (N29)? address_i[156] : 1'b0;
  assign N1110 = (N27)? address_i[27] : 
                 (N28)? address_i[91] : 
                 (N29)? address_i[155] : 1'b0;
  assign N1111 = (N27)? address_i[26] : 
                 (N28)? address_i[90] : 
                 (N29)? address_i[154] : 1'b0;
  assign N1112 = (N27)? address_i[25] : 
                 (N28)? address_i[89] : 
                 (N29)? address_i[153] : 1'b0;
  assign N1113 = (N27)? address_i[24] : 
                 (N28)? address_i[88] : 
                 (N29)? address_i[152] : 1'b0;
  assign N1114 = (N27)? address_i[23] : 
                 (N28)? address_i[87] : 
                 (N29)? address_i[151] : 1'b0;
  assign N1115 = (N27)? address_i[22] : 
                 (N28)? address_i[86] : 
                 (N29)? address_i[150] : 1'b0;
  assign N1116 = (N27)? address_i[21] : 
                 (N28)? address_i[85] : 
                 (N29)? address_i[149] : 1'b0;
  assign N1117 = (N27)? address_i[20] : 
                 (N28)? address_i[84] : 
                 (N29)? address_i[148] : 1'b0;
  assign N1118 = (N27)? address_i[19] : 
                 (N28)? address_i[83] : 
                 (N29)? address_i[147] : 1'b0;
  assign N1119 = (N27)? address_i[18] : 
                 (N28)? address_i[82] : 
                 (N29)? address_i[146] : 1'b0;
  assign N1120 = (N27)? address_i[17] : 
                 (N28)? address_i[81] : 
                 (N29)? address_i[145] : 1'b0;
  assign N1121 = (N27)? address_i[16] : 
                 (N28)? address_i[80] : 
                 (N29)? address_i[144] : 1'b0;
  assign N1122 = (N27)? address_i[15] : 
                 (N28)? address_i[79] : 
                 (N29)? address_i[143] : 1'b0;
  assign N1123 = (N27)? address_i[14] : 
                 (N28)? address_i[78] : 
                 (N29)? address_i[142] : 1'b0;
  assign N1124 = (N27)? address_i[13] : 
                 (N28)? address_i[77] : 
                 (N29)? address_i[141] : 1'b0;
  assign N1125 = (N27)? address_i[12] : 
                 (N28)? address_i[76] : 
                 (N29)? address_i[140] : 1'b0;
  assign N1126 = (N27)? address_i[11] : 
                 (N28)? address_i[75] : 
                 (N29)? address_i[139] : 1'b0;
  assign N1127 = (N27)? address_i[10] : 
                 (N28)? address_i[74] : 
                 (N29)? address_i[138] : 1'b0;
  assign N1128 = (N27)? address_i[9] : 
                 (N28)? address_i[73] : 
                 (N29)? address_i[137] : 1'b0;
  assign N1129 = (N27)? address_i[8] : 
                 (N28)? address_i[72] : 
                 (N29)? address_i[136] : 1'b0;
  assign N1130 = (N27)? address_i[7] : 
                 (N28)? address_i[71] : 
                 (N29)? address_i[135] : 1'b0;
  assign N1131 = (N27)? address_i[6] : 
                 (N28)? address_i[70] : 
                 (N29)? address_i[134] : 1'b0;
  assign N1132 = (N27)? address_i[5] : 
                 (N28)? address_i[69] : 
                 (N29)? address_i[133] : 1'b0;
  assign N1133 = (N27)? address_i[4] : 
                 (N28)? address_i[68] : 
                 (N29)? address_i[132] : 1'b0;
  assign N1134 = (N27)? address_i[3] : 
                 (N28)? address_i[67] : 
                 (N29)? address_i[131] : 1'b0;
  assign N1135 = (N27)? address_i[2] : 
                 (N28)? address_i[66] : 
                 (N29)? address_i[130] : 1'b0;
  assign N1136 = (N27)? address_i[1] : 
                 (N28)? address_i[65] : 
                 (N29)? address_i[129] : 1'b0;
  assign N1137 = (N27)? address_i[0] : 
                 (N28)? address_i[64] : 
                 (N29)? address_i[128] : 1'b0;
  assign N1139 = (N30)? data_wdata_i[63] : 
                 (N28)? data_wdata_i[127] : 
                 (N29)? data_wdata_i[191] : 1'b0;
  assign N30 = N1138;
  assign N1140 = (N30)? data_wdata_i[62] : 
                 (N28)? data_wdata_i[126] : 
                 (N29)? data_wdata_i[190] : 1'b0;
  assign N1141 = (N30)? data_wdata_i[61] : 
                 (N28)? data_wdata_i[125] : 
                 (N29)? data_wdata_i[189] : 1'b0;
  assign N1142 = (N30)? data_wdata_i[60] : 
                 (N28)? data_wdata_i[124] : 
                 (N29)? data_wdata_i[188] : 1'b0;
  assign N1143 = (N30)? data_wdata_i[59] : 
                 (N28)? data_wdata_i[123] : 
                 (N29)? data_wdata_i[187] : 1'b0;
  assign N1144 = (N30)? data_wdata_i[58] : 
                 (N28)? data_wdata_i[122] : 
                 (N29)? data_wdata_i[186] : 1'b0;
  assign N1145 = (N30)? data_wdata_i[57] : 
                 (N28)? data_wdata_i[121] : 
                 (N29)? data_wdata_i[185] : 1'b0;
  assign N1146 = (N30)? data_wdata_i[56] : 
                 (N28)? data_wdata_i[120] : 
                 (N29)? data_wdata_i[184] : 1'b0;
  assign N1147 = (N30)? data_wdata_i[55] : 
                 (N28)? data_wdata_i[119] : 
                 (N29)? data_wdata_i[183] : 1'b0;
  assign N1148 = (N30)? data_wdata_i[54] : 
                 (N28)? data_wdata_i[118] : 
                 (N29)? data_wdata_i[182] : 1'b0;
  assign N1149 = (N30)? data_wdata_i[53] : 
                 (N28)? data_wdata_i[117] : 
                 (N29)? data_wdata_i[181] : 1'b0;
  assign N1150 = (N30)? data_wdata_i[52] : 
                 (N28)? data_wdata_i[116] : 
                 (N29)? data_wdata_i[180] : 1'b0;
  assign N1151 = (N30)? data_wdata_i[51] : 
                 (N28)? data_wdata_i[115] : 
                 (N29)? data_wdata_i[179] : 1'b0;
  assign N1152 = (N30)? data_wdata_i[50] : 
                 (N28)? data_wdata_i[114] : 
                 (N29)? data_wdata_i[178] : 1'b0;
  assign N1153 = (N30)? data_wdata_i[49] : 
                 (N28)? data_wdata_i[113] : 
                 (N29)? data_wdata_i[177] : 1'b0;
  assign N1154 = (N30)? data_wdata_i[48] : 
                 (N28)? data_wdata_i[112] : 
                 (N29)? data_wdata_i[176] : 1'b0;
  assign N1155 = (N30)? data_wdata_i[47] : 
                 (N28)? data_wdata_i[111] : 
                 (N29)? data_wdata_i[175] : 1'b0;
  assign N1156 = (N30)? data_wdata_i[46] : 
                 (N28)? data_wdata_i[110] : 
                 (N29)? data_wdata_i[174] : 1'b0;
  assign N1157 = (N30)? data_wdata_i[45] : 
                 (N28)? data_wdata_i[109] : 
                 (N29)? data_wdata_i[173] : 1'b0;
  assign N1158 = (N30)? data_wdata_i[44] : 
                 (N28)? data_wdata_i[108] : 
                 (N29)? data_wdata_i[172] : 1'b0;
  assign N1159 = (N30)? data_wdata_i[43] : 
                 (N28)? data_wdata_i[107] : 
                 (N29)? data_wdata_i[171] : 1'b0;
  assign N1160 = (N30)? data_wdata_i[42] : 
                 (N28)? data_wdata_i[106] : 
                 (N29)? data_wdata_i[170] : 1'b0;
  assign N1161 = (N30)? data_wdata_i[41] : 
                 (N28)? data_wdata_i[105] : 
                 (N29)? data_wdata_i[169] : 1'b0;
  assign N1162 = (N30)? data_wdata_i[40] : 
                 (N28)? data_wdata_i[104] : 
                 (N29)? data_wdata_i[168] : 1'b0;
  assign N1163 = (N30)? data_wdata_i[39] : 
                 (N28)? data_wdata_i[103] : 
                 (N29)? data_wdata_i[167] : 1'b0;
  assign N1164 = (N30)? data_wdata_i[38] : 
                 (N28)? data_wdata_i[102] : 
                 (N29)? data_wdata_i[166] : 1'b0;
  assign N1165 = (N30)? data_wdata_i[37] : 
                 (N28)? data_wdata_i[101] : 
                 (N29)? data_wdata_i[165] : 1'b0;
  assign N1166 = (N30)? data_wdata_i[36] : 
                 (N28)? data_wdata_i[100] : 
                 (N29)? data_wdata_i[164] : 1'b0;
  assign N1167 = (N30)? data_wdata_i[35] : 
                 (N28)? data_wdata_i[99] : 
                 (N29)? data_wdata_i[163] : 1'b0;
  assign N1168 = (N30)? data_wdata_i[34] : 
                 (N28)? data_wdata_i[98] : 
                 (N29)? data_wdata_i[162] : 1'b0;
  assign N1169 = (N30)? data_wdata_i[33] : 
                 (N28)? data_wdata_i[97] : 
                 (N29)? data_wdata_i[161] : 1'b0;
  assign N1170 = (N30)? data_wdata_i[32] : 
                 (N28)? data_wdata_i[96] : 
                 (N29)? data_wdata_i[160] : 1'b0;
  assign N1171 = (N30)? data_wdata_i[31] : 
                 (N28)? data_wdata_i[95] : 
                 (N29)? data_wdata_i[159] : 1'b0;
  assign N1172 = (N30)? data_wdata_i[30] : 
                 (N28)? data_wdata_i[94] : 
                 (N29)? data_wdata_i[158] : 1'b0;
  assign N1173 = (N30)? data_wdata_i[29] : 
                 (N28)? data_wdata_i[93] : 
                 (N29)? data_wdata_i[157] : 1'b0;
  assign N1174 = (N30)? data_wdata_i[28] : 
                 (N28)? data_wdata_i[92] : 
                 (N29)? data_wdata_i[156] : 1'b0;
  assign N1175 = (N30)? data_wdata_i[27] : 
                 (N28)? data_wdata_i[91] : 
                 (N29)? data_wdata_i[155] : 1'b0;
  assign N1176 = (N30)? data_wdata_i[26] : 
                 (N28)? data_wdata_i[90] : 
                 (N29)? data_wdata_i[154] : 1'b0;
  assign N1177 = (N30)? data_wdata_i[25] : 
                 (N28)? data_wdata_i[89] : 
                 (N29)? data_wdata_i[153] : 1'b0;
  assign N1178 = (N30)? data_wdata_i[24] : 
                 (N28)? data_wdata_i[88] : 
                 (N29)? data_wdata_i[152] : 1'b0;
  assign N1179 = (N30)? data_wdata_i[23] : 
                 (N28)? data_wdata_i[87] : 
                 (N29)? data_wdata_i[151] : 1'b0;
  assign N1180 = (N30)? data_wdata_i[22] : 
                 (N28)? data_wdata_i[86] : 
                 (N29)? data_wdata_i[150] : 1'b0;
  assign N1181 = (N30)? data_wdata_i[21] : 
                 (N28)? data_wdata_i[85] : 
                 (N29)? data_wdata_i[149] : 1'b0;
  assign N1182 = (N30)? data_wdata_i[20] : 
                 (N28)? data_wdata_i[84] : 
                 (N29)? data_wdata_i[148] : 1'b0;
  assign N1183 = (N30)? data_wdata_i[19] : 
                 (N28)? data_wdata_i[83] : 
                 (N29)? data_wdata_i[147] : 1'b0;
  assign N1184 = (N30)? data_wdata_i[18] : 
                 (N28)? data_wdata_i[82] : 
                 (N29)? data_wdata_i[146] : 1'b0;
  assign N1185 = (N30)? data_wdata_i[17] : 
                 (N28)? data_wdata_i[81] : 
                 (N29)? data_wdata_i[145] : 1'b0;
  assign N1186 = (N30)? data_wdata_i[16] : 
                 (N28)? data_wdata_i[80] : 
                 (N29)? data_wdata_i[144] : 1'b0;
  assign N1187 = (N30)? data_wdata_i[15] : 
                 (N28)? data_wdata_i[79] : 
                 (N29)? data_wdata_i[143] : 1'b0;
  assign N1188 = (N30)? data_wdata_i[14] : 
                 (N28)? data_wdata_i[78] : 
                 (N29)? data_wdata_i[142] : 1'b0;
  assign N1189 = (N30)? data_wdata_i[13] : 
                 (N28)? data_wdata_i[77] : 
                 (N29)? data_wdata_i[141] : 1'b0;
  assign N1190 = (N30)? data_wdata_i[12] : 
                 (N28)? data_wdata_i[76] : 
                 (N29)? data_wdata_i[140] : 1'b0;
  assign N1191 = (N30)? data_wdata_i[11] : 
                 (N28)? data_wdata_i[75] : 
                 (N29)? data_wdata_i[139] : 1'b0;
  assign N1192 = (N30)? data_wdata_i[10] : 
                 (N28)? data_wdata_i[74] : 
                 (N29)? data_wdata_i[138] : 1'b0;
  assign N1193 = (N30)? data_wdata_i[9] : 
                 (N28)? data_wdata_i[73] : 
                 (N29)? data_wdata_i[137] : 1'b0;
  assign N1194 = (N30)? data_wdata_i[8] : 
                 (N28)? data_wdata_i[72] : 
                 (N29)? data_wdata_i[136] : 1'b0;
  assign N1195 = (N30)? data_wdata_i[7] : 
                 (N28)? data_wdata_i[71] : 
                 (N29)? data_wdata_i[135] : 1'b0;
  assign N1196 = (N30)? data_wdata_i[6] : 
                 (N28)? data_wdata_i[70] : 
                 (N29)? data_wdata_i[134] : 1'b0;
  assign N1197 = (N30)? data_wdata_i[5] : 
                 (N28)? data_wdata_i[69] : 
                 (N29)? data_wdata_i[133] : 1'b0;
  assign N1198 = (N30)? data_wdata_i[4] : 
                 (N28)? data_wdata_i[68] : 
                 (N29)? data_wdata_i[132] : 1'b0;
  assign N1199 = (N30)? data_wdata_i[3] : 
                 (N28)? data_wdata_i[67] : 
                 (N29)? data_wdata_i[131] : 1'b0;
  assign N1200 = (N30)? data_wdata_i[2] : 
                 (N28)? data_wdata_i[66] : 
                 (N29)? data_wdata_i[130] : 1'b0;
  assign N1201 = (N30)? data_wdata_i[1] : 
                 (N28)? data_wdata_i[65] : 
                 (N29)? data_wdata_i[129] : 1'b0;
  assign N1202 = (N30)? data_wdata_i[0] : 
                 (N28)? data_wdata_i[64] : 
                 (N29)? data_wdata_i[128] : 1'b0;
  assign N1203 = (N27)? data_be_i[7] : 
                 (N28)? data_be_i[15] : 
                 (N29)? data_be_i[23] : 1'b0;
  assign N1204 = (N27)? data_be_i[6] : 
                 (N28)? data_be_i[14] : 
                 (N29)? data_be_i[22] : 1'b0;
  assign N1205 = (N27)? data_be_i[5] : 
                 (N28)? data_be_i[13] : 
                 (N29)? data_be_i[21] : 1'b0;
  assign N1206 = (N27)? data_be_i[4] : 
                 (N28)? data_be_i[12] : 
                 (N29)? data_be_i[20] : 1'b0;
  assign N1207 = (N27)? data_be_i[3] : 
                 (N28)? data_be_i[11] : 
                 (N29)? data_be_i[19] : 1'b0;
  assign N1208 = (N27)? data_be_i[2] : 
                 (N28)? data_be_i[10] : 
                 (N29)? data_be_i[18] : 1'b0;
  assign N1209 = (N27)? data_be_i[1] : 
                 (N28)? data_be_i[9] : 
                 (N29)? data_be_i[17] : 1'b0;
  assign N1210 = (N27)? data_be_i[0] : 
                 (N28)? data_be_i[8] : 
                 (N29)? data_be_i[16] : 1'b0;
  assign N1211 = (N27)? data_size_i[1] : 
                 (N28)? data_size_i[3] : 
                 (N29)? data_size_i[5] : 1'b0;
  assign N1212 = (N27)? data_size_i[0] : 
                 (N28)? data_size_i[2] : 
                 (N29)? data_size_i[4] : 1'b0;
  assign N1215 = (N27)? data_we_i[0] : 
                 (N28)? data_we_i[1] : 
                 (N29)? data_we_i[2] : 1'b0;
  assign N34 = ~N31;
  assign N35 = ~N32;
  assign N36 = ~N33;
  assign N37 = ~state_q[1];
  assign N38 = ~state_q[0];
  assign N41 = ~N40;
  assign N42 = ~data_req_i[0];
  assign N188 = ~data_req_i[0];
  assign N189 = ~data_req_i[1];
  assign N336 = ~N335;
  assign N337 = ~data_req_i[2];
  assign N484 = ~N335;
  assign N1216 = ~data_rvalid_i;
  assign N1223 = ~rst_ni;
  assign N1224 = N41 | state_q[0];
  assign N1225 = ~N1224;
  assign N1226 = N41 | state_q[0];
  assign N1227 = ~N1226;
  assign N1228 = N1216 & N41;
  assign N1229 = N1228 | state_q[0];
  assign N1230 = ~N1229;

endmodule