module bsg_mux_one_hot_128_05
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [639:0] data_i;
  input [4:0] sel_one_hot_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383;
  wire [639:0] data_masked;
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[3];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[3];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[3];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[3];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[3];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[3];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[3];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[3];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[3];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[3];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[3];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[3];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[3];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[3];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[3];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[3];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[3];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[4];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[4];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[4];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[4];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[4];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[4];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[4];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[4];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[4];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[4];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[4];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[4];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[4];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[4];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[4];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[4];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[4];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[4];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[4];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[4];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[4];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[4];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[4];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[4];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[4];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[4];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[4];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[4];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[4];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[4];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[4];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[4];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[4];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[4];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[4];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[4];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[4];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[4];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[4];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[4];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[4];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[4];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[4];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[4];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[4];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[4];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[4];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[4];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[4];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[4];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[4];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[4];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[4];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[4];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[4];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[4];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[4];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[4];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[4];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[4];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[4];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[4];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[4];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[4];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[4];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[4];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[4];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[4];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[4];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[4];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[4];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[4];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[4];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[4];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[4];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[4];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[4];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[4];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[4];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[4];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[4];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[4];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[4];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[4];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[4];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[4];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[4];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[4];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[4];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[4];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[4];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[4];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[4];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[4];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[4];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[4];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[4];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[4];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[4];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[4];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[4];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[4];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[4];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[4];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[4];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[4];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[4];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[4];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[4];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[4];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[4];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[4];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[4];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[4];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[4];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[4];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[4];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[4];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[4];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[4];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[4];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[4];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[4];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[4];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[4];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[4];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[4];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[4];
  assign data_o[0] = N2 | data_masked[0];
  assign N2 = N1 | data_masked[128];
  assign N1 = N0 | data_masked[256];
  assign N0 = data_masked[512] | data_masked[384];
  assign data_o[1] = N5 | data_masked[1];
  assign N5 = N4 | data_masked[129];
  assign N4 = N3 | data_masked[257];
  assign N3 = data_masked[513] | data_masked[385];
  assign data_o[2] = N8 | data_masked[2];
  assign N8 = N7 | data_masked[130];
  assign N7 = N6 | data_masked[258];
  assign N6 = data_masked[514] | data_masked[386];
  assign data_o[3] = N11 | data_masked[3];
  assign N11 = N10 | data_masked[131];
  assign N10 = N9 | data_masked[259];
  assign N9 = data_masked[515] | data_masked[387];
  assign data_o[4] = N14 | data_masked[4];
  assign N14 = N13 | data_masked[132];
  assign N13 = N12 | data_masked[260];
  assign N12 = data_masked[516] | data_masked[388];
  assign data_o[5] = N17 | data_masked[5];
  assign N17 = N16 | data_masked[133];
  assign N16 = N15 | data_masked[261];
  assign N15 = data_masked[517] | data_masked[389];
  assign data_o[6] = N20 | data_masked[6];
  assign N20 = N19 | data_masked[134];
  assign N19 = N18 | data_masked[262];
  assign N18 = data_masked[518] | data_masked[390];
  assign data_o[7] = N23 | data_masked[7];
  assign N23 = N22 | data_masked[135];
  assign N22 = N21 | data_masked[263];
  assign N21 = data_masked[519] | data_masked[391];
  assign data_o[8] = N26 | data_masked[8];
  assign N26 = N25 | data_masked[136];
  assign N25 = N24 | data_masked[264];
  assign N24 = data_masked[520] | data_masked[392];
  assign data_o[9] = N29 | data_masked[9];
  assign N29 = N28 | data_masked[137];
  assign N28 = N27 | data_masked[265];
  assign N27 = data_masked[521] | data_masked[393];
  assign data_o[10] = N32 | data_masked[10];
  assign N32 = N31 | data_masked[138];
  assign N31 = N30 | data_masked[266];
  assign N30 = data_masked[522] | data_masked[394];
  assign data_o[11] = N35 | data_masked[11];
  assign N35 = N34 | data_masked[139];
  assign N34 = N33 | data_masked[267];
  assign N33 = data_masked[523] | data_masked[395];
  assign data_o[12] = N38 | data_masked[12];
  assign N38 = N37 | data_masked[140];
  assign N37 = N36 | data_masked[268];
  assign N36 = data_masked[524] | data_masked[396];
  assign data_o[13] = N41 | data_masked[13];
  assign N41 = N40 | data_masked[141];
  assign N40 = N39 | data_masked[269];
  assign N39 = data_masked[525] | data_masked[397];
  assign data_o[14] = N44 | data_masked[14];
  assign N44 = N43 | data_masked[142];
  assign N43 = N42 | data_masked[270];
  assign N42 = data_masked[526] | data_masked[398];
  assign data_o[15] = N47 | data_masked[15];
  assign N47 = N46 | data_masked[143];
  assign N46 = N45 | data_masked[271];
  assign N45 = data_masked[527] | data_masked[399];
  assign data_o[16] = N50 | data_masked[16];
  assign N50 = N49 | data_masked[144];
  assign N49 = N48 | data_masked[272];
  assign N48 = data_masked[528] | data_masked[400];
  assign data_o[17] = N53 | data_masked[17];
  assign N53 = N52 | data_masked[145];
  assign N52 = N51 | data_masked[273];
  assign N51 = data_masked[529] | data_masked[401];
  assign data_o[18] = N56 | data_masked[18];
  assign N56 = N55 | data_masked[146];
  assign N55 = N54 | data_masked[274];
  assign N54 = data_masked[530] | data_masked[402];
  assign data_o[19] = N59 | data_masked[19];
  assign N59 = N58 | data_masked[147];
  assign N58 = N57 | data_masked[275];
  assign N57 = data_masked[531] | data_masked[403];
  assign data_o[20] = N62 | data_masked[20];
  assign N62 = N61 | data_masked[148];
  assign N61 = N60 | data_masked[276];
  assign N60 = data_masked[532] | data_masked[404];
  assign data_o[21] = N65 | data_masked[21];
  assign N65 = N64 | data_masked[149];
  assign N64 = N63 | data_masked[277];
  assign N63 = data_masked[533] | data_masked[405];
  assign data_o[22] = N68 | data_masked[22];
  assign N68 = N67 | data_masked[150];
  assign N67 = N66 | data_masked[278];
  assign N66 = data_masked[534] | data_masked[406];
  assign data_o[23] = N71 | data_masked[23];
  assign N71 = N70 | data_masked[151];
  assign N70 = N69 | data_masked[279];
  assign N69 = data_masked[535] | data_masked[407];
  assign data_o[24] = N74 | data_masked[24];
  assign N74 = N73 | data_masked[152];
  assign N73 = N72 | data_masked[280];
  assign N72 = data_masked[536] | data_masked[408];
  assign data_o[25] = N77 | data_masked[25];
  assign N77 = N76 | data_masked[153];
  assign N76 = N75 | data_masked[281];
  assign N75 = data_masked[537] | data_masked[409];
  assign data_o[26] = N80 | data_masked[26];
  assign N80 = N79 | data_masked[154];
  assign N79 = N78 | data_masked[282];
  assign N78 = data_masked[538] | data_masked[410];
  assign data_o[27] = N83 | data_masked[27];
  assign N83 = N82 | data_masked[155];
  assign N82 = N81 | data_masked[283];
  assign N81 = data_masked[539] | data_masked[411];
  assign data_o[28] = N86 | data_masked[28];
  assign N86 = N85 | data_masked[156];
  assign N85 = N84 | data_masked[284];
  assign N84 = data_masked[540] | data_masked[412];
  assign data_o[29] = N89 | data_masked[29];
  assign N89 = N88 | data_masked[157];
  assign N88 = N87 | data_masked[285];
  assign N87 = data_masked[541] | data_masked[413];
  assign data_o[30] = N92 | data_masked[30];
  assign N92 = N91 | data_masked[158];
  assign N91 = N90 | data_masked[286];
  assign N90 = data_masked[542] | data_masked[414];
  assign data_o[31] = N95 | data_masked[31];
  assign N95 = N94 | data_masked[159];
  assign N94 = N93 | data_masked[287];
  assign N93 = data_masked[543] | data_masked[415];
  assign data_o[32] = N98 | data_masked[32];
  assign N98 = N97 | data_masked[160];
  assign N97 = N96 | data_masked[288];
  assign N96 = data_masked[544] | data_masked[416];
  assign data_o[33] = N101 | data_masked[33];
  assign N101 = N100 | data_masked[161];
  assign N100 = N99 | data_masked[289];
  assign N99 = data_masked[545] | data_masked[417];
  assign data_o[34] = N104 | data_masked[34];
  assign N104 = N103 | data_masked[162];
  assign N103 = N102 | data_masked[290];
  assign N102 = data_masked[546] | data_masked[418];
  assign data_o[35] = N107 | data_masked[35];
  assign N107 = N106 | data_masked[163];
  assign N106 = N105 | data_masked[291];
  assign N105 = data_masked[547] | data_masked[419];
  assign data_o[36] = N110 | data_masked[36];
  assign N110 = N109 | data_masked[164];
  assign N109 = N108 | data_masked[292];
  assign N108 = data_masked[548] | data_masked[420];
  assign data_o[37] = N113 | data_masked[37];
  assign N113 = N112 | data_masked[165];
  assign N112 = N111 | data_masked[293];
  assign N111 = data_masked[549] | data_masked[421];
  assign data_o[38] = N116 | data_masked[38];
  assign N116 = N115 | data_masked[166];
  assign N115 = N114 | data_masked[294];
  assign N114 = data_masked[550] | data_masked[422];
  assign data_o[39] = N119 | data_masked[39];
  assign N119 = N118 | data_masked[167];
  assign N118 = N117 | data_masked[295];
  assign N117 = data_masked[551] | data_masked[423];
  assign data_o[40] = N122 | data_masked[40];
  assign N122 = N121 | data_masked[168];
  assign N121 = N120 | data_masked[296];
  assign N120 = data_masked[552] | data_masked[424];
  assign data_o[41] = N125 | data_masked[41];
  assign N125 = N124 | data_masked[169];
  assign N124 = N123 | data_masked[297];
  assign N123 = data_masked[553] | data_masked[425];
  assign data_o[42] = N128 | data_masked[42];
  assign N128 = N127 | data_masked[170];
  assign N127 = N126 | data_masked[298];
  assign N126 = data_masked[554] | data_masked[426];
  assign data_o[43] = N131 | data_masked[43];
  assign N131 = N130 | data_masked[171];
  assign N130 = N129 | data_masked[299];
  assign N129 = data_masked[555] | data_masked[427];
  assign data_o[44] = N134 | data_masked[44];
  assign N134 = N133 | data_masked[172];
  assign N133 = N132 | data_masked[300];
  assign N132 = data_masked[556] | data_masked[428];
  assign data_o[45] = N137 | data_masked[45];
  assign N137 = N136 | data_masked[173];
  assign N136 = N135 | data_masked[301];
  assign N135 = data_masked[557] | data_masked[429];
  assign data_o[46] = N140 | data_masked[46];
  assign N140 = N139 | data_masked[174];
  assign N139 = N138 | data_masked[302];
  assign N138 = data_masked[558] | data_masked[430];
  assign data_o[47] = N143 | data_masked[47];
  assign N143 = N142 | data_masked[175];
  assign N142 = N141 | data_masked[303];
  assign N141 = data_masked[559] | data_masked[431];
  assign data_o[48] = N146 | data_masked[48];
  assign N146 = N145 | data_masked[176];
  assign N145 = N144 | data_masked[304];
  assign N144 = data_masked[560] | data_masked[432];
  assign data_o[49] = N149 | data_masked[49];
  assign N149 = N148 | data_masked[177];
  assign N148 = N147 | data_masked[305];
  assign N147 = data_masked[561] | data_masked[433];
  assign data_o[50] = N152 | data_masked[50];
  assign N152 = N151 | data_masked[178];
  assign N151 = N150 | data_masked[306];
  assign N150 = data_masked[562] | data_masked[434];
  assign data_o[51] = N155 | data_masked[51];
  assign N155 = N154 | data_masked[179];
  assign N154 = N153 | data_masked[307];
  assign N153 = data_masked[563] | data_masked[435];
  assign data_o[52] = N158 | data_masked[52];
  assign N158 = N157 | data_masked[180];
  assign N157 = N156 | data_masked[308];
  assign N156 = data_masked[564] | data_masked[436];
  assign data_o[53] = N161 | data_masked[53];
  assign N161 = N160 | data_masked[181];
  assign N160 = N159 | data_masked[309];
  assign N159 = data_masked[565] | data_masked[437];
  assign data_o[54] = N164 | data_masked[54];
  assign N164 = N163 | data_masked[182];
  assign N163 = N162 | data_masked[310];
  assign N162 = data_masked[566] | data_masked[438];
  assign data_o[55] = N167 | data_masked[55];
  assign N167 = N166 | data_masked[183];
  assign N166 = N165 | data_masked[311];
  assign N165 = data_masked[567] | data_masked[439];
  assign data_o[56] = N170 | data_masked[56];
  assign N170 = N169 | data_masked[184];
  assign N169 = N168 | data_masked[312];
  assign N168 = data_masked[568] | data_masked[440];
  assign data_o[57] = N173 | data_masked[57];
  assign N173 = N172 | data_masked[185];
  assign N172 = N171 | data_masked[313];
  assign N171 = data_masked[569] | data_masked[441];
  assign data_o[58] = N176 | data_masked[58];
  assign N176 = N175 | data_masked[186];
  assign N175 = N174 | data_masked[314];
  assign N174 = data_masked[570] | data_masked[442];
  assign data_o[59] = N179 | data_masked[59];
  assign N179 = N178 | data_masked[187];
  assign N178 = N177 | data_masked[315];
  assign N177 = data_masked[571] | data_masked[443];
  assign data_o[60] = N182 | data_masked[60];
  assign N182 = N181 | data_masked[188];
  assign N181 = N180 | data_masked[316];
  assign N180 = data_masked[572] | data_masked[444];
  assign data_o[61] = N185 | data_masked[61];
  assign N185 = N184 | data_masked[189];
  assign N184 = N183 | data_masked[317];
  assign N183 = data_masked[573] | data_masked[445];
  assign data_o[62] = N188 | data_masked[62];
  assign N188 = N187 | data_masked[190];
  assign N187 = N186 | data_masked[318];
  assign N186 = data_masked[574] | data_masked[446];
  assign data_o[63] = N191 | data_masked[63];
  assign N191 = N190 | data_masked[191];
  assign N190 = N189 | data_masked[319];
  assign N189 = data_masked[575] | data_masked[447];
  assign data_o[64] = N194 | data_masked[64];
  assign N194 = N193 | data_masked[192];
  assign N193 = N192 | data_masked[320];
  assign N192 = data_masked[576] | data_masked[448];
  assign data_o[65] = N197 | data_masked[65];
  assign N197 = N196 | data_masked[193];
  assign N196 = N195 | data_masked[321];
  assign N195 = data_masked[577] | data_masked[449];
  assign data_o[66] = N200 | data_masked[66];
  assign N200 = N199 | data_masked[194];
  assign N199 = N198 | data_masked[322];
  assign N198 = data_masked[578] | data_masked[450];
  assign data_o[67] = N203 | data_masked[67];
  assign N203 = N202 | data_masked[195];
  assign N202 = N201 | data_masked[323];
  assign N201 = data_masked[579] | data_masked[451];
  assign data_o[68] = N206 | data_masked[68];
  assign N206 = N205 | data_masked[196];
  assign N205 = N204 | data_masked[324];
  assign N204 = data_masked[580] | data_masked[452];
  assign data_o[69] = N209 | data_masked[69];
  assign N209 = N208 | data_masked[197];
  assign N208 = N207 | data_masked[325];
  assign N207 = data_masked[581] | data_masked[453];
  assign data_o[70] = N212 | data_masked[70];
  assign N212 = N211 | data_masked[198];
  assign N211 = N210 | data_masked[326];
  assign N210 = data_masked[582] | data_masked[454];
  assign data_o[71] = N215 | data_masked[71];
  assign N215 = N214 | data_masked[199];
  assign N214 = N213 | data_masked[327];
  assign N213 = data_masked[583] | data_masked[455];
  assign data_o[72] = N218 | data_masked[72];
  assign N218 = N217 | data_masked[200];
  assign N217 = N216 | data_masked[328];
  assign N216 = data_masked[584] | data_masked[456];
  assign data_o[73] = N221 | data_masked[73];
  assign N221 = N220 | data_masked[201];
  assign N220 = N219 | data_masked[329];
  assign N219 = data_masked[585] | data_masked[457];
  assign data_o[74] = N224 | data_masked[74];
  assign N224 = N223 | data_masked[202];
  assign N223 = N222 | data_masked[330];
  assign N222 = data_masked[586] | data_masked[458];
  assign data_o[75] = N227 | data_masked[75];
  assign N227 = N226 | data_masked[203];
  assign N226 = N225 | data_masked[331];
  assign N225 = data_masked[587] | data_masked[459];
  assign data_o[76] = N230 | data_masked[76];
  assign N230 = N229 | data_masked[204];
  assign N229 = N228 | data_masked[332];
  assign N228 = data_masked[588] | data_masked[460];
  assign data_o[77] = N233 | data_masked[77];
  assign N233 = N232 | data_masked[205];
  assign N232 = N231 | data_masked[333];
  assign N231 = data_masked[589] | data_masked[461];
  assign data_o[78] = N236 | data_masked[78];
  assign N236 = N235 | data_masked[206];
  assign N235 = N234 | data_masked[334];
  assign N234 = data_masked[590] | data_masked[462];
  assign data_o[79] = N239 | data_masked[79];
  assign N239 = N238 | data_masked[207];
  assign N238 = N237 | data_masked[335];
  assign N237 = data_masked[591] | data_masked[463];
  assign data_o[80] = N242 | data_masked[80];
  assign N242 = N241 | data_masked[208];
  assign N241 = N240 | data_masked[336];
  assign N240 = data_masked[592] | data_masked[464];
  assign data_o[81] = N245 | data_masked[81];
  assign N245 = N244 | data_masked[209];
  assign N244 = N243 | data_masked[337];
  assign N243 = data_masked[593] | data_masked[465];
  assign data_o[82] = N248 | data_masked[82];
  assign N248 = N247 | data_masked[210];
  assign N247 = N246 | data_masked[338];
  assign N246 = data_masked[594] | data_masked[466];
  assign data_o[83] = N251 | data_masked[83];
  assign N251 = N250 | data_masked[211];
  assign N250 = N249 | data_masked[339];
  assign N249 = data_masked[595] | data_masked[467];
  assign data_o[84] = N254 | data_masked[84];
  assign N254 = N253 | data_masked[212];
  assign N253 = N252 | data_masked[340];
  assign N252 = data_masked[596] | data_masked[468];
  assign data_o[85] = N257 | data_masked[85];
  assign N257 = N256 | data_masked[213];
  assign N256 = N255 | data_masked[341];
  assign N255 = data_masked[597] | data_masked[469];
  assign data_o[86] = N260 | data_masked[86];
  assign N260 = N259 | data_masked[214];
  assign N259 = N258 | data_masked[342];
  assign N258 = data_masked[598] | data_masked[470];
  assign data_o[87] = N263 | data_masked[87];
  assign N263 = N262 | data_masked[215];
  assign N262 = N261 | data_masked[343];
  assign N261 = data_masked[599] | data_masked[471];
  assign data_o[88] = N266 | data_masked[88];
  assign N266 = N265 | data_masked[216];
  assign N265 = N264 | data_masked[344];
  assign N264 = data_masked[600] | data_masked[472];
  assign data_o[89] = N269 | data_masked[89];
  assign N269 = N268 | data_masked[217];
  assign N268 = N267 | data_masked[345];
  assign N267 = data_masked[601] | data_masked[473];
  assign data_o[90] = N272 | data_masked[90];
  assign N272 = N271 | data_masked[218];
  assign N271 = N270 | data_masked[346];
  assign N270 = data_masked[602] | data_masked[474];
  assign data_o[91] = N275 | data_masked[91];
  assign N275 = N274 | data_masked[219];
  assign N274 = N273 | data_masked[347];
  assign N273 = data_masked[603] | data_masked[475];
  assign data_o[92] = N278 | data_masked[92];
  assign N278 = N277 | data_masked[220];
  assign N277 = N276 | data_masked[348];
  assign N276 = data_masked[604] | data_masked[476];
  assign data_o[93] = N281 | data_masked[93];
  assign N281 = N280 | data_masked[221];
  assign N280 = N279 | data_masked[349];
  assign N279 = data_masked[605] | data_masked[477];
  assign data_o[94] = N284 | data_masked[94];
  assign N284 = N283 | data_masked[222];
  assign N283 = N282 | data_masked[350];
  assign N282 = data_masked[606] | data_masked[478];
  assign data_o[95] = N287 | data_masked[95];
  assign N287 = N286 | data_masked[223];
  assign N286 = N285 | data_masked[351];
  assign N285 = data_masked[607] | data_masked[479];
  assign data_o[96] = N290 | data_masked[96];
  assign N290 = N289 | data_masked[224];
  assign N289 = N288 | data_masked[352];
  assign N288 = data_masked[608] | data_masked[480];
  assign data_o[97] = N293 | data_masked[97];
  assign N293 = N292 | data_masked[225];
  assign N292 = N291 | data_masked[353];
  assign N291 = data_masked[609] | data_masked[481];
  assign data_o[98] = N296 | data_masked[98];
  assign N296 = N295 | data_masked[226];
  assign N295 = N294 | data_masked[354];
  assign N294 = data_masked[610] | data_masked[482];
  assign data_o[99] = N299 | data_masked[99];
  assign N299 = N298 | data_masked[227];
  assign N298 = N297 | data_masked[355];
  assign N297 = data_masked[611] | data_masked[483];
  assign data_o[100] = N302 | data_masked[100];
  assign N302 = N301 | data_masked[228];
  assign N301 = N300 | data_masked[356];
  assign N300 = data_masked[612] | data_masked[484];
  assign data_o[101] = N305 | data_masked[101];
  assign N305 = N304 | data_masked[229];
  assign N304 = N303 | data_masked[357];
  assign N303 = data_masked[613] | data_masked[485];
  assign data_o[102] = N308 | data_masked[102];
  assign N308 = N307 | data_masked[230];
  assign N307 = N306 | data_masked[358];
  assign N306 = data_masked[614] | data_masked[486];
  assign data_o[103] = N311 | data_masked[103];
  assign N311 = N310 | data_masked[231];
  assign N310 = N309 | data_masked[359];
  assign N309 = data_masked[615] | data_masked[487];
  assign data_o[104] = N314 | data_masked[104];
  assign N314 = N313 | data_masked[232];
  assign N313 = N312 | data_masked[360];
  assign N312 = data_masked[616] | data_masked[488];
  assign data_o[105] = N317 | data_masked[105];
  assign N317 = N316 | data_masked[233];
  assign N316 = N315 | data_masked[361];
  assign N315 = data_masked[617] | data_masked[489];
  assign data_o[106] = N320 | data_masked[106];
  assign N320 = N319 | data_masked[234];
  assign N319 = N318 | data_masked[362];
  assign N318 = data_masked[618] | data_masked[490];
  assign data_o[107] = N323 | data_masked[107];
  assign N323 = N322 | data_masked[235];
  assign N322 = N321 | data_masked[363];
  assign N321 = data_masked[619] | data_masked[491];
  assign data_o[108] = N326 | data_masked[108];
  assign N326 = N325 | data_masked[236];
  assign N325 = N324 | data_masked[364];
  assign N324 = data_masked[620] | data_masked[492];
  assign data_o[109] = N329 | data_masked[109];
  assign N329 = N328 | data_masked[237];
  assign N328 = N327 | data_masked[365];
  assign N327 = data_masked[621] | data_masked[493];
  assign data_o[110] = N332 | data_masked[110];
  assign N332 = N331 | data_masked[238];
  assign N331 = N330 | data_masked[366];
  assign N330 = data_masked[622] | data_masked[494];
  assign data_o[111] = N335 | data_masked[111];
  assign N335 = N334 | data_masked[239];
  assign N334 = N333 | data_masked[367];
  assign N333 = data_masked[623] | data_masked[495];
  assign data_o[112] = N338 | data_masked[112];
  assign N338 = N337 | data_masked[240];
  assign N337 = N336 | data_masked[368];
  assign N336 = data_masked[624] | data_masked[496];
  assign data_o[113] = N341 | data_masked[113];
  assign N341 = N340 | data_masked[241];
  assign N340 = N339 | data_masked[369];
  assign N339 = data_masked[625] | data_masked[497];
  assign data_o[114] = N344 | data_masked[114];
  assign N344 = N343 | data_masked[242];
  assign N343 = N342 | data_masked[370];
  assign N342 = data_masked[626] | data_masked[498];
  assign data_o[115] = N347 | data_masked[115];
  assign N347 = N346 | data_masked[243];
  assign N346 = N345 | data_masked[371];
  assign N345 = data_masked[627] | data_masked[499];
  assign data_o[116] = N350 | data_masked[116];
  assign N350 = N349 | data_masked[244];
  assign N349 = N348 | data_masked[372];
  assign N348 = data_masked[628] | data_masked[500];
  assign data_o[117] = N353 | data_masked[117];
  assign N353 = N352 | data_masked[245];
  assign N352 = N351 | data_masked[373];
  assign N351 = data_masked[629] | data_masked[501];
  assign data_o[118] = N356 | data_masked[118];
  assign N356 = N355 | data_masked[246];
  assign N355 = N354 | data_masked[374];
  assign N354 = data_masked[630] | data_masked[502];
  assign data_o[119] = N359 | data_masked[119];
  assign N359 = N358 | data_masked[247];
  assign N358 = N357 | data_masked[375];
  assign N357 = data_masked[631] | data_masked[503];
  assign data_o[120] = N362 | data_masked[120];
  assign N362 = N361 | data_masked[248];
  assign N361 = N360 | data_masked[376];
  assign N360 = data_masked[632] | data_masked[504];
  assign data_o[121] = N365 | data_masked[121];
  assign N365 = N364 | data_masked[249];
  assign N364 = N363 | data_masked[377];
  assign N363 = data_masked[633] | data_masked[505];
  assign data_o[122] = N368 | data_masked[122];
  assign N368 = N367 | data_masked[250];
  assign N367 = N366 | data_masked[378];
  assign N366 = data_masked[634] | data_masked[506];
  assign data_o[123] = N371 | data_masked[123];
  assign N371 = N370 | data_masked[251];
  assign N370 = N369 | data_masked[379];
  assign N369 = data_masked[635] | data_masked[507];
  assign data_o[124] = N374 | data_masked[124];
  assign N374 = N373 | data_masked[252];
  assign N373 = N372 | data_masked[380];
  assign N372 = data_masked[636] | data_masked[508];
  assign data_o[125] = N377 | data_masked[125];
  assign N377 = N376 | data_masked[253];
  assign N376 = N375 | data_masked[381];
  assign N375 = data_masked[637] | data_masked[509];
  assign data_o[126] = N380 | data_masked[126];
  assign N380 = N379 | data_masked[254];
  assign N379 = N378 | data_masked[382];
  assign N378 = data_masked[638] | data_masked[510];
  assign data_o[127] = N383 | data_masked[127];
  assign N383 = N382 | data_masked[255];
  assign N382 = N381 | data_masked[383];
  assign N381 = data_masked[639] | data_masked[511];

endmodule