module control_3_bf8b4530d8d246dd74ac53a13471bba17941dff7(clk, rst, \complete_in.tag , \complete_in.valid , valid_in, repeated, flush_in, busy_in, deferred, sgl_pipe_in, stop_mark_in, gpr_write_valid_in, gpr_write_in, gpr_a_read_valid_in, gpr_a_read_in, gpr_b_read_valid_in, gpr_b_read_in, gpr_c_read_valid_in, gpr_c_read_in, \execute_next_tag.tag , \execute_next_tag.valid , \execute_next_cr_tag.tag , \execute_next_cr_tag.valid , cr_read_in, cr_write_in, valid_out, stall_out, stopped_out, gpr_bypass_a, gpr_bypass_b, gpr_bypass_c, cr_bypass, \instr_tag_out.tag , \instr_tag_out.valid );
  wire [9:0] _000_;
  wire [9:0] _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire [9:0] _012_;
  wire _013_;
  wire [7:0] _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire [9:0] _026_;
  wire _027_;
  wire [7:0] _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire [9:0] _040_;
  wire _041_;
  wire [7:0] _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire [9:0] _054_;
  wire _055_;
  wire [7:0] _056_;
  wire _057_;
  wire [1:0] _058_;
  wire [1:0] _059_;
  wire [1:0] _060_;
  reg [5:0] _061_ = 6'h00;
  reg [39:0] _062_;
  reg [1:0] _063_;
  reg [1:0] _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire [2:0] _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire [2:0] _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire [2:0] _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire [2:0] _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire [1:0] _089_;
  wire [1:0] _090_;
  wire [1:0] _091_;
  wire [1:0] _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire [2:0] _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire [2:0] _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire [2:0] _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire [2:0] _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire [1:0] _117_;
  wire [1:0] _118_;
  wire [1:0] _119_;
  wire [1:0] _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire [2:0] _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire [2:0] _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire [2:0] _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire [2:0] _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire [1:0] _145_;
  wire [1:0] _146_;
  wire [1:0] _147_;
  wire [1:0] _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire [31:0] _174_;
  wire [1:0] _175_;
  wire [1:0] _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire [31:0] _191_;
  wire [3:0] _192_;
  wire [3:0] _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire [5:0] _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire [1:0] _203_;
  wire _204_;
  wire _205_;
  wire [1:0] _206_;
  wire [1:0] _207_;
  wire _208_;
  wire [1:0] _209_;
  wire [1:0] _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire [1:0] _214_;
  wire [1:0] _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire [3:0] _219_;
  wire _220_;
  wire [1:0] _221_;
  wire _222_;
  wire _223_;
  wire [1:0] _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire [1:0] _228_;
  wire [1:0] _229_;
  wire _230_;
  wire _231_;
  wire [1:0] _232_;
  wire [3:0] _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire [31:0] _240_;
  wire [3:0] _241_;
  wire _242_;
  wire [9:0] _243_;
  input busy_in;
  wire busy_in;
  input clk;
  wire clk;
  input [1:0] \complete_in.tag ;
  wire [1:0] \complete_in.tag ;
  input \complete_in.valid ;
  wire \complete_in.valid ;
  output cr_bypass;
  wire cr_bypass;
  input cr_read_in;
  wire cr_read_in;
  wire cr_tag_stall;
  input cr_write_in;
  wire cr_write_in;
  wire cr_write_valid;
  wire [1:0] curr_cr_tag;
  wire [1:0] curr_tag;
  input deferred;
  wire deferred;
  input [1:0] \execute_next_cr_tag.tag ;
  wire [1:0] \execute_next_cr_tag.tag ;
  input \execute_next_cr_tag.valid ;
  wire \execute_next_cr_tag.valid ;
  input [1:0] \execute_next_tag.tag ;
  wire [1:0] \execute_next_tag.tag ;
  input \execute_next_tag.valid ;
  wire \execute_next_tag.valid ;
  input flush_in;
  wire flush_in;
  input [6:0] gpr_a_read_in;
  wire [6:0] gpr_a_read_in;
  input gpr_a_read_valid_in;
  wire gpr_a_read_valid_in;
  input [6:0] gpr_b_read_in;
  wire [6:0] gpr_b_read_in;
  input gpr_b_read_valid_in;
  wire gpr_b_read_valid_in;
  output gpr_bypass_a;
  wire gpr_bypass_a;
  output gpr_bypass_b;
  wire gpr_bypass_b;
  output gpr_bypass_c;
  wire gpr_bypass_c;
  input [6:0] gpr_c_read_in;
  wire [6:0] gpr_c_read_in;
  input gpr_c_read_valid_in;
  wire gpr_c_read_valid_in;
  wire gpr_tag_stall;
  input [6:0] gpr_write_in;
  wire [6:0] gpr_write_in;
  wire gpr_write_valid;
  input gpr_write_valid_in;
  wire gpr_write_valid_in;
  wire [2:0] instr_tag;
  output [1:0] \instr_tag_out.tag ;
  wire [1:0] \instr_tag_out.tag ;
  output \instr_tag_out.valid ;
  wire \instr_tag_out.valid ;
  wire [1:0] next_tag;
  wire [5:0] r_int;
  input repeated;
  wire repeated;
  wire [5:0] rin_int;
  input rst;
  wire rst;
  input sgl_pipe_in;
  wire sgl_pipe_in;
  output stall_out;
  wire stall_out;
  input stop_mark_in;
  wire stop_mark_in;
  output stopped_out;
  wire stopped_out;
  wire [39:0] tag_regs;
  input valid_in;
  wire valid_in;
  output valid_out;
  wire valid_out;
  assign _000_ = _176_[0] ? tag_regs[19:10] : tag_regs[9:0];
  assign _001_ = _176_[0] ? tag_regs[39:30] : tag_regs[29:20];
  assign _243_ = _176_[1] ? _001_ : _000_;
  assign _002_ = rst | flush_in;
  assign _003_ = 32'd0 == { 30'h00000000, \complete_in.tag  };
  assign _004_ = \complete_in.valid  & _003_;
  assign _005_ = _004_ ? 1'h0 : tag_regs[30];
  assign _006_ = _004_ ? 1'h0 : tag_regs[39];
  assign _007_ = tag_regs[37:31] == gpr_write_in;
  assign _008_ = gpr_write_valid & _007_;
  assign _009_ = _008_ ? 1'h0 : tag_regs[38];
  assign _010_ = 32'd0 == { 30'h00000000, instr_tag[1:0] };
  assign _011_ = instr_tag[2] & _010_;
  assign _012_ = _011_ ? { cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid } : { _006_, _009_, tag_regs[37:31], _005_ };
  assign _013_ = _002_ ? 1'h0 : _012_[0];
  assign _014_ = _002_ ? tag_regs[38:31] : _012_[8:1];
  assign _015_ = _002_ ? 1'h0 : _012_[9];
  assign _016_ = rst | flush_in;
  assign _017_ = 32'd1 == { 30'h00000000, \complete_in.tag  };
  assign _018_ = \complete_in.valid  & _017_;
  assign _019_ = _018_ ? 1'h0 : tag_regs[20];
  assign _020_ = _018_ ? 1'h0 : tag_regs[29];
  assign _021_ = tag_regs[27:21] == gpr_write_in;
  assign _022_ = gpr_write_valid & _021_;
  assign _023_ = _022_ ? 1'h0 : tag_regs[28];
  assign _024_ = 32'd1 == { 30'h00000000, instr_tag[1:0] };
  assign _025_ = instr_tag[2] & _024_;
  assign _026_ = _025_ ? { cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid } : { _020_, _023_, tag_regs[27:21], _019_ };
  assign _027_ = _016_ ? 1'h0 : _026_[0];
  assign _028_ = _016_ ? tag_regs[28:21] : _026_[8:1];
  assign _029_ = _016_ ? 1'h0 : _026_[9];
  assign _030_ = rst | flush_in;
  assign _031_ = 32'd2 == { 30'h00000000, \complete_in.tag  };
  assign _032_ = \complete_in.valid  & _031_;
  assign _033_ = _032_ ? 1'h0 : tag_regs[10];
  assign _034_ = _032_ ? 1'h0 : tag_regs[19];
  assign _035_ = tag_regs[17:11] == gpr_write_in;
  assign _036_ = gpr_write_valid & _035_;
  assign _037_ = _036_ ? 1'h0 : tag_regs[18];
  assign _038_ = 32'd2 == { 30'h00000000, instr_tag[1:0] };
  assign _039_ = instr_tag[2] & _038_;
  assign _040_ = _039_ ? { cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid } : { _034_, _037_, tag_regs[17:11], _033_ };
  assign _041_ = _030_ ? 1'h0 : _040_[0];
  assign _042_ = _030_ ? tag_regs[18:11] : _040_[8:1];
  assign _043_ = _030_ ? 1'h0 : _040_[9];
  assign _044_ = rst | flush_in;
  assign _045_ = 32'd3 == { 30'h00000000, \complete_in.tag  };
  assign _046_ = \complete_in.valid  & _045_;
  assign _047_ = _046_ ? 1'h0 : tag_regs[0];
  assign _048_ = _046_ ? 1'h0 : tag_regs[9];
  assign _049_ = tag_regs[7:1] == gpr_write_in;
  assign _050_ = gpr_write_valid & _049_;
  assign _051_ = _050_ ? 1'h0 : tag_regs[8];
  assign _052_ = 32'd3 == { 30'h00000000, instr_tag[1:0] };
  assign _053_ = instr_tag[2] & _052_;
  assign _054_ = _053_ ? { cr_write_valid, gpr_write_valid, gpr_write_in, gpr_write_valid } : { _048_, _051_, tag_regs[7:1], _047_ };
  assign _055_ = _044_ ? 1'h0 : _054_[0];
  assign _056_ = _044_ ? tag_regs[8:1] : _054_[8:1];
  assign _057_ = _044_ ? 1'h0 : _054_[9];
  assign _058_ = cr_write_valid ? instr_tag[1:0] : curr_cr_tag;
  assign _059_ = rst ? 2'h0 : next_tag;
  assign _060_ = rst ? 2'h0 : _058_;
  always @(posedge clk)
    _061_ <= rin_int;
  always @(posedge clk)
    _062_ <= { _015_, _014_, _013_, _029_, _028_, _027_, _043_, _042_, _041_, _057_, _056_, _055_ };
  always @(posedge clk)
    _063_ <= _059_;
  always @(posedge clk)
    _064_ <= _060_;
  assign _065_ = tag_regs[30] & tag_regs[38];
  assign _066_ = tag_regs[37:31] == gpr_a_read_in;
  assign _067_ = _065_ & _066_;
  assign _068_ = _067_ ? { gpr_a_read_valid_in, 2'h0 } : 3'h0;
  assign _069_ = tag_regs[20] & tag_regs[28];
  assign _070_ = tag_regs[27:21] == gpr_a_read_in;
  assign _071_ = _069_ & _070_;
  assign _072_ = _071_ ? { gpr_a_read_valid_in, 2'h1 } : _068_;
  assign _073_ = tag_regs[10] & tag_regs[18];
  assign _074_ = tag_regs[17:11] == gpr_a_read_in;
  assign _075_ = _073_ & _074_;
  assign _076_ = _075_ ? { gpr_a_read_valid_in, 2'h2 } : _072_;
  assign _077_ = tag_regs[0] & tag_regs[8];
  assign _078_ = tag_regs[7:1] == gpr_a_read_in;
  assign _079_ = _077_ & _078_;
  assign _080_ = _079_ ? { gpr_a_read_valid_in, 2'h3 } : _076_;
  assign _081_ = _080_[2] & \complete_in.valid ;
  assign _082_ = { 30'h00000000, _080_[1:0] } == { 30'h00000000, \complete_in.tag  };
  assign _083_ = _081_ & _082_;
  assign _084_ = _067_ ? gpr_a_read_valid_in : 1'h0;
  assign _085_ = _071_ ? gpr_a_read_valid_in : _084_;
  assign _086_ = _075_ ? gpr_a_read_valid_in : _085_;
  assign _087_ = _079_ ? gpr_a_read_valid_in : _086_;
  assign _088_ = _083_ ? 1'h0 : _087_;
  assign _089_ = _067_ ? 2'h0 : 2'h0;
  assign _090_ = _071_ ? 2'h1 : _089_;
  assign _091_ = _075_ ? 2'h2 : _090_;
  assign _092_ = _079_ ? 2'h3 : _091_;
  assign _093_ = tag_regs[30] & tag_regs[38];
  assign _094_ = tag_regs[37:31] == gpr_b_read_in;
  assign _095_ = _093_ & _094_;
  assign _096_ = _095_ ? { gpr_b_read_valid_in, 2'h0 } : 3'h0;
  assign _097_ = tag_regs[20] & tag_regs[28];
  assign _098_ = tag_regs[27:21] == gpr_b_read_in;
  assign _099_ = _097_ & _098_;
  assign _100_ = _099_ ? { gpr_b_read_valid_in, 2'h1 } : _096_;
  assign _101_ = tag_regs[10] & tag_regs[18];
  assign _102_ = tag_regs[17:11] == gpr_b_read_in;
  assign _103_ = _101_ & _102_;
  assign _104_ = _103_ ? { gpr_b_read_valid_in, 2'h2 } : _100_;
  assign _105_ = tag_regs[0] & tag_regs[8];
  assign _106_ = tag_regs[7:1] == gpr_b_read_in;
  assign _107_ = _105_ & _106_;
  assign _108_ = _107_ ? { gpr_b_read_valid_in, 2'h3 } : _104_;
  assign _109_ = _108_[2] & \complete_in.valid ;
  assign _110_ = { 30'h00000000, _108_[1:0] } == { 30'h00000000, \complete_in.tag  };
  assign _111_ = _109_ & _110_;
  assign _112_ = _095_ ? gpr_b_read_valid_in : 1'h0;
  assign _113_ = _099_ ? gpr_b_read_valid_in : _112_;
  assign _114_ = _103_ ? gpr_b_read_valid_in : _113_;
  assign _115_ = _107_ ? gpr_b_read_valid_in : _114_;
  assign _116_ = _111_ ? 1'h0 : _115_;
  assign _117_ = _095_ ? 2'h0 : 2'h0;
  assign _118_ = _099_ ? 2'h1 : _117_;
  assign _119_ = _103_ ? 2'h2 : _118_;
  assign _120_ = _107_ ? 2'h3 : _119_;
  assign _121_ = tag_regs[30] & tag_regs[38];
  assign _122_ = tag_regs[37:31] == gpr_c_read_in;
  assign _123_ = _121_ & _122_;
  assign _124_ = _123_ ? { gpr_c_read_valid_in, 2'h0 } : 3'h0;
  assign _125_ = tag_regs[20] & tag_regs[28];
  assign _126_ = tag_regs[27:21] == gpr_c_read_in;
  assign _127_ = _125_ & _126_;
  assign _128_ = _127_ ? { gpr_c_read_valid_in, 2'h1 } : _124_;
  assign _129_ = tag_regs[10] & tag_regs[18];
  assign _130_ = tag_regs[17:11] == gpr_c_read_in;
  assign _131_ = _129_ & _130_;
  assign _132_ = _131_ ? { gpr_c_read_valid_in, 2'h2 } : _128_;
  assign _133_ = tag_regs[0] & tag_regs[8];
  assign _134_ = tag_regs[7:1] == gpr_c_read_in;
  assign _135_ = _133_ & _134_;
  assign _136_ = _135_ ? { gpr_c_read_valid_in, 2'h3 } : _132_;
  assign _137_ = _136_[2] & \complete_in.valid ;
  assign _138_ = { 30'h00000000, _136_[1:0] } == { 30'h00000000, \complete_in.tag  };
  assign _139_ = _137_ & _138_;
  assign _140_ = _123_ ? gpr_c_read_valid_in : 1'h0;
  assign _141_ = _127_ ? gpr_c_read_valid_in : _140_;
  assign _142_ = _131_ ? gpr_c_read_valid_in : _141_;
  assign _143_ = _135_ ? gpr_c_read_valid_in : _142_;
  assign _144_ = _139_ ? 1'h0 : _143_;
  assign _145_ = _123_ ? 2'h0 : 2'h0;
  assign _146_ = _127_ ? 2'h1 : _145_;
  assign _147_ = _131_ ? 2'h2 : _146_;
  assign _148_ = _135_ ? 2'h3 : _147_;
  assign _149_ = \execute_next_tag.valid  & _088_;
  assign _150_ = { 30'h00000000, \execute_next_tag.tag  } == { 30'h00000000, _092_ };
  assign _151_ = _149_ & _150_;
  assign _152_ = 1'h1 & _151_;
  assign _153_ = _152_ ? 1'h1 : 1'h0;
  assign _154_ = \execute_next_tag.valid  & _116_;
  assign _155_ = { 30'h00000000, \execute_next_tag.tag  } == { 30'h00000000, _120_ };
  assign _156_ = _154_ & _155_;
  assign _157_ = 1'h1 & _156_;
  assign _158_ = _157_ ? 1'h1 : 1'h0;
  assign _159_ = \execute_next_tag.valid  & _144_;
  assign _160_ = { 30'h00000000, \execute_next_tag.tag  } == { 30'h00000000, _148_ };
  assign _161_ = _159_ & _160_;
  assign _162_ = 1'h1 & _161_;
  assign _163_ = _162_ ? 1'h1 : 1'h0;
  assign _164_ = ~ _153_;
  assign _165_ = _088_ & _164_;
  assign _166_ = ~ _158_;
  assign _167_ = _116_ & _166_;
  assign _168_ = _165_ | _167_;
  assign _169_ = ~ _163_;
  assign _170_ = _144_ & _169_;
  assign _171_ = _168_ | _170_;
  assign _172_ = ~ deferred;
  assign _173_ = _235_ & _172_;
  assign _174_ = { 30'h00000000, curr_tag } + 32'd1;
  assign _175_ = instr_tag[2] ? _174_[1:0] : curr_tag;
  assign _176_ = 2'h3 - curr_cr_tag;
  assign _177_ = cr_read_in & _243_[9];
  assign _178_ = _177_ & \complete_in.valid ;
  assign _179_ = { 30'h00000000, curr_cr_tag } == { 30'h00000000, \complete_in.tag  };
  assign _180_ = _178_ & _179_;
  assign _181_ = _180_ ? 1'h0 : _177_;
  assign _182_ = \execute_next_cr_tag.valid  & _181_;
  assign _183_ = { 30'h00000000, \execute_next_cr_tag.tag  } == { 30'h00000000, curr_cr_tag };
  assign _184_ = _182_ & _183_;
  assign _185_ = 1'h1 & _184_;
  assign _186_ = _185_ ? 1'h1 : 1'h0;
  assign _187_ = ~ _186_;
  assign _188_ = _181_ & _187_;
  assign _189_ = ~ flush_in;
  assign _190_ = valid_in & _189_;
  assign _191_ = { r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5:2] } - 32'd1;
  assign _192_ = \complete_in.valid  ? _191_[3:0] : r_int[5:2];
  assign _193_ = flush_in ? 4'h0 : _192_;
  assign _194_ = $signed({ r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5], r_int[5:2] }) >= $signed(32'd4);
  assign _195_ = _194_ ? 1'h0 : _190_;
  assign _196_ = _194_ ? 1'h1 : 1'h0;
  assign _197_ = rst ? 6'h00 : { _193_, r_int[1:0] };
  assign _198_ = rst ? 1'h0 : _195_;
  assign _199_ = { _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5:2] } == 32'd0;
  assign _200_ = stop_mark_in & _199_;
  assign _201_ = _200_ ? 1'h1 : 1'h0;
  assign _202_ = { _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5:2] } != 32'd0;
  assign _203_ = _202_ ? 2'h1 : 2'h2;
  assign _204_ = _202_ ? 1'h1 : _196_;
  assign _205_ = gpr_tag_stall | cr_tag_stall;
  assign _206_ = rst ? 2'h0 : r_int[1:0];
  assign _207_ = sgl_pipe_in ? _203_ : _206_;
  assign _208_ = sgl_pipe_in ? _204_ : _205_;
  assign _209_ = rst ? 2'h0 : r_int[1:0];
  assign _210_ = _198_ ? _207_ : _209_;
  assign _211_ = _198_ ? _208_ : _196_;
  assign _212_ = r_int[1:0] == 2'h0;
  assign _213_ = { _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5:2] } == 32'd0;
  assign _214_ = rst ? 2'h0 : r_int[1:0];
  assign _215_ = _213_ ? 2'h2 : _214_;
  assign _216_ = _213_ ? _196_ : 1'h1;
  assign _217_ = r_int[1:0] == 2'h1;
  assign _218_ = { _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5], _197_[5:2] } == 32'd0;
  assign _219_ = rst ? 4'h0 : _193_;
  assign _220_ = { _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_[3], _219_ } != 32'd0;
  assign _221_ = _220_ ? 2'h1 : 2'h2;
  assign _222_ = _220_ ? 1'h1 : _196_;
  assign _223_ = gpr_tag_stall | cr_tag_stall;
  assign _224_ = _226_ ? _221_ : 2'h0;
  assign _225_ = sgl_pipe_in ? _222_ : _223_;
  assign _226_ = _198_ & sgl_pipe_in;
  assign _227_ = _198_ ? _225_ : _196_;
  assign _228_ = rst ? 2'h0 : r_int[1:0];
  assign _229_ = _218_ ? _224_ : _228_;
  assign _230_ = _218_ ? _227_ : 1'h1;
  assign _231_ = r_int[1:0] == 2'h2;
  function [1:0] \27760 ;
    input [1:0] a;
    input [5:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \27760  = b[1:0];
      3'b?1?:
        \27760  = b[3:2];
      3'b1??:
        \27760  = b[5:4];
      default:
        \27760  = a;
    endcase
  endfunction
  assign _232_ = \27760 (2'hx, { _229_, _215_, _210_ }, { _231_, _217_, _212_ });
  assign _233_ = rst ? 4'h0 : _193_;
  function [0:0] \27765 ;
    input [0:0] a;
    input [2:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \27765  = b[0:0];
      3'b?1?:
        \27765  = b[1:1];
      3'b1??:
        \27765  = b[2:2];
      default:
        \27765  = a;
    endcase
  endfunction
  assign _234_ = \27765 (1'hx, { _230_, _216_, _211_ }, { _231_, _217_, _212_ });
  assign _235_ = _234_ ? 1'h0 : _198_;
  assign _236_ = gpr_write_valid_in & _235_;
  assign _237_ = cr_write_in & _235_;
  assign _238_ = ~ deferred;
  assign _239_ = _235_ & _238_;
  assign _240_ = { _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_[3], _233_ } + 32'd1;
  assign _241_ = _239_ ? _240_[3:0] : _233_;
  assign _242_ = _234_ | deferred;
  assign r_int = _061_;
  assign rin_int = { _241_, _232_ };
  assign gpr_write_valid = _236_;
  assign cr_write_valid = _237_;
  assign tag_regs = _062_;
  assign instr_tag = { _173_, curr_tag };
  assign gpr_tag_stall = _171_;
  assign cr_tag_stall = _188_;
  assign curr_tag = _063_;
  assign next_tag = _175_;
  assign curr_cr_tag = _064_;
  assign valid_out = _235_;
  assign stall_out = _242_;
  assign stopped_out = _201_;
  assign gpr_bypass_a = _153_;
  assign gpr_bypass_b = _158_;
  assign gpr_bypass_c = _163_;
  assign cr_bypass = _186_;
  assign \instr_tag_out.tag  = instr_tag[1:0];
  assign \instr_tag_out.valid  = instr_tag[2];
endmodule