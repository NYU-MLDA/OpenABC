module pipe_reg_simple_Depth1
(
  clk_i,
  rst_ni,
  d_i,
  d_o
);

  input [196:0] d_i;
  output [196:0] d_o;
  input clk_i;
  input rst_ni;
  wire N0;
  reg [196:0] d_o;

  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[196] <= 1'b0;
    end else if(1'b1) begin
      d_o[196] <= d_i[196];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[195] <= 1'b0;
    end else if(1'b1) begin
      d_o[195] <= d_i[195];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[194] <= 1'b0;
    end else if(1'b1) begin
      d_o[194] <= d_i[194];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[193] <= 1'b0;
    end else if(1'b1) begin
      d_o[193] <= d_i[193];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[192] <= 1'b0;
    end else if(1'b1) begin
      d_o[192] <= d_i[192];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[191] <= 1'b0;
    end else if(1'b1) begin
      d_o[191] <= d_i[191];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[190] <= 1'b0;
    end else if(1'b1) begin
      d_o[190] <= d_i[190];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[189] <= 1'b0;
    end else if(1'b1) begin
      d_o[189] <= d_i[189];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[188] <= 1'b0;
    end else if(1'b1) begin
      d_o[188] <= d_i[188];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[187] <= 1'b0;
    end else if(1'b1) begin
      d_o[187] <= d_i[187];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[186] <= 1'b0;
    end else if(1'b1) begin
      d_o[186] <= d_i[186];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[185] <= 1'b0;
    end else if(1'b1) begin
      d_o[185] <= d_i[185];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[184] <= 1'b0;
    end else if(1'b1) begin
      d_o[184] <= d_i[184];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[183] <= 1'b0;
    end else if(1'b1) begin
      d_o[183] <= d_i[183];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[182] <= 1'b0;
    end else if(1'b1) begin
      d_o[182] <= d_i[182];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[181] <= 1'b0;
    end else if(1'b1) begin
      d_o[181] <= d_i[181];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[180] <= 1'b0;
    end else if(1'b1) begin
      d_o[180] <= d_i[180];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[179] <= 1'b0;
    end else if(1'b1) begin
      d_o[179] <= d_i[179];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[178] <= 1'b0;
    end else if(1'b1) begin
      d_o[178] <= d_i[178];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[177] <= 1'b0;
    end else if(1'b1) begin
      d_o[177] <= d_i[177];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[176] <= 1'b0;
    end else if(1'b1) begin
      d_o[176] <= d_i[176];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[175] <= 1'b0;
    end else if(1'b1) begin
      d_o[175] <= d_i[175];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[174] <= 1'b0;
    end else if(1'b1) begin
      d_o[174] <= d_i[174];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[173] <= 1'b0;
    end else if(1'b1) begin
      d_o[173] <= d_i[173];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[172] <= 1'b0;
    end else if(1'b1) begin
      d_o[172] <= d_i[172];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[171] <= 1'b0;
    end else if(1'b1) begin
      d_o[171] <= d_i[171];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[170] <= 1'b0;
    end else if(1'b1) begin
      d_o[170] <= d_i[170];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[169] <= 1'b0;
    end else if(1'b1) begin
      d_o[169] <= d_i[169];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[168] <= 1'b0;
    end else if(1'b1) begin
      d_o[168] <= d_i[168];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[167] <= 1'b0;
    end else if(1'b1) begin
      d_o[167] <= d_i[167];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[166] <= 1'b0;
    end else if(1'b1) begin
      d_o[166] <= d_i[166];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[165] <= 1'b0;
    end else if(1'b1) begin
      d_o[165] <= d_i[165];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[164] <= 1'b0;
    end else if(1'b1) begin
      d_o[164] <= d_i[164];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[163] <= 1'b0;
    end else if(1'b1) begin
      d_o[163] <= d_i[163];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[162] <= 1'b0;
    end else if(1'b1) begin
      d_o[162] <= d_i[162];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[161] <= 1'b0;
    end else if(1'b1) begin
      d_o[161] <= d_i[161];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[160] <= 1'b0;
    end else if(1'b1) begin
      d_o[160] <= d_i[160];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[159] <= 1'b0;
    end else if(1'b1) begin
      d_o[159] <= d_i[159];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[158] <= 1'b0;
    end else if(1'b1) begin
      d_o[158] <= d_i[158];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[157] <= 1'b0;
    end else if(1'b1) begin
      d_o[157] <= d_i[157];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[156] <= 1'b0;
    end else if(1'b1) begin
      d_o[156] <= d_i[156];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[155] <= 1'b0;
    end else if(1'b1) begin
      d_o[155] <= d_i[155];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[154] <= 1'b0;
    end else if(1'b1) begin
      d_o[154] <= d_i[154];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[153] <= 1'b0;
    end else if(1'b1) begin
      d_o[153] <= d_i[153];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[152] <= 1'b0;
    end else if(1'b1) begin
      d_o[152] <= d_i[152];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[151] <= 1'b0;
    end else if(1'b1) begin
      d_o[151] <= d_i[151];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[150] <= 1'b0;
    end else if(1'b1) begin
      d_o[150] <= d_i[150];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[149] <= 1'b0;
    end else if(1'b1) begin
      d_o[149] <= d_i[149];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[148] <= 1'b0;
    end else if(1'b1) begin
      d_o[148] <= d_i[148];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[147] <= 1'b0;
    end else if(1'b1) begin
      d_o[147] <= d_i[147];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[146] <= 1'b0;
    end else if(1'b1) begin
      d_o[146] <= d_i[146];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[145] <= 1'b0;
    end else if(1'b1) begin
      d_o[145] <= d_i[145];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[144] <= 1'b0;
    end else if(1'b1) begin
      d_o[144] <= d_i[144];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[143] <= 1'b0;
    end else if(1'b1) begin
      d_o[143] <= d_i[143];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[142] <= 1'b0;
    end else if(1'b1) begin
      d_o[142] <= d_i[142];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[141] <= 1'b0;
    end else if(1'b1) begin
      d_o[141] <= d_i[141];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[140] <= 1'b0;
    end else if(1'b1) begin
      d_o[140] <= d_i[140];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[139] <= 1'b0;
    end else if(1'b1) begin
      d_o[139] <= d_i[139];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[138] <= 1'b0;
    end else if(1'b1) begin
      d_o[138] <= d_i[138];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[137] <= 1'b0;
    end else if(1'b1) begin
      d_o[137] <= d_i[137];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[136] <= 1'b0;
    end else if(1'b1) begin
      d_o[136] <= d_i[136];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[135] <= 1'b0;
    end else if(1'b1) begin
      d_o[135] <= d_i[135];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[134] <= 1'b0;
    end else if(1'b1) begin
      d_o[134] <= d_i[134];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[133] <= 1'b0;
    end else if(1'b1) begin
      d_o[133] <= d_i[133];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[132] <= 1'b0;
    end else if(1'b1) begin
      d_o[132] <= d_i[132];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[131] <= 1'b0;
    end else if(1'b1) begin
      d_o[131] <= d_i[131];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[130] <= 1'b0;
    end else if(1'b1) begin
      d_o[130] <= d_i[130];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[129] <= 1'b0;
    end else if(1'b1) begin
      d_o[129] <= d_i[129];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[128] <= 1'b0;
    end else if(1'b1) begin
      d_o[128] <= d_i[128];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[127] <= 1'b0;
    end else if(1'b1) begin
      d_o[127] <= d_i[127];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[126] <= 1'b0;
    end else if(1'b1) begin
      d_o[126] <= d_i[126];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[125] <= 1'b0;
    end else if(1'b1) begin
      d_o[125] <= d_i[125];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[124] <= 1'b0;
    end else if(1'b1) begin
      d_o[124] <= d_i[124];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[123] <= 1'b0;
    end else if(1'b1) begin
      d_o[123] <= d_i[123];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[122] <= 1'b0;
    end else if(1'b1) begin
      d_o[122] <= d_i[122];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[121] <= 1'b0;
    end else if(1'b1) begin
      d_o[121] <= d_i[121];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[120] <= 1'b0;
    end else if(1'b1) begin
      d_o[120] <= d_i[120];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[119] <= 1'b0;
    end else if(1'b1) begin
      d_o[119] <= d_i[119];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[118] <= 1'b0;
    end else if(1'b1) begin
      d_o[118] <= d_i[118];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[117] <= 1'b0;
    end else if(1'b1) begin
      d_o[117] <= d_i[117];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[116] <= 1'b0;
    end else if(1'b1) begin
      d_o[116] <= d_i[116];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[115] <= 1'b0;
    end else if(1'b1) begin
      d_o[115] <= d_i[115];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[114] <= 1'b0;
    end else if(1'b1) begin
      d_o[114] <= d_i[114];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[113] <= 1'b0;
    end else if(1'b1) begin
      d_o[113] <= d_i[113];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[112] <= 1'b0;
    end else if(1'b1) begin
      d_o[112] <= d_i[112];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[111] <= 1'b0;
    end else if(1'b1) begin
      d_o[111] <= d_i[111];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[110] <= 1'b0;
    end else if(1'b1) begin
      d_o[110] <= d_i[110];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[109] <= 1'b0;
    end else if(1'b1) begin
      d_o[109] <= d_i[109];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[108] <= 1'b0;
    end else if(1'b1) begin
      d_o[108] <= d_i[108];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[107] <= 1'b0;
    end else if(1'b1) begin
      d_o[107] <= d_i[107];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[106] <= 1'b0;
    end else if(1'b1) begin
      d_o[106] <= d_i[106];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[105] <= 1'b0;
    end else if(1'b1) begin
      d_o[105] <= d_i[105];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[104] <= 1'b0;
    end else if(1'b1) begin
      d_o[104] <= d_i[104];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[103] <= 1'b0;
    end else if(1'b1) begin
      d_o[103] <= d_i[103];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[102] <= 1'b0;
    end else if(1'b1) begin
      d_o[102] <= d_i[102];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[101] <= 1'b0;
    end else if(1'b1) begin
      d_o[101] <= d_i[101];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[100] <= 1'b0;
    end else if(1'b1) begin
      d_o[100] <= d_i[100];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[99] <= 1'b0;
    end else if(1'b1) begin
      d_o[99] <= d_i[99];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[98] <= 1'b0;
    end else if(1'b1) begin
      d_o[98] <= d_i[98];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[97] <= 1'b0;
    end else if(1'b1) begin
      d_o[97] <= d_i[97];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[96] <= 1'b0;
    end else if(1'b1) begin
      d_o[96] <= d_i[96];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[95] <= 1'b0;
    end else if(1'b1) begin
      d_o[95] <= d_i[95];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[94] <= 1'b0;
    end else if(1'b1) begin
      d_o[94] <= d_i[94];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[93] <= 1'b0;
    end else if(1'b1) begin
      d_o[93] <= d_i[93];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[92] <= 1'b0;
    end else if(1'b1) begin
      d_o[92] <= d_i[92];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[91] <= 1'b0;
    end else if(1'b1) begin
      d_o[91] <= d_i[91];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[90] <= 1'b0;
    end else if(1'b1) begin
      d_o[90] <= d_i[90];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[89] <= 1'b0;
    end else if(1'b1) begin
      d_o[89] <= d_i[89];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[88] <= 1'b0;
    end else if(1'b1) begin
      d_o[88] <= d_i[88];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[87] <= 1'b0;
    end else if(1'b1) begin
      d_o[87] <= d_i[87];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[86] <= 1'b0;
    end else if(1'b1) begin
      d_o[86] <= d_i[86];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[85] <= 1'b0;
    end else if(1'b1) begin
      d_o[85] <= d_i[85];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[84] <= 1'b0;
    end else if(1'b1) begin
      d_o[84] <= d_i[84];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[83] <= 1'b0;
    end else if(1'b1) begin
      d_o[83] <= d_i[83];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[82] <= 1'b0;
    end else if(1'b1) begin
      d_o[82] <= d_i[82];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[81] <= 1'b0;
    end else if(1'b1) begin
      d_o[81] <= d_i[81];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[80] <= 1'b0;
    end else if(1'b1) begin
      d_o[80] <= d_i[80];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[79] <= 1'b0;
    end else if(1'b1) begin
      d_o[79] <= d_i[79];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[78] <= 1'b0;
    end else if(1'b1) begin
      d_o[78] <= d_i[78];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[77] <= 1'b0;
    end else if(1'b1) begin
      d_o[77] <= d_i[77];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[76] <= 1'b0;
    end else if(1'b1) begin
      d_o[76] <= d_i[76];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[75] <= 1'b0;
    end else if(1'b1) begin
      d_o[75] <= d_i[75];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[74] <= 1'b0;
    end else if(1'b1) begin
      d_o[74] <= d_i[74];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[73] <= 1'b0;
    end else if(1'b1) begin
      d_o[73] <= d_i[73];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[72] <= 1'b0;
    end else if(1'b1) begin
      d_o[72] <= d_i[72];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[71] <= 1'b0;
    end else if(1'b1) begin
      d_o[71] <= d_i[71];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[70] <= 1'b0;
    end else if(1'b1) begin
      d_o[70] <= d_i[70];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[69] <= 1'b0;
    end else if(1'b1) begin
      d_o[69] <= d_i[69];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[68] <= 1'b0;
    end else if(1'b1) begin
      d_o[68] <= d_i[68];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[67] <= 1'b0;
    end else if(1'b1) begin
      d_o[67] <= d_i[67];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[66] <= 1'b0;
    end else if(1'b1) begin
      d_o[66] <= d_i[66];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[65] <= 1'b0;
    end else if(1'b1) begin
      d_o[65] <= d_i[65];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[64] <= 1'b0;
    end else if(1'b1) begin
      d_o[64] <= d_i[64];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[63] <= 1'b0;
    end else if(1'b1) begin
      d_o[63] <= d_i[63];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[62] <= 1'b0;
    end else if(1'b1) begin
      d_o[62] <= d_i[62];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[61] <= 1'b0;
    end else if(1'b1) begin
      d_o[61] <= d_i[61];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[60] <= 1'b0;
    end else if(1'b1) begin
      d_o[60] <= d_i[60];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[59] <= 1'b0;
    end else if(1'b1) begin
      d_o[59] <= d_i[59];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[58] <= 1'b0;
    end else if(1'b1) begin
      d_o[58] <= d_i[58];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[57] <= 1'b0;
    end else if(1'b1) begin
      d_o[57] <= d_i[57];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[56] <= 1'b0;
    end else if(1'b1) begin
      d_o[56] <= d_i[56];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[55] <= 1'b0;
    end else if(1'b1) begin
      d_o[55] <= d_i[55];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[54] <= 1'b0;
    end else if(1'b1) begin
      d_o[54] <= d_i[54];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[53] <= 1'b0;
    end else if(1'b1) begin
      d_o[53] <= d_i[53];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[52] <= 1'b0;
    end else if(1'b1) begin
      d_o[52] <= d_i[52];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[51] <= 1'b0;
    end else if(1'b1) begin
      d_o[51] <= d_i[51];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[50] <= 1'b0;
    end else if(1'b1) begin
      d_o[50] <= d_i[50];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[49] <= 1'b0;
    end else if(1'b1) begin
      d_o[49] <= d_i[49];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[48] <= 1'b0;
    end else if(1'b1) begin
      d_o[48] <= d_i[48];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[47] <= 1'b0;
    end else if(1'b1) begin
      d_o[47] <= d_i[47];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[46] <= 1'b0;
    end else if(1'b1) begin
      d_o[46] <= d_i[46];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[45] <= 1'b0;
    end else if(1'b1) begin
      d_o[45] <= d_i[45];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[44] <= 1'b0;
    end else if(1'b1) begin
      d_o[44] <= d_i[44];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[43] <= 1'b0;
    end else if(1'b1) begin
      d_o[43] <= d_i[43];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[42] <= 1'b0;
    end else if(1'b1) begin
      d_o[42] <= d_i[42];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[41] <= 1'b0;
    end else if(1'b1) begin
      d_o[41] <= d_i[41];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[40] <= 1'b0;
    end else if(1'b1) begin
      d_o[40] <= d_i[40];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[39] <= 1'b0;
    end else if(1'b1) begin
      d_o[39] <= d_i[39];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[38] <= 1'b0;
    end else if(1'b1) begin
      d_o[38] <= d_i[38];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[37] <= 1'b0;
    end else if(1'b1) begin
      d_o[37] <= d_i[37];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[36] <= 1'b0;
    end else if(1'b1) begin
      d_o[36] <= d_i[36];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[35] <= 1'b0;
    end else if(1'b1) begin
      d_o[35] <= d_i[35];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[34] <= 1'b0;
    end else if(1'b1) begin
      d_o[34] <= d_i[34];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[33] <= 1'b0;
    end else if(1'b1) begin
      d_o[33] <= d_i[33];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[32] <= 1'b0;
    end else if(1'b1) begin
      d_o[32] <= d_i[32];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[31] <= 1'b0;
    end else if(1'b1) begin
      d_o[31] <= d_i[31];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[30] <= 1'b0;
    end else if(1'b1) begin
      d_o[30] <= d_i[30];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[29] <= 1'b0;
    end else if(1'b1) begin
      d_o[29] <= d_i[29];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[28] <= 1'b0;
    end else if(1'b1) begin
      d_o[28] <= d_i[28];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[27] <= 1'b0;
    end else if(1'b1) begin
      d_o[27] <= d_i[27];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[26] <= 1'b0;
    end else if(1'b1) begin
      d_o[26] <= d_i[26];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[25] <= 1'b0;
    end else if(1'b1) begin
      d_o[25] <= d_i[25];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[24] <= 1'b0;
    end else if(1'b1) begin
      d_o[24] <= d_i[24];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[23] <= 1'b0;
    end else if(1'b1) begin
      d_o[23] <= d_i[23];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[22] <= 1'b0;
    end else if(1'b1) begin
      d_o[22] <= d_i[22];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[21] <= 1'b0;
    end else if(1'b1) begin
      d_o[21] <= d_i[21];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[20] <= 1'b0;
    end else if(1'b1) begin
      d_o[20] <= d_i[20];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[19] <= 1'b0;
    end else if(1'b1) begin
      d_o[19] <= d_i[19];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[18] <= 1'b0;
    end else if(1'b1) begin
      d_o[18] <= d_i[18];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[17] <= 1'b0;
    end else if(1'b1) begin
      d_o[17] <= d_i[17];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[16] <= 1'b0;
    end else if(1'b1) begin
      d_o[16] <= d_i[16];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[15] <= 1'b0;
    end else if(1'b1) begin
      d_o[15] <= d_i[15];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[14] <= 1'b0;
    end else if(1'b1) begin
      d_o[14] <= d_i[14];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[13] <= 1'b0;
    end else if(1'b1) begin
      d_o[13] <= d_i[13];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[12] <= 1'b0;
    end else if(1'b1) begin
      d_o[12] <= d_i[12];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[11] <= 1'b0;
    end else if(1'b1) begin
      d_o[11] <= d_i[11];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[10] <= 1'b0;
    end else if(1'b1) begin
      d_o[10] <= d_i[10];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[9] <= 1'b0;
    end else if(1'b1) begin
      d_o[9] <= d_i[9];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[8] <= 1'b0;
    end else if(1'b1) begin
      d_o[8] <= d_i[8];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[7] <= 1'b0;
    end else if(1'b1) begin
      d_o[7] <= d_i[7];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[6] <= 1'b0;
    end else if(1'b1) begin
      d_o[6] <= d_i[6];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[5] <= 1'b0;
    end else if(1'b1) begin
      d_o[5] <= d_i[5];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[4] <= 1'b0;
    end else if(1'b1) begin
      d_o[4] <= d_i[4];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[3] <= 1'b0;
    end else if(1'b1) begin
      d_o[3] <= d_i[3];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[2] <= 1'b0;
    end else if(1'b1) begin
      d_o[2] <= d_i[2];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[1] <= 1'b0;
    end else if(1'b1) begin
      d_o[1] <= d_i[1];
    end 
  end


  always @(posedge clk_i or posedge N0) begin
    if(N0) begin
      d_o[0] <= 1'b0;
    end else if(1'b1) begin
      d_o[0] <= d_i[0];
    end 
  end

  assign N0 = ~rst_ni;

endmodule