module bp_cce_msg_uncached_05
(
  clk_i,
  reset_i,
  cce_id_i,
  lce_req_i,
  lce_req_v_i,
  lce_req_yumi_o,
  lce_cmd_o,
  lce_cmd_v_o,
  lce_cmd_ready_i,
  mem_resp_i,
  mem_resp_v_i,
  mem_resp_yumi_o,
  mem_cmd_o,
  mem_cmd_v_o,
  mem_cmd_ready_i
);

  input [3:0] cce_id_i;
  input [118:0] lce_req_i;
  output [567:0] lce_cmd_o;
  input [571:0] mem_resp_i;
  output [571:0] mem_cmd_o;
  input clk_i;
  input reset_i;
  input lce_req_v_i;
  input lce_cmd_ready_i;
  input mem_resp_v_i;
  input mem_cmd_ready_i;
  output lce_req_yumi_o;
  output lce_cmd_v_o;
  output mem_resp_yumi_o;
  output mem_cmd_v_o;
  wire [567:0] lce_cmd_o;
  wire [571:0] mem_cmd_o;
  wire lce_req_yumi_o,lce_cmd_v_o,mem_resp_yumi_o,mem_cmd_v_o,N0,N1,N2,N3,N4,N5,N6,N7,
  N8,N9,N10,N11,N12,N13,lce_req_r_msg__65_,lce_req_r_msg__64_,lce_req_r_msg__63_,
  lce_req_r_msg__62_,lce_req_r_msg__61_,lce_req_r_msg__60_,lce_req_r_msg__59_,
  lce_req_r_msg__58_,lce_req_r_msg__57_,lce_req_r_msg__56_,lce_req_r_msg__55_,
  lce_req_r_msg__54_,lce_req_r_msg__53_,lce_req_r_msg__52_,lce_req_r_msg__51_,
  lce_req_r_msg__50_,lce_req_r_msg__49_,lce_req_r_msg__48_,lce_req_r_msg__47_,
  lce_req_r_msg__46_,lce_req_r_msg__45_,lce_req_r_msg__44_,lce_req_r_msg__43_,lce_req_r_msg__42_,
  lce_req_r_msg__41_,lce_req_r_msg__40_,lce_req_r_msg__39_,lce_req_r_msg__38_,
  lce_req_r_msg__37_,lce_req_r_msg__36_,lce_req_r_msg__35_,lce_req_r_msg__34_,
  lce_req_r_msg__33_,lce_req_r_msg__32_,lce_req_r_msg__31_,lce_req_r_msg__30_,
  lce_req_r_msg__29_,lce_req_r_msg__28_,lce_req_r_msg__27_,lce_req_r_msg__26_,lce_req_r_msg__25_,
  lce_req_r_msg__24_,lce_req_r_msg__23_,lce_req_r_msg__22_,lce_req_r_msg__21_,
  lce_req_r_msg__20_,lce_req_r_msg__19_,lce_req_r_msg__18_,lce_req_r_msg__17_,
  lce_req_r_msg__16_,lce_req_r_msg__15_,lce_req_r_msg__14_,lce_req_r_msg__13_,
  lce_req_r_msg__12_,lce_req_r_msg__11_,lce_req_r_msg__10_,lce_req_r_msg__9_,
  lce_req_r_msg__8_,lce_req_r_msg__7_,lce_req_r_msg__6_,lce_req_r_msg__5_,lce_req_r_msg__4_,
  lce_req_r_msg__3_,lce_req_r_msg__2_,lce_req_r_msg__1_,lce_req_r_msg__0_,
  lce_req_r_addr__39_,lce_req_r_addr__38_,lce_req_r_addr__37_,lce_req_r_addr__36_,
  lce_req_r_addr__35_,lce_req_r_addr__34_,lce_req_r_addr__33_,lce_req_r_addr__32_,
  lce_req_r_addr__31_,lce_req_r_addr__30_,lce_req_r_addr__29_,lce_req_r_addr__28_,
  lce_req_r_addr__27_,lce_req_r_addr__26_,lce_req_r_addr__25_,lce_req_r_addr__24_,
  lce_req_r_addr__23_,lce_req_r_addr__22_,lce_req_r_addr__21_,lce_req_r_addr__20_,
  lce_req_r_addr__19_,lce_req_r_addr__18_,lce_req_r_addr__17_,lce_req_r_addr__16_,
  lce_req_r_addr__15_,lce_req_r_addr__14_,lce_req_r_addr__13_,lce_req_r_addr__12_,
  lce_req_r_addr__11_,lce_req_r_addr__10_,lce_req_r_addr__9_,lce_req_r_addr__8_,
  lce_req_r_addr__7_,lce_req_r_addr__6_,lce_req_r_addr__5_,lce_req_r_addr__4_,lce_req_r_addr__3_,
  lce_req_r_addr__2_,lce_req_r_addr__1_,lce_req_r_addr__0_,lce_req_r_src_id__5_,
  lce_req_r_src_id__4_,lce_req_r_src_id__3_,lce_req_r_src_id__2_,lce_req_r_src_id__1_,
  lce_req_r_src_id__0_,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,
  N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,
  N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,
  N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,
  N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,
  N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,
  N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,
  N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,
  N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,
  N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,
  N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,
  N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,
  N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,
  N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,
  N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,
  N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,
  N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,
  N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,
  N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,
  N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,
  N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,
  N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,
  N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,
  N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,
  N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,
  N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,
  N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,
  N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,
  N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,
  N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,
  N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,
  N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,
  N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,
  N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,
  N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,
  N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,
  N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,
  N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,
  N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,
  N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,
  N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,
  N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,
  N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,
  N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,
  N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,
  N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,
  N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,
  N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,
  N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,
  N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,
  N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,
  N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,
  N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,
  N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,
  N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,
  N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,
  N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,
  N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,
  N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,
  N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,
  N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,
  N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,
  N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,
  N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,
  N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,
  N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,
  N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,
  N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,
  N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,
  N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,
  N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,
  N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,
  N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,
  N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,
  N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,
  N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,
  N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,
  N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,
  N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,
  N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,
  N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,
  N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,
  N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,
  N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,
  N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,
  N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,
  N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,
  N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,
  N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,
  N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,
  N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,
  N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,
  N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,
  N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,
  N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,
  N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,
  N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,
  N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,
  N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,
  N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,
  N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,
  N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
  N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,
  N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
  N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,
  N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,
  N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,
  N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,
  N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,
  N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,
  N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,
  N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,
  N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,
  N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,
  N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,
  N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743;
  wire [1:0] uc_state,uc_state_n;
  reg lce_req_r_msg__65__sv2v_reg,lce_req_r_msg__64__sv2v_reg,
  lce_req_r_msg__63__sv2v_reg,lce_req_r_msg__62__sv2v_reg,lce_req_r_msg__61__sv2v_reg,
  lce_req_r_msg__60__sv2v_reg,lce_req_r_msg__59__sv2v_reg,lce_req_r_msg__58__sv2v_reg,
  lce_req_r_msg__57__sv2v_reg,lce_req_r_msg__56__sv2v_reg,lce_req_r_msg__55__sv2v_reg,
  lce_req_r_msg__54__sv2v_reg,lce_req_r_msg__53__sv2v_reg,lce_req_r_msg__52__sv2v_reg,
  lce_req_r_msg__51__sv2v_reg,lce_req_r_msg__50__sv2v_reg,lce_req_r_msg__49__sv2v_reg,
  lce_req_r_msg__48__sv2v_reg,lce_req_r_msg__47__sv2v_reg,lce_req_r_msg__46__sv2v_reg,
  lce_req_r_msg__45__sv2v_reg,lce_req_r_msg__44__sv2v_reg,
  lce_req_r_msg__43__sv2v_reg,lce_req_r_msg__42__sv2v_reg,lce_req_r_msg__41__sv2v_reg,
  lce_req_r_msg__40__sv2v_reg,lce_req_r_msg__39__sv2v_reg,lce_req_r_msg__38__sv2v_reg,
  lce_req_r_msg__37__sv2v_reg,lce_req_r_msg__36__sv2v_reg,lce_req_r_msg__35__sv2v_reg,
  lce_req_r_msg__34__sv2v_reg,lce_req_r_msg__33__sv2v_reg,lce_req_r_msg__32__sv2v_reg,
  lce_req_r_msg__31__sv2v_reg,lce_req_r_msg__30__sv2v_reg,lce_req_r_msg__29__sv2v_reg,
  lce_req_r_msg__28__sv2v_reg,lce_req_r_msg__27__sv2v_reg,lce_req_r_msg__26__sv2v_reg,
  lce_req_r_msg__25__sv2v_reg,lce_req_r_msg__24__sv2v_reg,
  lce_req_r_msg__23__sv2v_reg,lce_req_r_msg__22__sv2v_reg,lce_req_r_msg__21__sv2v_reg,
  lce_req_r_msg__20__sv2v_reg,lce_req_r_msg__19__sv2v_reg,lce_req_r_msg__18__sv2v_reg,
  lce_req_r_msg__17__sv2v_reg,lce_req_r_msg__16__sv2v_reg,lce_req_r_msg__15__sv2v_reg,
  lce_req_r_msg__14__sv2v_reg,lce_req_r_msg__13__sv2v_reg,lce_req_r_msg__12__sv2v_reg,
  lce_req_r_msg__11__sv2v_reg,lce_req_r_msg__10__sv2v_reg,lce_req_r_msg__9__sv2v_reg,
  lce_req_r_msg__8__sv2v_reg,lce_req_r_msg__7__sv2v_reg,lce_req_r_msg__6__sv2v_reg,
  lce_req_r_msg__5__sv2v_reg,lce_req_r_msg__4__sv2v_reg,lce_req_r_msg__3__sv2v_reg,
  lce_req_r_msg__2__sv2v_reg,lce_req_r_msg__1__sv2v_reg,lce_req_r_msg__0__sv2v_reg,
  lce_req_r_addr__39__sv2v_reg,lce_req_r_addr__38__sv2v_reg,
  lce_req_r_addr__37__sv2v_reg,lce_req_r_addr__36__sv2v_reg,lce_req_r_addr__35__sv2v_reg,
  lce_req_r_addr__34__sv2v_reg,lce_req_r_addr__33__sv2v_reg,lce_req_r_addr__32__sv2v_reg,
  lce_req_r_addr__31__sv2v_reg,lce_req_r_addr__30__sv2v_reg,lce_req_r_addr__29__sv2v_reg,
  lce_req_r_addr__28__sv2v_reg,lce_req_r_addr__27__sv2v_reg,
  lce_req_r_addr__26__sv2v_reg,lce_req_r_addr__25__sv2v_reg,lce_req_r_addr__24__sv2v_reg,
  lce_req_r_addr__23__sv2v_reg,lce_req_r_addr__22__sv2v_reg,lce_req_r_addr__21__sv2v_reg,
  lce_req_r_addr__20__sv2v_reg,lce_req_r_addr__19__sv2v_reg,lce_req_r_addr__18__sv2v_reg,
  lce_req_r_addr__17__sv2v_reg,lce_req_r_addr__16__sv2v_reg,
  lce_req_r_addr__15__sv2v_reg,lce_req_r_addr__14__sv2v_reg,lce_req_r_addr__13__sv2v_reg,
  lce_req_r_addr__12__sv2v_reg,lce_req_r_addr__11__sv2v_reg,lce_req_r_addr__10__sv2v_reg,
  lce_req_r_addr__9__sv2v_reg,lce_req_r_addr__8__sv2v_reg,lce_req_r_addr__7__sv2v_reg,
  lce_req_r_addr__6__sv2v_reg,lce_req_r_addr__5__sv2v_reg,lce_req_r_addr__4__sv2v_reg,
  lce_req_r_addr__3__sv2v_reg,lce_req_r_addr__2__sv2v_reg,lce_req_r_addr__1__sv2v_reg,
  lce_req_r_addr__0__sv2v_reg,lce_req_r_src_id__5__sv2v_reg,
  lce_req_r_src_id__4__sv2v_reg,lce_req_r_src_id__3__sv2v_reg,lce_req_r_src_id__2__sv2v_reg,
  lce_req_r_src_id__1__sv2v_reg,lce_req_r_src_id__0__sv2v_reg,uc_state_1_sv2v_reg,
  uc_state_0_sv2v_reg;
  assign lce_req_r_msg__65_ = lce_req_r_msg__65__sv2v_reg;
  assign lce_req_r_msg__64_ = lce_req_r_msg__64__sv2v_reg;
  assign lce_req_r_msg__63_ = lce_req_r_msg__63__sv2v_reg;
  assign lce_req_r_msg__62_ = lce_req_r_msg__62__sv2v_reg;
  assign lce_req_r_msg__61_ = lce_req_r_msg__61__sv2v_reg;
  assign lce_req_r_msg__60_ = lce_req_r_msg__60__sv2v_reg;
  assign lce_req_r_msg__59_ = lce_req_r_msg__59__sv2v_reg;
  assign lce_req_r_msg__58_ = lce_req_r_msg__58__sv2v_reg;
  assign lce_req_r_msg__57_ = lce_req_r_msg__57__sv2v_reg;
  assign lce_req_r_msg__56_ = lce_req_r_msg__56__sv2v_reg;
  assign lce_req_r_msg__55_ = lce_req_r_msg__55__sv2v_reg;
  assign lce_req_r_msg__54_ = lce_req_r_msg__54__sv2v_reg;
  assign lce_req_r_msg__53_ = lce_req_r_msg__53__sv2v_reg;
  assign lce_req_r_msg__52_ = lce_req_r_msg__52__sv2v_reg;
  assign lce_req_r_msg__51_ = lce_req_r_msg__51__sv2v_reg;
  assign lce_req_r_msg__50_ = lce_req_r_msg__50__sv2v_reg;
  assign lce_req_r_msg__49_ = lce_req_r_msg__49__sv2v_reg;
  assign lce_req_r_msg__48_ = lce_req_r_msg__48__sv2v_reg;
  assign lce_req_r_msg__47_ = lce_req_r_msg__47__sv2v_reg;
  assign lce_req_r_msg__46_ = lce_req_r_msg__46__sv2v_reg;
  assign lce_req_r_msg__45_ = lce_req_r_msg__45__sv2v_reg;
  assign lce_req_r_msg__44_ = lce_req_r_msg__44__sv2v_reg;
  assign lce_req_r_msg__43_ = lce_req_r_msg__43__sv2v_reg;
  assign lce_req_r_msg__42_ = lce_req_r_msg__42__sv2v_reg;
  assign lce_req_r_msg__41_ = lce_req_r_msg__41__sv2v_reg;
  assign lce_req_r_msg__40_ = lce_req_r_msg__40__sv2v_reg;
  assign lce_req_r_msg__39_ = lce_req_r_msg__39__sv2v_reg;
  assign lce_req_r_msg__38_ = lce_req_r_msg__38__sv2v_reg;
  assign lce_req_r_msg__37_ = lce_req_r_msg__37__sv2v_reg;
  assign lce_req_r_msg__36_ = lce_req_r_msg__36__sv2v_reg;
  assign lce_req_r_msg__35_ = lce_req_r_msg__35__sv2v_reg;
  assign lce_req_r_msg__34_ = lce_req_r_msg__34__sv2v_reg;
  assign lce_req_r_msg__33_ = lce_req_r_msg__33__sv2v_reg;
  assign lce_req_r_msg__32_ = lce_req_r_msg__32__sv2v_reg;
  assign lce_req_r_msg__31_ = lce_req_r_msg__31__sv2v_reg;
  assign lce_req_r_msg__30_ = lce_req_r_msg__30__sv2v_reg;
  assign lce_req_r_msg__29_ = lce_req_r_msg__29__sv2v_reg;
  assign lce_req_r_msg__28_ = lce_req_r_msg__28__sv2v_reg;
  assign lce_req_r_msg__27_ = lce_req_r_msg__27__sv2v_reg;
  assign lce_req_r_msg__26_ = lce_req_r_msg__26__sv2v_reg;
  assign lce_req_r_msg__25_ = lce_req_r_msg__25__sv2v_reg;
  assign lce_req_r_msg__24_ = lce_req_r_msg__24__sv2v_reg;
  assign lce_req_r_msg__23_ = lce_req_r_msg__23__sv2v_reg;
  assign lce_req_r_msg__22_ = lce_req_r_msg__22__sv2v_reg;
  assign lce_req_r_msg__21_ = lce_req_r_msg__21__sv2v_reg;
  assign lce_req_r_msg__20_ = lce_req_r_msg__20__sv2v_reg;
  assign lce_req_r_msg__19_ = lce_req_r_msg__19__sv2v_reg;
  assign lce_req_r_msg__18_ = lce_req_r_msg__18__sv2v_reg;
  assign lce_req_r_msg__17_ = lce_req_r_msg__17__sv2v_reg;
  assign lce_req_r_msg__16_ = lce_req_r_msg__16__sv2v_reg;
  assign lce_req_r_msg__15_ = lce_req_r_msg__15__sv2v_reg;
  assign lce_req_r_msg__14_ = lce_req_r_msg__14__sv2v_reg;
  assign lce_req_r_msg__13_ = lce_req_r_msg__13__sv2v_reg;
  assign lce_req_r_msg__12_ = lce_req_r_msg__12__sv2v_reg;
  assign lce_req_r_msg__11_ = lce_req_r_msg__11__sv2v_reg;
  assign lce_req_r_msg__10_ = lce_req_r_msg__10__sv2v_reg;
  assign lce_req_r_msg__9_ = lce_req_r_msg__9__sv2v_reg;
  assign lce_req_r_msg__8_ = lce_req_r_msg__8__sv2v_reg;
  assign lce_req_r_msg__7_ = lce_req_r_msg__7__sv2v_reg;
  assign lce_req_r_msg__6_ = lce_req_r_msg__6__sv2v_reg;
  assign lce_req_r_msg__5_ = lce_req_r_msg__5__sv2v_reg;
  assign lce_req_r_msg__4_ = lce_req_r_msg__4__sv2v_reg;
  assign lce_req_r_msg__3_ = lce_req_r_msg__3__sv2v_reg;
  assign lce_req_r_msg__2_ = lce_req_r_msg__2__sv2v_reg;
  assign lce_req_r_msg__1_ = lce_req_r_msg__1__sv2v_reg;
  assign lce_req_r_msg__0_ = lce_req_r_msg__0__sv2v_reg;
  assign lce_req_r_addr__39_ = lce_req_r_addr__39__sv2v_reg;
  assign lce_req_r_addr__38_ = lce_req_r_addr__38__sv2v_reg;
  assign lce_req_r_addr__37_ = lce_req_r_addr__37__sv2v_reg;
  assign lce_req_r_addr__36_ = lce_req_r_addr__36__sv2v_reg;
  assign lce_req_r_addr__35_ = lce_req_r_addr__35__sv2v_reg;
  assign lce_req_r_addr__34_ = lce_req_r_addr__34__sv2v_reg;
  assign lce_req_r_addr__33_ = lce_req_r_addr__33__sv2v_reg;
  assign lce_req_r_addr__32_ = lce_req_r_addr__32__sv2v_reg;
  assign lce_req_r_addr__31_ = lce_req_r_addr__31__sv2v_reg;
  assign lce_req_r_addr__30_ = lce_req_r_addr__30__sv2v_reg;
  assign lce_req_r_addr__29_ = lce_req_r_addr__29__sv2v_reg;
  assign lce_req_r_addr__28_ = lce_req_r_addr__28__sv2v_reg;
  assign lce_req_r_addr__27_ = lce_req_r_addr__27__sv2v_reg;
  assign lce_req_r_addr__26_ = lce_req_r_addr__26__sv2v_reg;
  assign lce_req_r_addr__25_ = lce_req_r_addr__25__sv2v_reg;
  assign lce_req_r_addr__24_ = lce_req_r_addr__24__sv2v_reg;
  assign lce_req_r_addr__23_ = lce_req_r_addr__23__sv2v_reg;
  assign lce_req_r_addr__22_ = lce_req_r_addr__22__sv2v_reg;
  assign lce_req_r_addr__21_ = lce_req_r_addr__21__sv2v_reg;
  assign lce_req_r_addr__20_ = lce_req_r_addr__20__sv2v_reg;
  assign lce_req_r_addr__19_ = lce_req_r_addr__19__sv2v_reg;
  assign lce_req_r_addr__18_ = lce_req_r_addr__18__sv2v_reg;
  assign lce_req_r_addr__17_ = lce_req_r_addr__17__sv2v_reg;
  assign lce_req_r_addr__16_ = lce_req_r_addr__16__sv2v_reg;
  assign lce_req_r_addr__15_ = lce_req_r_addr__15__sv2v_reg;
  assign lce_req_r_addr__14_ = lce_req_r_addr__14__sv2v_reg;
  assign lce_req_r_addr__13_ = lce_req_r_addr__13__sv2v_reg;
  assign lce_req_r_addr__12_ = lce_req_r_addr__12__sv2v_reg;
  assign lce_req_r_addr__11_ = lce_req_r_addr__11__sv2v_reg;
  assign lce_req_r_addr__10_ = lce_req_r_addr__10__sv2v_reg;
  assign lce_req_r_addr__9_ = lce_req_r_addr__9__sv2v_reg;
  assign lce_req_r_addr__8_ = lce_req_r_addr__8__sv2v_reg;
  assign lce_req_r_addr__7_ = lce_req_r_addr__7__sv2v_reg;
  assign lce_req_r_addr__6_ = lce_req_r_addr__6__sv2v_reg;
  assign lce_req_r_addr__5_ = lce_req_r_addr__5__sv2v_reg;
  assign lce_req_r_addr__4_ = lce_req_r_addr__4__sv2v_reg;
  assign lce_req_r_addr__3_ = lce_req_r_addr__3__sv2v_reg;
  assign lce_req_r_addr__2_ = lce_req_r_addr__2__sv2v_reg;
  assign lce_req_r_addr__1_ = lce_req_r_addr__1__sv2v_reg;
  assign lce_req_r_addr__0_ = lce_req_r_addr__0__sv2v_reg;
  assign lce_req_r_src_id__5_ = lce_req_r_src_id__5__sv2v_reg;
  assign lce_req_r_src_id__4_ = lce_req_r_src_id__4__sv2v_reg;
  assign lce_req_r_src_id__3_ = lce_req_r_src_id__3__sv2v_reg;
  assign lce_req_r_src_id__2_ = lce_req_r_src_id__2__sv2v_reg;
  assign lce_req_r_src_id__1_ = lce_req_r_src_id__1__sv2v_reg;
  assign lce_req_r_src_id__0_ = lce_req_r_src_id__0__sv2v_reg;
  assign uc_state[1] = uc_state_1_sv2v_reg;
  assign uc_state[0] = uc_state_0_sv2v_reg;
  assign mem_cmd_o[2] = 1'b0;
  assign mem_cmd_o[3] = 1'b0;
  assign mem_cmd_o[46] = 1'b0;
  assign mem_cmd_o[47] = 1'b0;
  assign mem_cmd_o[48] = 1'b0;
  assign mem_cmd_o[49] = 1'b0;
  assign mem_cmd_o[50] = 1'b0;
  assign mem_cmd_o[51] = 1'b0;
  assign mem_cmd_o[52] = 1'b0;
  assign mem_cmd_o[53] = 1'b0;
  assign mem_cmd_o[124] = 1'b0;
  assign mem_cmd_o[125] = 1'b0;
  assign mem_cmd_o[126] = 1'b0;
  assign mem_cmd_o[127] = 1'b0;
  assign mem_cmd_o[128] = 1'b0;
  assign mem_cmd_o[129] = 1'b0;
  assign mem_cmd_o[130] = 1'b0;
  assign mem_cmd_o[131] = 1'b0;
  assign mem_cmd_o[132] = 1'b0;
  assign mem_cmd_o[133] = 1'b0;
  assign mem_cmd_o[134] = 1'b0;
  assign mem_cmd_o[135] = 1'b0;
  assign mem_cmd_o[136] = 1'b0;
  assign mem_cmd_o[137] = 1'b0;
  assign mem_cmd_o[138] = 1'b0;
  assign mem_cmd_o[139] = 1'b0;
  assign mem_cmd_o[140] = 1'b0;
  assign mem_cmd_o[141] = 1'b0;
  assign mem_cmd_o[142] = 1'b0;
  assign mem_cmd_o[143] = 1'b0;
  assign mem_cmd_o[144] = 1'b0;
  assign mem_cmd_o[145] = 1'b0;
  assign mem_cmd_o[146] = 1'b0;
  assign mem_cmd_o[147] = 1'b0;
  assign mem_cmd_o[148] = 1'b0;
  assign mem_cmd_o[149] = 1'b0;
  assign mem_cmd_o[150] = 1'b0;
  assign mem_cmd_o[151] = 1'b0;
  assign mem_cmd_o[152] = 1'b0;
  assign mem_cmd_o[153] = 1'b0;
  assign mem_cmd_o[154] = 1'b0;
  assign mem_cmd_o[155] = 1'b0;
  assign mem_cmd_o[156] = 1'b0;
  assign mem_cmd_o[157] = 1'b0;
  assign mem_cmd_o[158] = 1'b0;
  assign mem_cmd_o[159] = 1'b0;
  assign mem_cmd_o[160] = 1'b0;
  assign mem_cmd_o[161] = 1'b0;
  assign mem_cmd_o[162] = 1'b0;
  assign mem_cmd_o[163] = 1'b0;
  assign mem_cmd_o[164] = 1'b0;
  assign mem_cmd_o[165] = 1'b0;
  assign mem_cmd_o[166] = 1'b0;
  assign mem_cmd_o[167] = 1'b0;
  assign mem_cmd_o[168] = 1'b0;
  assign mem_cmd_o[169] = 1'b0;
  assign mem_cmd_o[170] = 1'b0;
  assign mem_cmd_o[171] = 1'b0;
  assign mem_cmd_o[172] = 1'b0;
  assign mem_cmd_o[173] = 1'b0;
  assign mem_cmd_o[174] = 1'b0;
  assign mem_cmd_o[175] = 1'b0;
  assign mem_cmd_o[176] = 1'b0;
  assign mem_cmd_o[177] = 1'b0;
  assign mem_cmd_o[178] = 1'b0;
  assign mem_cmd_o[179] = 1'b0;
  assign mem_cmd_o[180] = 1'b0;
  assign mem_cmd_o[181] = 1'b0;
  assign mem_cmd_o[182] = 1'b0;
  assign mem_cmd_o[183] = 1'b0;
  assign mem_cmd_o[184] = 1'b0;
  assign mem_cmd_o[185] = 1'b0;
  assign mem_cmd_o[186] = 1'b0;
  assign mem_cmd_o[187] = 1'b0;
  assign mem_cmd_o[188] = 1'b0;
  assign mem_cmd_o[189] = 1'b0;
  assign mem_cmd_o[190] = 1'b0;
  assign mem_cmd_o[191] = 1'b0;
  assign mem_cmd_o[192] = 1'b0;
  assign mem_cmd_o[193] = 1'b0;
  assign mem_cmd_o[194] = 1'b0;
  assign mem_cmd_o[195] = 1'b0;
  assign mem_cmd_o[196] = 1'b0;
  assign mem_cmd_o[197] = 1'b0;
  assign mem_cmd_o[198] = 1'b0;
  assign mem_cmd_o[199] = 1'b0;
  assign mem_cmd_o[200] = 1'b0;
  assign mem_cmd_o[201] = 1'b0;
  assign mem_cmd_o[202] = 1'b0;
  assign mem_cmd_o[203] = 1'b0;
  assign mem_cmd_o[204] = 1'b0;
  assign mem_cmd_o[205] = 1'b0;
  assign mem_cmd_o[206] = 1'b0;
  assign mem_cmd_o[207] = 1'b0;
  assign mem_cmd_o[208] = 1'b0;
  assign mem_cmd_o[209] = 1'b0;
  assign mem_cmd_o[210] = 1'b0;
  assign mem_cmd_o[211] = 1'b0;
  assign mem_cmd_o[212] = 1'b0;
  assign mem_cmd_o[213] = 1'b0;
  assign mem_cmd_o[214] = 1'b0;
  assign mem_cmd_o[215] = 1'b0;
  assign mem_cmd_o[216] = 1'b0;
  assign mem_cmd_o[217] = 1'b0;
  assign mem_cmd_o[218] = 1'b0;
  assign mem_cmd_o[219] = 1'b0;
  assign mem_cmd_o[220] = 1'b0;
  assign mem_cmd_o[221] = 1'b0;
  assign mem_cmd_o[222] = 1'b0;
  assign mem_cmd_o[223] = 1'b0;
  assign mem_cmd_o[224] = 1'b0;
  assign mem_cmd_o[225] = 1'b0;
  assign mem_cmd_o[226] = 1'b0;
  assign mem_cmd_o[227] = 1'b0;
  assign mem_cmd_o[228] = 1'b0;
  assign mem_cmd_o[229] = 1'b0;
  assign mem_cmd_o[230] = 1'b0;
  assign mem_cmd_o[231] = 1'b0;
  assign mem_cmd_o[232] = 1'b0;
  assign mem_cmd_o[233] = 1'b0;
  assign mem_cmd_o[234] = 1'b0;
  assign mem_cmd_o[235] = 1'b0;
  assign mem_cmd_o[236] = 1'b0;
  assign mem_cmd_o[237] = 1'b0;
  assign mem_cmd_o[238] = 1'b0;
  assign mem_cmd_o[239] = 1'b0;
  assign mem_cmd_o[240] = 1'b0;
  assign mem_cmd_o[241] = 1'b0;
  assign mem_cmd_o[242] = 1'b0;
  assign mem_cmd_o[243] = 1'b0;
  assign mem_cmd_o[244] = 1'b0;
  assign mem_cmd_o[245] = 1'b0;
  assign mem_cmd_o[246] = 1'b0;
  assign mem_cmd_o[247] = 1'b0;
  assign mem_cmd_o[248] = 1'b0;
  assign mem_cmd_o[249] = 1'b0;
  assign mem_cmd_o[250] = 1'b0;
  assign mem_cmd_o[251] = 1'b0;
  assign mem_cmd_o[252] = 1'b0;
  assign mem_cmd_o[253] = 1'b0;
  assign mem_cmd_o[254] = 1'b0;
  assign mem_cmd_o[255] = 1'b0;
  assign mem_cmd_o[256] = 1'b0;
  assign mem_cmd_o[257] = 1'b0;
  assign mem_cmd_o[258] = 1'b0;
  assign mem_cmd_o[259] = 1'b0;
  assign mem_cmd_o[260] = 1'b0;
  assign mem_cmd_o[261] = 1'b0;
  assign mem_cmd_o[262] = 1'b0;
  assign mem_cmd_o[263] = 1'b0;
  assign mem_cmd_o[264] = 1'b0;
  assign mem_cmd_o[265] = 1'b0;
  assign mem_cmd_o[266] = 1'b0;
  assign mem_cmd_o[267] = 1'b0;
  assign mem_cmd_o[268] = 1'b0;
  assign mem_cmd_o[269] = 1'b0;
  assign mem_cmd_o[270] = 1'b0;
  assign mem_cmd_o[271] = 1'b0;
  assign mem_cmd_o[272] = 1'b0;
  assign mem_cmd_o[273] = 1'b0;
  assign mem_cmd_o[274] = 1'b0;
  assign mem_cmd_o[275] = 1'b0;
  assign mem_cmd_o[276] = 1'b0;
  assign mem_cmd_o[277] = 1'b0;
  assign mem_cmd_o[278] = 1'b0;
  assign mem_cmd_o[279] = 1'b0;
  assign mem_cmd_o[280] = 1'b0;
  assign mem_cmd_o[281] = 1'b0;
  assign mem_cmd_o[282] = 1'b0;
  assign mem_cmd_o[283] = 1'b0;
  assign mem_cmd_o[284] = 1'b0;
  assign mem_cmd_o[285] = 1'b0;
  assign mem_cmd_o[286] = 1'b0;
  assign mem_cmd_o[287] = 1'b0;
  assign mem_cmd_o[288] = 1'b0;
  assign mem_cmd_o[289] = 1'b0;
  assign mem_cmd_o[290] = 1'b0;
  assign mem_cmd_o[291] = 1'b0;
  assign mem_cmd_o[292] = 1'b0;
  assign mem_cmd_o[293] = 1'b0;
  assign mem_cmd_o[294] = 1'b0;
  assign mem_cmd_o[295] = 1'b0;
  assign mem_cmd_o[296] = 1'b0;
  assign mem_cmd_o[297] = 1'b0;
  assign mem_cmd_o[298] = 1'b0;
  assign mem_cmd_o[299] = 1'b0;
  assign mem_cmd_o[300] = 1'b0;
  assign mem_cmd_o[301] = 1'b0;
  assign mem_cmd_o[302] = 1'b0;
  assign mem_cmd_o[303] = 1'b0;
  assign mem_cmd_o[304] = 1'b0;
  assign mem_cmd_o[305] = 1'b0;
  assign mem_cmd_o[306] = 1'b0;
  assign mem_cmd_o[307] = 1'b0;
  assign mem_cmd_o[308] = 1'b0;
  assign mem_cmd_o[309] = 1'b0;
  assign mem_cmd_o[310] = 1'b0;
  assign mem_cmd_o[311] = 1'b0;
  assign mem_cmd_o[312] = 1'b0;
  assign mem_cmd_o[313] = 1'b0;
  assign mem_cmd_o[314] = 1'b0;
  assign mem_cmd_o[315] = 1'b0;
  assign mem_cmd_o[316] = 1'b0;
  assign mem_cmd_o[317] = 1'b0;
  assign mem_cmd_o[318] = 1'b0;
  assign mem_cmd_o[319] = 1'b0;
  assign mem_cmd_o[320] = 1'b0;
  assign mem_cmd_o[321] = 1'b0;
  assign mem_cmd_o[322] = 1'b0;
  assign mem_cmd_o[323] = 1'b0;
  assign mem_cmd_o[324] = 1'b0;
  assign mem_cmd_o[325] = 1'b0;
  assign mem_cmd_o[326] = 1'b0;
  assign mem_cmd_o[327] = 1'b0;
  assign mem_cmd_o[328] = 1'b0;
  assign mem_cmd_o[329] = 1'b0;
  assign mem_cmd_o[330] = 1'b0;
  assign mem_cmd_o[331] = 1'b0;
  assign mem_cmd_o[332] = 1'b0;
  assign mem_cmd_o[333] = 1'b0;
  assign mem_cmd_o[334] = 1'b0;
  assign mem_cmd_o[335] = 1'b0;
  assign mem_cmd_o[336] = 1'b0;
  assign mem_cmd_o[337] = 1'b0;
  assign mem_cmd_o[338] = 1'b0;
  assign mem_cmd_o[339] = 1'b0;
  assign mem_cmd_o[340] = 1'b0;
  assign mem_cmd_o[341] = 1'b0;
  assign mem_cmd_o[342] = 1'b0;
  assign mem_cmd_o[343] = 1'b0;
  assign mem_cmd_o[344] = 1'b0;
  assign mem_cmd_o[345] = 1'b0;
  assign mem_cmd_o[346] = 1'b0;
  assign mem_cmd_o[347] = 1'b0;
  assign mem_cmd_o[348] = 1'b0;
  assign mem_cmd_o[349] = 1'b0;
  assign mem_cmd_o[350] = 1'b0;
  assign mem_cmd_o[351] = 1'b0;
  assign mem_cmd_o[352] = 1'b0;
  assign mem_cmd_o[353] = 1'b0;
  assign mem_cmd_o[354] = 1'b0;
  assign mem_cmd_o[355] = 1'b0;
  assign mem_cmd_o[356] = 1'b0;
  assign mem_cmd_o[357] = 1'b0;
  assign mem_cmd_o[358] = 1'b0;
  assign mem_cmd_o[359] = 1'b0;
  assign mem_cmd_o[360] = 1'b0;
  assign mem_cmd_o[361] = 1'b0;
  assign mem_cmd_o[362] = 1'b0;
  assign mem_cmd_o[363] = 1'b0;
  assign mem_cmd_o[364] = 1'b0;
  assign mem_cmd_o[365] = 1'b0;
  assign mem_cmd_o[366] = 1'b0;
  assign mem_cmd_o[367] = 1'b0;
  assign mem_cmd_o[368] = 1'b0;
  assign mem_cmd_o[369] = 1'b0;
  assign mem_cmd_o[370] = 1'b0;
  assign mem_cmd_o[371] = 1'b0;
  assign mem_cmd_o[372] = 1'b0;
  assign mem_cmd_o[373] = 1'b0;
  assign mem_cmd_o[374] = 1'b0;
  assign mem_cmd_o[375] = 1'b0;
  assign mem_cmd_o[376] = 1'b0;
  assign mem_cmd_o[377] = 1'b0;
  assign mem_cmd_o[378] = 1'b0;
  assign mem_cmd_o[379] = 1'b0;
  assign mem_cmd_o[380] = 1'b0;
  assign mem_cmd_o[381] = 1'b0;
  assign mem_cmd_o[382] = 1'b0;
  assign mem_cmd_o[383] = 1'b0;
  assign mem_cmd_o[384] = 1'b0;
  assign mem_cmd_o[385] = 1'b0;
  assign mem_cmd_o[386] = 1'b0;
  assign mem_cmd_o[387] = 1'b0;
  assign mem_cmd_o[388] = 1'b0;
  assign mem_cmd_o[389] = 1'b0;
  assign mem_cmd_o[390] = 1'b0;
  assign mem_cmd_o[391] = 1'b0;
  assign mem_cmd_o[392] = 1'b0;
  assign mem_cmd_o[393] = 1'b0;
  assign mem_cmd_o[394] = 1'b0;
  assign mem_cmd_o[395] = 1'b0;
  assign mem_cmd_o[396] = 1'b0;
  assign mem_cmd_o[397] = 1'b0;
  assign mem_cmd_o[398] = 1'b0;
  assign mem_cmd_o[399] = 1'b0;
  assign mem_cmd_o[400] = 1'b0;
  assign mem_cmd_o[401] = 1'b0;
  assign mem_cmd_o[402] = 1'b0;
  assign mem_cmd_o[403] = 1'b0;
  assign mem_cmd_o[404] = 1'b0;
  assign mem_cmd_o[405] = 1'b0;
  assign mem_cmd_o[406] = 1'b0;
  assign mem_cmd_o[407] = 1'b0;
  assign mem_cmd_o[408] = 1'b0;
  assign mem_cmd_o[409] = 1'b0;
  assign mem_cmd_o[410] = 1'b0;
  assign mem_cmd_o[411] = 1'b0;
  assign mem_cmd_o[412] = 1'b0;
  assign mem_cmd_o[413] = 1'b0;
  assign mem_cmd_o[414] = 1'b0;
  assign mem_cmd_o[415] = 1'b0;
  assign mem_cmd_o[416] = 1'b0;
  assign mem_cmd_o[417] = 1'b0;
  assign mem_cmd_o[418] = 1'b0;
  assign mem_cmd_o[419] = 1'b0;
  assign mem_cmd_o[420] = 1'b0;
  assign mem_cmd_o[421] = 1'b0;
  assign mem_cmd_o[422] = 1'b0;
  assign mem_cmd_o[423] = 1'b0;
  assign mem_cmd_o[424] = 1'b0;
  assign mem_cmd_o[425] = 1'b0;
  assign mem_cmd_o[426] = 1'b0;
  assign mem_cmd_o[427] = 1'b0;
  assign mem_cmd_o[428] = 1'b0;
  assign mem_cmd_o[429] = 1'b0;
  assign mem_cmd_o[430] = 1'b0;
  assign mem_cmd_o[431] = 1'b0;
  assign mem_cmd_o[432] = 1'b0;
  assign mem_cmd_o[433] = 1'b0;
  assign mem_cmd_o[434] = 1'b0;
  assign mem_cmd_o[435] = 1'b0;
  assign mem_cmd_o[436] = 1'b0;
  assign mem_cmd_o[437] = 1'b0;
  assign mem_cmd_o[438] = 1'b0;
  assign mem_cmd_o[439] = 1'b0;
  assign mem_cmd_o[440] = 1'b0;
  assign mem_cmd_o[441] = 1'b0;
  assign mem_cmd_o[442] = 1'b0;
  assign mem_cmd_o[443] = 1'b0;
  assign mem_cmd_o[444] = 1'b0;
  assign mem_cmd_o[445] = 1'b0;
  assign mem_cmd_o[446] = 1'b0;
  assign mem_cmd_o[447] = 1'b0;
  assign mem_cmd_o[448] = 1'b0;
  assign mem_cmd_o[449] = 1'b0;
  assign mem_cmd_o[450] = 1'b0;
  assign mem_cmd_o[451] = 1'b0;
  assign mem_cmd_o[452] = 1'b0;
  assign mem_cmd_o[453] = 1'b0;
  assign mem_cmd_o[454] = 1'b0;
  assign mem_cmd_o[455] = 1'b0;
  assign mem_cmd_o[456] = 1'b0;
  assign mem_cmd_o[457] = 1'b0;
  assign mem_cmd_o[458] = 1'b0;
  assign mem_cmd_o[459] = 1'b0;
  assign mem_cmd_o[460] = 1'b0;
  assign mem_cmd_o[461] = 1'b0;
  assign mem_cmd_o[462] = 1'b0;
  assign mem_cmd_o[463] = 1'b0;
  assign mem_cmd_o[464] = 1'b0;
  assign mem_cmd_o[465] = 1'b0;
  assign mem_cmd_o[466] = 1'b0;
  assign mem_cmd_o[467] = 1'b0;
  assign mem_cmd_o[468] = 1'b0;
  assign mem_cmd_o[469] = 1'b0;
  assign mem_cmd_o[470] = 1'b0;
  assign mem_cmd_o[471] = 1'b0;
  assign mem_cmd_o[472] = 1'b0;
  assign mem_cmd_o[473] = 1'b0;
  assign mem_cmd_o[474] = 1'b0;
  assign mem_cmd_o[475] = 1'b0;
  assign mem_cmd_o[476] = 1'b0;
  assign mem_cmd_o[477] = 1'b0;
  assign mem_cmd_o[478] = 1'b0;
  assign mem_cmd_o[479] = 1'b0;
  assign mem_cmd_o[480] = 1'b0;
  assign mem_cmd_o[481] = 1'b0;
  assign mem_cmd_o[482] = 1'b0;
  assign mem_cmd_o[483] = 1'b0;
  assign mem_cmd_o[484] = 1'b0;
  assign mem_cmd_o[485] = 1'b0;
  assign mem_cmd_o[486] = 1'b0;
  assign mem_cmd_o[487] = 1'b0;
  assign mem_cmd_o[488] = 1'b0;
  assign mem_cmd_o[489] = 1'b0;
  assign mem_cmd_o[490] = 1'b0;
  assign mem_cmd_o[491] = 1'b0;
  assign mem_cmd_o[492] = 1'b0;
  assign mem_cmd_o[493] = 1'b0;
  assign mem_cmd_o[494] = 1'b0;
  assign mem_cmd_o[495] = 1'b0;
  assign mem_cmd_o[496] = 1'b0;
  assign mem_cmd_o[497] = 1'b0;
  assign mem_cmd_o[498] = 1'b0;
  assign mem_cmd_o[499] = 1'b0;
  assign mem_cmd_o[500] = 1'b0;
  assign mem_cmd_o[501] = 1'b0;
  assign mem_cmd_o[502] = 1'b0;
  assign mem_cmd_o[503] = 1'b0;
  assign mem_cmd_o[504] = 1'b0;
  assign mem_cmd_o[505] = 1'b0;
  assign mem_cmd_o[506] = 1'b0;
  assign mem_cmd_o[507] = 1'b0;
  assign mem_cmd_o[508] = 1'b0;
  assign mem_cmd_o[509] = 1'b0;
  assign mem_cmd_o[510] = 1'b0;
  assign mem_cmd_o[511] = 1'b0;
  assign mem_cmd_o[512] = 1'b0;
  assign mem_cmd_o[513] = 1'b0;
  assign mem_cmd_o[514] = 1'b0;
  assign mem_cmd_o[515] = 1'b0;
  assign mem_cmd_o[516] = 1'b0;
  assign mem_cmd_o[517] = 1'b0;
  assign mem_cmd_o[518] = 1'b0;
  assign mem_cmd_o[519] = 1'b0;
  assign mem_cmd_o[520] = 1'b0;
  assign mem_cmd_o[521] = 1'b0;
  assign mem_cmd_o[522] = 1'b0;
  assign mem_cmd_o[523] = 1'b0;
  assign mem_cmd_o[524] = 1'b0;
  assign mem_cmd_o[525] = 1'b0;
  assign mem_cmd_o[526] = 1'b0;
  assign mem_cmd_o[527] = 1'b0;
  assign mem_cmd_o[528] = 1'b0;
  assign mem_cmd_o[529] = 1'b0;
  assign mem_cmd_o[530] = 1'b0;
  assign mem_cmd_o[531] = 1'b0;
  assign mem_cmd_o[532] = 1'b0;
  assign mem_cmd_o[533] = 1'b0;
  assign mem_cmd_o[534] = 1'b0;
  assign mem_cmd_o[535] = 1'b0;
  assign mem_cmd_o[536] = 1'b0;
  assign mem_cmd_o[537] = 1'b0;
  assign mem_cmd_o[538] = 1'b0;
  assign mem_cmd_o[539] = 1'b0;
  assign mem_cmd_o[540] = 1'b0;
  assign mem_cmd_o[541] = 1'b0;
  assign mem_cmd_o[542] = 1'b0;
  assign mem_cmd_o[543] = 1'b0;
  assign mem_cmd_o[544] = 1'b0;
  assign mem_cmd_o[545] = 1'b0;
  assign mem_cmd_o[546] = 1'b0;
  assign mem_cmd_o[547] = 1'b0;
  assign mem_cmd_o[548] = 1'b0;
  assign mem_cmd_o[549] = 1'b0;
  assign mem_cmd_o[550] = 1'b0;
  assign mem_cmd_o[551] = 1'b0;
  assign mem_cmd_o[552] = 1'b0;
  assign mem_cmd_o[553] = 1'b0;
  assign mem_cmd_o[554] = 1'b0;
  assign mem_cmd_o[555] = 1'b0;
  assign mem_cmd_o[556] = 1'b0;
  assign mem_cmd_o[557] = 1'b0;
  assign mem_cmd_o[558] = 1'b0;
  assign mem_cmd_o[559] = 1'b0;
  assign mem_cmd_o[560] = 1'b0;
  assign mem_cmd_o[561] = 1'b0;
  assign mem_cmd_o[562] = 1'b0;
  assign mem_cmd_o[563] = 1'b0;
  assign mem_cmd_o[564] = 1'b0;
  assign mem_cmd_o[565] = 1'b0;
  assign mem_cmd_o[566] = 1'b0;
  assign mem_cmd_o[567] = 1'b0;
  assign mem_cmd_o[568] = 1'b0;
  assign mem_cmd_o[569] = 1'b0;
  assign mem_cmd_o[570] = 1'b0;
  assign mem_cmd_o[571] = 1'b0;
  assign lce_cmd_o[10] = 1'b0;
  assign lce_cmd_o[11] = 1'b0;
  assign lce_cmd_o[12] = 1'b0;

  always @(posedge clk_i) begin
    if(N1650) begin
      lce_req_r_msg__65__sv2v_reg <= N127;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__64__sv2v_reg <= N126;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__63__sv2v_reg <= N125;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__62__sv2v_reg <= N124;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__61__sv2v_reg <= N123;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__60__sv2v_reg <= N122;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__59__sv2v_reg <= N121;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__58__sv2v_reg <= N120;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__57__sv2v_reg <= N119;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__56__sv2v_reg <= N118;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__55__sv2v_reg <= N117;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__54__sv2v_reg <= N116;
    end 
  end


  always @(posedge clk_i) begin
    if(N1664) begin
      lce_req_r_msg__53__sv2v_reg <= N115;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__52__sv2v_reg <= N114;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__51__sv2v_reg <= N113;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__50__sv2v_reg <= N112;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__49__sv2v_reg <= N111;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__48__sv2v_reg <= N110;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__47__sv2v_reg <= N109;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__46__sv2v_reg <= N108;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__45__sv2v_reg <= N107;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__44__sv2v_reg <= N106;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__43__sv2v_reg <= N105;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__42__sv2v_reg <= N104;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__41__sv2v_reg <= N103;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__40__sv2v_reg <= N102;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__39__sv2v_reg <= N101;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__38__sv2v_reg <= N100;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__37__sv2v_reg <= N99;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__36__sv2v_reg <= N98;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__35__sv2v_reg <= N97;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__34__sv2v_reg <= N96;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__33__sv2v_reg <= N95;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__32__sv2v_reg <= N94;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__31__sv2v_reg <= N93;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__30__sv2v_reg <= N92;
    end 
  end


  always @(posedge clk_i) begin
    if(N1675) begin
      lce_req_r_msg__29__sv2v_reg <= N91;
    end 
  end


  always @(posedge clk_i) begin
    if(N1679) begin
      lce_req_r_msg__28__sv2v_reg <= N90;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__27__sv2v_reg <= N89;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__26__sv2v_reg <= N88;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__25__sv2v_reg <= N87;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__24__sv2v_reg <= N86;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__23__sv2v_reg <= N85;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__22__sv2v_reg <= N84;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__21__sv2v_reg <= N83;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__20__sv2v_reg <= N82;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__19__sv2v_reg <= N81;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__18__sv2v_reg <= N80;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__17__sv2v_reg <= N79;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__16__sv2v_reg <= N78;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__15__sv2v_reg <= N77;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__14__sv2v_reg <= N76;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__13__sv2v_reg <= N75;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__12__sv2v_reg <= N74;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__11__sv2v_reg <= N73;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__10__sv2v_reg <= N72;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__9__sv2v_reg <= N71;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__8__sv2v_reg <= N70;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__7__sv2v_reg <= N69;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__6__sv2v_reg <= N68;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__5__sv2v_reg <= N67;
    end 
  end


  always @(posedge clk_i) begin
    if(N1688) begin
      lce_req_r_msg__4__sv2v_reg <= N66;
    end 
  end


  always @(posedge clk_i) begin
    if(N1695) begin
      lce_req_r_msg__3__sv2v_reg <= N65;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_msg__2__sv2v_reg <= N64;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_msg__1__sv2v_reg <= N63;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_msg__0__sv2v_reg <= N62;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__39__sv2v_reg <= N61;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__38__sv2v_reg <= N60;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__37__sv2v_reg <= N59;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__36__sv2v_reg <= N58;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__35__sv2v_reg <= N57;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__34__sv2v_reg <= N56;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__33__sv2v_reg <= N55;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__32__sv2v_reg <= N54;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__31__sv2v_reg <= N53;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__30__sv2v_reg <= N52;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__29__sv2v_reg <= N51;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__28__sv2v_reg <= N50;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__27__sv2v_reg <= N49;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__26__sv2v_reg <= N48;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__25__sv2v_reg <= N47;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__24__sv2v_reg <= N46;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__23__sv2v_reg <= N45;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__22__sv2v_reg <= N44;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__21__sv2v_reg <= N43;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__20__sv2v_reg <= N42;
    end 
  end


  always @(posedge clk_i) begin
    if(N1702) begin
      lce_req_r_addr__19__sv2v_reg <= N41;
    end 
  end


  always @(posedge clk_i) begin
    if(N1712) begin
      lce_req_r_addr__18__sv2v_reg <= N40;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__17__sv2v_reg <= N39;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__16__sv2v_reg <= N38;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__15__sv2v_reg <= N37;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__14__sv2v_reg <= N36;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__13__sv2v_reg <= N35;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__12__sv2v_reg <= N34;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__11__sv2v_reg <= N33;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__10__sv2v_reg <= N32;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__9__sv2v_reg <= N31;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__8__sv2v_reg <= N30;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__7__sv2v_reg <= N29;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__6__sv2v_reg <= N28;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__5__sv2v_reg <= N27;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__4__sv2v_reg <= N26;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__3__sv2v_reg <= N25;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__2__sv2v_reg <= N24;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__1__sv2v_reg <= N23;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_addr__0__sv2v_reg <= N22;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__5__sv2v_reg <= N21;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__4__sv2v_reg <= N20;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__3__sv2v_reg <= N19;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__2__sv2v_reg <= N18;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__1__sv2v_reg <= N17;
    end 
  end


  always @(posedge clk_i) begin
    if(N1717) begin
      lce_req_r_src_id__0__sv2v_reg <= N16;
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      uc_state_1_sv2v_reg <= N15;
    end 
  end


  always @(posedge clk_i) begin
    if(1'b1) begin
      uc_state_0_sv2v_reg <= N14;
    end 
  end

  assign N131 = N129 & N130;
  assign N132 = uc_state[1] | N130;
  assign N134 = N129 | uc_state[0];
  assign N136 = uc_state[1] & uc_state[0];
  assign N1718 = ~lce_req_r_msg__1_;
  assign N1719 = lce_req_r_msg__0_ | N1718;
  assign N1720 = ~N1719;
  assign N1721 = lce_req_r_msg__0_ | N1718;
  assign N1722 = ~N1721;
  assign N1723 = ~lce_req_r_msg__0_;
  assign N1724 = N1723 | lce_req_r_msg__1_;
  assign N1725 = ~N1724;
  assign N1726 = lce_req_r_msg__0_ | lce_req_r_msg__1_;
  assign N1727 = ~N1726;
  assign N1728 = N1723 | lce_req_r_msg__1_;
  assign N1729 = ~N1728;
  assign N1730 = lce_req_r_msg__0_ | lce_req_r_msg__1_;
  assign N1731 = ~N1730;
  assign N1732 = ~lce_req_i[11];
  assign N1733 = N1732 | lce_req_i[12];
  assign N1734 = lce_req_i[10] | N1733;
  assign N1735 = ~N1734;
  assign N1736 = mem_resp_i[0] | N1741;
  assign N1737 = ~N1736;
  assign N1738 = ~mem_resp_i[1];
  assign N1739 = ~mem_resp_i[0];
  assign N1740 = mem_resp_i[2] | mem_resp_i[3];
  assign N1741 = N1738 | N1740;
  assign N1742 = N1739 | N1741;
  assign N1743 = ~N1742;
  assign { N15, N14 } = (N0)? { 1'b0, 1'b0 } : 
                        (N1)? uc_state_n : 1'b0;
  assign N0 = reset_i;
  assign N1 = N128;
  assign { N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N1)? { N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403 } : 1'b0;
  assign N143 = (N2)? lce_cmd_ready_i : 
                (N1630)? lce_cmd_ready_i : 
                (N142)? 1'b0 : 
                (N3)? 1'b0 : 1'b0;
  assign N2 = N137;
  assign N3 = 1'b0;
  assign { N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N151, N150, N149, N148, N147, N146, N145, N144 } = (N2)? { mem_resp_i[60:60], 1'b0, 1'b0, 1'b0, mem_resp_i[43:4], 1'b0, 1'b1, mem_resp_i[59:54] } : 
                                                                                                                                                                                                                                                                                                                                      (N1630)? { mem_resp_i[43:4], cce_id_i, 1'b1, 1'b1, mem_resp_i[59:54] } : 
                                                                                                                                                                                                                                                                                                                                      (N142)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                      (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N153 } = (N2)? { mem_resp_i[571:61], 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N152)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709 } = (N1630)? { lce_req_r_msg__65_, lce_req_r_msg__64_, lce_req_r_msg__63_, lce_req_r_msg__62_, lce_req_r_msg__61_, lce_req_r_msg__60_, lce_req_r_msg__59_, lce_req_r_msg__58_, lce_req_r_msg__57_, lce_req_r_msg__56_, lce_req_r_msg__55_, lce_req_r_msg__54_, lce_req_r_msg__53_, lce_req_r_msg__52_, lce_req_r_msg__51_, lce_req_r_msg__50_, lce_req_r_msg__49_, lce_req_r_msg__48_, lce_req_r_msg__47_, lce_req_r_msg__46_, lce_req_r_msg__45_, lce_req_r_msg__44_, lce_req_r_msg__43_, lce_req_r_msg__42_, lce_req_r_msg__41_, lce_req_r_msg__40_, lce_req_r_msg__39_, lce_req_r_msg__38_, lce_req_r_msg__37_, lce_req_r_msg__36_, lce_req_r_msg__35_, lce_req_r_msg__34_, lce_req_r_msg__33_, lce_req_r_msg__32_, lce_req_r_msg__31_, lce_req_r_msg__30_, lce_req_r_msg__29_, lce_req_r_msg__28_, lce_req_r_msg__27_, lce_req_r_msg__26_, lce_req_r_msg__25_, lce_req_r_msg__24_, lce_req_r_msg__23_, lce_req_r_msg__22_, lce_req_r_msg__21_, lce_req_r_msg__20_, lce_req_r_msg__19_, lce_req_r_msg__18_, lce_req_r_msg__17_, lce_req_r_msg__16_, lce_req_r_msg__15_, lce_req_r_msg__14_, lce_req_r_msg__13_, lce_req_r_msg__12_, lce_req_r_msg__11_, lce_req_r_msg__10_, lce_req_r_msg__9_, lce_req_r_msg__8_, lce_req_r_msg__7_, lce_req_r_msg__6_, lce_req_r_msg__5_, lce_req_r_msg__4_, lce_req_r_msg__3_, lce_req_r_msg__2_, lce_req_r_msg__1_, lce_req_r_msg__0_, lce_req_r_addr__39_, lce_req_r_addr__38_, lce_req_r_addr__37_, lce_req_r_addr__36_, lce_req_r_addr__35_, lce_req_r_addr__34_, lce_req_r_addr__33_, lce_req_r_addr__32_, lce_req_r_addr__31_, lce_req_r_addr__30_, lce_req_r_addr__29_, lce_req_r_addr__28_, lce_req_r_addr__27_, lce_req_r_addr__26_, lce_req_r_addr__25_, lce_req_r_addr__24_, lce_req_r_addr__23_, lce_req_r_addr__22_, lce_req_r_addr__21_, lce_req_r_addr__20_, lce_req_r_addr__19_, lce_req_r_addr__18_, lce_req_r_addr__17_, lce_req_r_addr__16_, lce_req_r_addr__15_, lce_req_r_addr__14_, lce_req_r_addr__13_, lce_req_r_addr__12_, lce_req_r_addr__11_, lce_req_r_addr__10_, lce_req_r_addr__9_, lce_req_r_addr__8_, lce_req_r_addr__7_, lce_req_r_addr__6_, lce_req_r_addr__5_, lce_req_r_addr__4_, lce_req_r_addr__3_, lce_req_r_addr__2_, lce_req_r_addr__1_, lce_req_r_addr__0_, lce_req_r_src_id__5_, lce_req_r_src_id__4_, lce_req_r_src_id__3_, lce_req_r_src_id__2_, lce_req_r_src_id__1_, lce_req_r_src_id__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1633)? { lce_req_i[118:13], lce_req_i[9:4] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N141)? { lce_req_r_msg__65_, lce_req_r_msg__64_, lce_req_r_msg__63_, lce_req_r_msg__62_, lce_req_r_msg__61_, lce_req_r_msg__60_, lce_req_r_msg__59_, lce_req_r_msg__58_, lce_req_r_msg__57_, lce_req_r_msg__56_, lce_req_r_msg__55_, lce_req_r_msg__54_, lce_req_r_msg__53_, lce_req_r_msg__52_, lce_req_r_msg__51_, lce_req_r_msg__50_, lce_req_r_msg__49_, lce_req_r_msg__48_, lce_req_r_msg__47_, lce_req_r_msg__46_, lce_req_r_msg__45_, lce_req_r_msg__44_, lce_req_r_msg__43_, lce_req_r_msg__42_, lce_req_r_msg__41_, lce_req_r_msg__40_, lce_req_r_msg__39_, lce_req_r_msg__38_, lce_req_r_msg__37_, lce_req_r_msg__36_, lce_req_r_msg__35_, lce_req_r_msg__34_, lce_req_r_msg__33_, lce_req_r_msg__32_, lce_req_r_msg__31_, lce_req_r_msg__30_, lce_req_r_msg__29_, lce_req_r_msg__28_, lce_req_r_msg__27_, lce_req_r_msg__26_, lce_req_r_msg__25_, lce_req_r_msg__24_, lce_req_r_msg__23_, lce_req_r_msg__22_, lce_req_r_msg__21_, lce_req_r_msg__20_, lce_req_r_msg__19_, lce_req_r_msg__18_, lce_req_r_msg__17_, lce_req_r_msg__16_, lce_req_r_msg__15_, lce_req_r_msg__14_, lce_req_r_msg__13_, lce_req_r_msg__12_, lce_req_r_msg__11_, lce_req_r_msg__10_, lce_req_r_msg__9_, lce_req_r_msg__8_, lce_req_r_msg__7_, lce_req_r_msg__6_, lce_req_r_msg__5_, lce_req_r_msg__4_, lce_req_r_msg__3_, lce_req_r_msg__2_, lce_req_r_msg__1_, lce_req_r_msg__0_, lce_req_r_addr__39_, lce_req_r_addr__38_, lce_req_r_addr__37_, lce_req_r_addr__36_, lce_req_r_addr__35_, lce_req_r_addr__34_, lce_req_r_addr__33_, lce_req_r_addr__32_, lce_req_r_addr__31_, lce_req_r_addr__30_, lce_req_r_addr__29_, lce_req_r_addr__28_, lce_req_r_addr__27_, lce_req_r_addr__26_, lce_req_r_addr__25_, lce_req_r_addr__24_, lce_req_r_addr__23_, lce_req_r_addr__22_, lce_req_r_addr__21_, lce_req_r_addr__20_, lce_req_r_addr__19_, lce_req_r_addr__18_, lce_req_r_addr__17_, lce_req_r_addr__16_, lce_req_r_addr__15_, lce_req_r_addr__14_, lce_req_r_addr__13_, lce_req_r_addr__12_, lce_req_r_addr__11_, lce_req_r_addr__10_, lce_req_r_addr__9_, lce_req_r_addr__8_, lce_req_r_addr__7_, lce_req_r_addr__6_, lce_req_r_addr__5_, lce_req_r_addr__4_, lce_req_r_addr__3_, lce_req_r_addr__2_, lce_req_r_addr__1_, lce_req_r_addr__0_, lce_req_r_src_id__5_, lce_req_r_src_id__4_, lce_req_r_src_id__3_, lce_req_r_src_id__2_, lce_req_r_src_id__1_, lce_req_r_src_id__0_ } : 1'b0;
  assign N821 = (N2)? 1'b0 : 
                (N1630)? 1'b0 : 
                (N1633)? lce_req_v_i : 
                (N141)? 1'b0 : 1'b0;
  assign { N823, N822 } = (N2)? { 1'b0, 1'b0 } : 
                          (N1630)? { 1'b0, 1'b0 } : 
                          (N1633)? { N1734, N1735 } : 
                          (N141)? { 1'b0, 1'b0 } : 1'b0;
  assign { N828, N827 } = (N4)? { 1'b0, 1'b0 } : 
                          (N5)? { 1'b0, 1'b1 } : 
                          (N6)? { 1'b1, 1'b0 } : 
                          (N826)? { 1'b1, 1'b1 } : 1'b0;
  assign N4 = N1727;
  assign N5 = N1725;
  assign N6 = N1720;
  assign { N833, N832 } = (N7)? { 1'b0, 1'b0 } : 
                          (N8)? { 1'b0, 1'b1 } : 
                          (N9)? { 1'b1, 1'b0 } : 
                          (N831)? { 1'b1, 1'b1 } : 1'b0;
  assign N7 = N1731;
  assign N8 = N1729;
  assign N9 = N1722;
  assign { N836, N835 } = (N10)? { N823, N822 } : 
                          (N11)? { 1'b0, N834 } : 
                          (N12)? { N834, 1'b0 } : 
                          (N13)? { 1'b0, 1'b0 } : 1'b0;
  assign N10 = N131;
  assign N11 = N133;
  assign N12 = N135;
  assign N13 = N136;
  assign N837 = (N10)? N821 : 
                (N11)? 1'b0 : 
                (N12)? 1'b0 : 
                (N13)? 1'b0 : 1'b0;
  assign N838 = (N10)? N143 : 
                (N11)? 1'b0 : 
                (N12)? 1'b0 : 
                (N13)? 1'b0 : 1'b0;
  assign { N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839 } = (N10)? { N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N151, N150, N149, N148, N147, N146, N145, N144 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403 } = (N10)? { N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1515 = (N10)? 1'b0 : 
                 (N11)? mem_cmd_ready_i : 
                 (N12)? mem_cmd_ready_i : 
                 (N13)? 1'b0 : 1'b0;
  assign { N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516 } = (N10)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_req_r_src_id__5_, lce_req_r_src_id__4_, lce_req_r_src_id__3_, lce_req_r_src_id__2_, lce_req_r_src_id__1_, lce_req_r_src_id__0_, N828, N827, lce_req_r_addr__39_, lce_req_r_addr__38_, lce_req_r_addr__37_, lce_req_r_addr__36_, lce_req_r_addr__35_, lce_req_r_addr__34_, lce_req_r_addr__33_, lce_req_r_addr__32_, lce_req_r_addr__31_, lce_req_r_addr__30_, lce_req_r_addr__29_, lce_req_r_addr__28_, lce_req_r_addr__27_, lce_req_r_addr__26_, lce_req_r_addr__25_, lce_req_r_addr__24_, lce_req_r_addr__23_, lce_req_r_addr__22_, lce_req_r_addr__21_, lce_req_r_addr__20_, lce_req_r_addr__19_, lce_req_r_addr__18_, lce_req_r_addr__17_, lce_req_r_addr__16_, lce_req_r_addr__15_, lce_req_r_addr__14_, lce_req_r_addr__13_, lce_req_r_addr__12_, lce_req_r_addr__11_, lce_req_r_addr__10_, lce_req_r_addr__9_, lce_req_r_addr__8_, lce_req_r_addr__7_, lce_req_r_addr__6_, lce_req_r_addr__5_, lce_req_r_addr__4_, lce_req_r_addr__3_, lce_req_r_addr__2_, lce_req_r_addr__1_, lce_req_r_addr__0_, 1'b1, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N12)? { lce_req_r_msg__65_, lce_req_r_msg__64_, lce_req_r_msg__63_, lce_req_r_msg__62_, lce_req_r_msg__61_, lce_req_r_msg__60_, lce_req_r_msg__59_, lce_req_r_msg__58_, lce_req_r_msg__57_, lce_req_r_msg__56_, lce_req_r_msg__55_, lce_req_r_msg__54_, lce_req_r_msg__53_, lce_req_r_msg__52_, lce_req_r_msg__51_, lce_req_r_msg__50_, lce_req_r_msg__49_, lce_req_r_msg__48_, lce_req_r_msg__47_, lce_req_r_msg__46_, lce_req_r_msg__45_, lce_req_r_msg__44_, lce_req_r_msg__43_, lce_req_r_msg__42_, lce_req_r_msg__41_, lce_req_r_msg__40_, lce_req_r_msg__39_, lce_req_r_msg__38_, lce_req_r_msg__37_, lce_req_r_msg__36_, lce_req_r_msg__35_, lce_req_r_msg__34_, lce_req_r_msg__33_, lce_req_r_msg__32_, lce_req_r_msg__31_, lce_req_r_msg__30_, lce_req_r_msg__29_, lce_req_r_msg__28_, lce_req_r_msg__27_, lce_req_r_msg__26_, lce_req_r_msg__25_, lce_req_r_msg__24_, lce_req_r_msg__23_, lce_req_r_msg__22_, lce_req_r_msg__21_, lce_req_r_msg__20_, lce_req_r_msg__19_, lce_req_r_msg__18_, lce_req_r_msg__17_, lce_req_r_msg__16_, lce_req_r_msg__15_, lce_req_r_msg__14_, lce_req_r_msg__13_, lce_req_r_msg__12_, lce_req_r_msg__11_, lce_req_r_msg__10_, lce_req_r_msg__9_, lce_req_r_msg__8_, lce_req_r_msg__7_, lce_req_r_msg__6_, lce_req_r_msg__5_, lce_req_r_msg__4_, lce_req_r_msg__3_, lce_req_r_msg__2_, lce_req_r_src_id__5_, lce_req_r_src_id__4_, lce_req_r_src_id__3_, lce_req_r_src_id__2_, lce_req_r_src_id__1_, lce_req_r_src_id__0_, N833, N832, lce_req_r_addr__39_, lce_req_r_addr__38_, lce_req_r_addr__37_, lce_req_r_addr__36_, lce_req_r_addr__35_, lce_req_r_addr__34_, lce_req_r_addr__33_, lce_req_r_addr__32_, lce_req_r_addr__31_, lce_req_r_addr__30_, lce_req_r_addr__29_, lce_req_r_addr__28_, lce_req_r_addr__27_, lce_req_r_addr__26_, lce_req_r_addr__25_, lce_req_r_addr__24_, lce_req_r_addr__23_, lce_req_r_addr__22_, lce_req_r_addr__21_, lce_req_r_addr__20_, lce_req_r_addr__19_, lce_req_r_addr__18_, lce_req_r_addr__17_, lce_req_r_addr__16_, lce_req_r_addr__15_, lce_req_r_addr__14_, lce_req_r_addr__13_, lce_req_r_addr__12_, lce_req_r_addr__11_, lce_req_r_addr__10_, lce_req_r_addr__9_, lce_req_r_addr__8_, lce_req_r_addr__7_, lce_req_r_addr__6_, lce_req_r_addr__5_, lce_req_r_addr__4_, lce_req_r_addr__3_, lce_req_r_addr__2_, lce_req_r_addr__1_, lce_req_r_addr__0_, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N13)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { mem_cmd_o[123:54], mem_cmd_o[45:4], mem_cmd_o[1:0] } = (N1)? { N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516 } : 
                                                                  (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign uc_state_n = (N1)? { N836, N835 } : 
                      (N0)? { 1'b0, 1'b0 } : 1'b0;
  assign lce_req_yumi_o = (N1)? N837 : 
                          (N0)? 1'b0 : 1'b0;
  assign lce_cmd_v_o = (N1)? N838 : 
                       (N0)? 1'b0 : 1'b0;
  assign { lce_cmd_o[567:13], lce_cmd_o[9:0] } = (N1)? { N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N846, N845, N844, N843, N842, N841, N840, N839 } : 
                                                 (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign mem_resp_yumi_o = (N1)? N838 : 
                           (N0)? 1'b0 : 1'b0;
  assign mem_cmd_v_o = (N1)? N1515 : 
                       (N0)? 1'b0 : 1'b0;
  assign N128 = ~reset_i;
  assign N129 = ~uc_state[1];
  assign N130 = ~uc_state[0];
  assign N133 = ~N132;
  assign N135 = ~N134;
  assign N137 = mem_resp_v_i & N1737;
  assign N138 = mem_resp_v_i & N1743;
  assign N139 = N138 | N137;
  assign N140 = lce_req_v_i | N139;
  assign N141 = ~N140;
  assign N142 = ~N139;
  assign N152 = ~N137;
  assign N824 = N1725 | N1727;
  assign N825 = N1720 | N824;
  assign N826 = ~N825;
  assign N829 = N1729 | N1731;
  assign N830 = N1722 | N829;
  assign N831 = ~N830;
  assign N834 = ~mem_cmd_ready_i;
  assign N1630 = N138 & N152;
  assign N1631 = ~N138;
  assign N1632 = N152 & N1631;
  assign N1633 = lce_req_v_i & N1632;
  assign N1634 = N128 & N128;
  assign N1635 = N131 & N1634;
  assign N1636 = N137 & N1635;
  assign N1637 = N128 & N128;
  assign N1638 = N133 & N1637;
  assign N1639 = N834 & N1638;
  assign N1640 = N1636 | N1639;
  assign N1641 = N128 & N128;
  assign N1642 = N135 & N1641;
  assign N1643 = N834 & N1642;
  assign N1644 = N1640 | N1643;
  assign N1645 = N128 & N128;
  assign N1646 = N136 & N1645;
  assign N1647 = N1644 | N1646;
  assign N1648 = reset_i & N128;
  assign N1649 = N1647 | N1648;
  assign N1650 = ~N1649;
  assign N1651 = N128 & N128;
  assign N1652 = N131 & N1651;
  assign N1653 = N137 & N1652;
  assign N1654 = N133 & N1651;
  assign N1655 = N834 & N1654;
  assign N1656 = N1653 | N1655;
  assign N1657 = N135 & N1651;
  assign N1658 = N834 & N1657;
  assign N1659 = N1656 | N1658;
  assign N1660 = N136 & N1651;
  assign N1661 = N1659 | N1660;
  assign N1662 = reset_i & N128;
  assign N1663 = N1661 | N1662;
  assign N1664 = ~N1663;
  assign N1665 = N131 & N1645;
  assign N1666 = N137 & N1665;
  assign N1667 = N133 & N1645;
  assign N1668 = N834 & N1667;
  assign N1669 = N1666 | N1668;
  assign N1670 = N135 & N1645;
  assign N1671 = N834 & N1670;
  assign N1672 = N1669 | N1671;
  assign N1673 = N1672 | N1646;
  assign N1674 = N1673 | N1648;
  assign N1675 = ~N1674;
  assign N1676 = N136 & N1641;
  assign N1677 = N1672 | N1676;
  assign N1678 = N1677 | N1648;
  assign N1679 = ~N1678;
  assign N1680 = N131 & N1641;
  assign N1681 = N137 & N1680;
  assign N1682 = N133 & N1641;
  assign N1683 = N834 & N1682;
  assign N1684 = N1681 | N1683;
  assign N1685 = N1684 | N1643;
  assign N1686 = N1685 | N1676;
  assign N1687 = N1686 | N1648;
  assign N1688 = ~N1687;
  assign N1689 = N135 & N1637;
  assign N1690 = N834 & N1689;
  assign N1691 = N1684 | N1690;
  assign N1692 = N136 & N1637;
  assign N1693 = N1691 | N1692;
  assign N1694 = N1693 | N1648;
  assign N1695 = ~N1694;
  assign N1696 = N131 & N1637;
  assign N1697 = N137 & N1696;
  assign N1698 = N1697 | N1639;
  assign N1699 = N1698 | N1690;
  assign N1700 = N1699 | N1692;
  assign N1701 = N1700 | N1648;
  assign N1702 = ~N1701;
  assign N1703 = N133 & N1634;
  assign N1704 = N834 & N1703;
  assign N1705 = N1697 | N1704;
  assign N1706 = N135 & N1634;
  assign N1707 = N834 & N1706;
  assign N1708 = N1705 | N1707;
  assign N1709 = N136 & N1634;
  assign N1710 = N1708 | N1709;
  assign N1711 = N1710 | N1648;
  assign N1712 = ~N1711;
  assign N1713 = N1636 | N1704;
  assign N1714 = N1713 | N1707;
  assign N1715 = N1714 | N1709;
  assign N1716 = N1715 | N1648;
  assign N1717 = ~N1716;

endmodule