module bsg_mux_one_hot_128_02
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [255:0] data_i;
  input [1:0] sel_one_hot_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire [255:0] data_masked;
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[128] | data_masked[0];
  assign data_o[1] = data_masked[129] | data_masked[1];
  assign data_o[2] = data_masked[130] | data_masked[2];
  assign data_o[3] = data_masked[131] | data_masked[3];
  assign data_o[4] = data_masked[132] | data_masked[4];
  assign data_o[5] = data_masked[133] | data_masked[5];
  assign data_o[6] = data_masked[134] | data_masked[6];
  assign data_o[7] = data_masked[135] | data_masked[7];
  assign data_o[8] = data_masked[136] | data_masked[8];
  assign data_o[9] = data_masked[137] | data_masked[9];
  assign data_o[10] = data_masked[138] | data_masked[10];
  assign data_o[11] = data_masked[139] | data_masked[11];
  assign data_o[12] = data_masked[140] | data_masked[12];
  assign data_o[13] = data_masked[141] | data_masked[13];
  assign data_o[14] = data_masked[142] | data_masked[14];
  assign data_o[15] = data_masked[143] | data_masked[15];
  assign data_o[16] = data_masked[144] | data_masked[16];
  assign data_o[17] = data_masked[145] | data_masked[17];
  assign data_o[18] = data_masked[146] | data_masked[18];
  assign data_o[19] = data_masked[147] | data_masked[19];
  assign data_o[20] = data_masked[148] | data_masked[20];
  assign data_o[21] = data_masked[149] | data_masked[21];
  assign data_o[22] = data_masked[150] | data_masked[22];
  assign data_o[23] = data_masked[151] | data_masked[23];
  assign data_o[24] = data_masked[152] | data_masked[24];
  assign data_o[25] = data_masked[153] | data_masked[25];
  assign data_o[26] = data_masked[154] | data_masked[26];
  assign data_o[27] = data_masked[155] | data_masked[27];
  assign data_o[28] = data_masked[156] | data_masked[28];
  assign data_o[29] = data_masked[157] | data_masked[29];
  assign data_o[30] = data_masked[158] | data_masked[30];
  assign data_o[31] = data_masked[159] | data_masked[31];
  assign data_o[32] = data_masked[160] | data_masked[32];
  assign data_o[33] = data_masked[161] | data_masked[33];
  assign data_o[34] = data_masked[162] | data_masked[34];
  assign data_o[35] = data_masked[163] | data_masked[35];
  assign data_o[36] = data_masked[164] | data_masked[36];
  assign data_o[37] = data_masked[165] | data_masked[37];
  assign data_o[38] = data_masked[166] | data_masked[38];
  assign data_o[39] = data_masked[167] | data_masked[39];
  assign data_o[40] = data_masked[168] | data_masked[40];
  assign data_o[41] = data_masked[169] | data_masked[41];
  assign data_o[42] = data_masked[170] | data_masked[42];
  assign data_o[43] = data_masked[171] | data_masked[43];
  assign data_o[44] = data_masked[172] | data_masked[44];
  assign data_o[45] = data_masked[173] | data_masked[45];
  assign data_o[46] = data_masked[174] | data_masked[46];
  assign data_o[47] = data_masked[175] | data_masked[47];
  assign data_o[48] = data_masked[176] | data_masked[48];
  assign data_o[49] = data_masked[177] | data_masked[49];
  assign data_o[50] = data_masked[178] | data_masked[50];
  assign data_o[51] = data_masked[179] | data_masked[51];
  assign data_o[52] = data_masked[180] | data_masked[52];
  assign data_o[53] = data_masked[181] | data_masked[53];
  assign data_o[54] = data_masked[182] | data_masked[54];
  assign data_o[55] = data_masked[183] | data_masked[55];
  assign data_o[56] = data_masked[184] | data_masked[56];
  assign data_o[57] = data_masked[185] | data_masked[57];
  assign data_o[58] = data_masked[186] | data_masked[58];
  assign data_o[59] = data_masked[187] | data_masked[59];
  assign data_o[60] = data_masked[188] | data_masked[60];
  assign data_o[61] = data_masked[189] | data_masked[61];
  assign data_o[62] = data_masked[190] | data_masked[62];
  assign data_o[63] = data_masked[191] | data_masked[63];
  assign data_o[64] = data_masked[192] | data_masked[64];
  assign data_o[65] = data_masked[193] | data_masked[65];
  assign data_o[66] = data_masked[194] | data_masked[66];
  assign data_o[67] = data_masked[195] | data_masked[67];
  assign data_o[68] = data_masked[196] | data_masked[68];
  assign data_o[69] = data_masked[197] | data_masked[69];
  assign data_o[70] = data_masked[198] | data_masked[70];
  assign data_o[71] = data_masked[199] | data_masked[71];
  assign data_o[72] = data_masked[200] | data_masked[72];
  assign data_o[73] = data_masked[201] | data_masked[73];
  assign data_o[74] = data_masked[202] | data_masked[74];
  assign data_o[75] = data_masked[203] | data_masked[75];
  assign data_o[76] = data_masked[204] | data_masked[76];
  assign data_o[77] = data_masked[205] | data_masked[77];
  assign data_o[78] = data_masked[206] | data_masked[78];
  assign data_o[79] = data_masked[207] | data_masked[79];
  assign data_o[80] = data_masked[208] | data_masked[80];
  assign data_o[81] = data_masked[209] | data_masked[81];
  assign data_o[82] = data_masked[210] | data_masked[82];
  assign data_o[83] = data_masked[211] | data_masked[83];
  assign data_o[84] = data_masked[212] | data_masked[84];
  assign data_o[85] = data_masked[213] | data_masked[85];
  assign data_o[86] = data_masked[214] | data_masked[86];
  assign data_o[87] = data_masked[215] | data_masked[87];
  assign data_o[88] = data_masked[216] | data_masked[88];
  assign data_o[89] = data_masked[217] | data_masked[89];
  assign data_o[90] = data_masked[218] | data_masked[90];
  assign data_o[91] = data_masked[219] | data_masked[91];
  assign data_o[92] = data_masked[220] | data_masked[92];
  assign data_o[93] = data_masked[221] | data_masked[93];
  assign data_o[94] = data_masked[222] | data_masked[94];
  assign data_o[95] = data_masked[223] | data_masked[95];
  assign data_o[96] = data_masked[224] | data_masked[96];
  assign data_o[97] = data_masked[225] | data_masked[97];
  assign data_o[98] = data_masked[226] | data_masked[98];
  assign data_o[99] = data_masked[227] | data_masked[99];
  assign data_o[100] = data_masked[228] | data_masked[100];
  assign data_o[101] = data_masked[229] | data_masked[101];
  assign data_o[102] = data_masked[230] | data_masked[102];
  assign data_o[103] = data_masked[231] | data_masked[103];
  assign data_o[104] = data_masked[232] | data_masked[104];
  assign data_o[105] = data_masked[233] | data_masked[105];
  assign data_o[106] = data_masked[234] | data_masked[106];
  assign data_o[107] = data_masked[235] | data_masked[107];
  assign data_o[108] = data_masked[236] | data_masked[108];
  assign data_o[109] = data_masked[237] | data_masked[109];
  assign data_o[110] = data_masked[238] | data_masked[110];
  assign data_o[111] = data_masked[239] | data_masked[111];
  assign data_o[112] = data_masked[240] | data_masked[112];
  assign data_o[113] = data_masked[241] | data_masked[113];
  assign data_o[114] = data_masked[242] | data_masked[114];
  assign data_o[115] = data_masked[243] | data_masked[115];
  assign data_o[116] = data_masked[244] | data_masked[116];
  assign data_o[117] = data_masked[245] | data_masked[117];
  assign data_o[118] = data_masked[246] | data_masked[118];
  assign data_o[119] = data_masked[247] | data_masked[119];
  assign data_o[120] = data_masked[248] | data_masked[120];
  assign data_o[121] = data_masked[249] | data_masked[121];
  assign data_o[122] = data_masked[250] | data_masked[122];
  assign data_o[123] = data_masked[251] | data_masked[123];
  assign data_o[124] = data_masked[252] | data_masked[124];
  assign data_o[125] = data_masked[253] | data_masked[125];
  assign data_o[126] = data_masked[254] | data_masked[126];
  assign data_o[127] = data_masked[255] | data_masked[127];

endmodule