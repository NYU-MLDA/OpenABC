module CSRFile( // @[:freechips.rocketchip.system.TinyConfig.fir@117976.2]
  input         clock, // @[:freechips.rocketchip.system.TinyConfig.fir@117977.4]
  input         reset, // @[:freechips.rocketchip.system.TinyConfig.fir@117978.4]
  input         io_ungated_clock, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_interrupts_debug, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_interrupts_mtip, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_interrupts_msip, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_interrupts_meip, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [11:0] io_rw_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [2:0]  io_rw_cmd, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_rw_rdata, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [31:0] io_rw_wdata, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [11:0] io_decode_0_csr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_decode_0_fp_illegal, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_decode_0_fp_csr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_decode_0_read_illegal, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_decode_0_write_illegal, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_decode_0_write_flush, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_csr_stall, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_eret, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_singleStep, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_debug, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_cease, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_status_isa, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_dprv, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_prv, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_sd, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [26:0] io_status_zero2, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_sxl, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_uxl, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_sd_rv32, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [7:0]  io_status_zero1, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_tsr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_tw, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_tvm, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_mxr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_sum, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_mprv, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_xs, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_fs, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_mpp, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_status_hpp, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_spp, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_mpie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_hpie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_spie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_upie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_mie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_hie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_sie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_status_uie, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_evec, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_exception, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input         io_retire, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [31:0] io_cause, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [31:0] io_pc, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [31:0] io_tval, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_time, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_interrupt, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_interrupt_cause, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_bp_0_control_action, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_bp_0_control_tmatch, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_bp_0_control_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_bp_0_control_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_bp_0_control_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_bp_0_address, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_0_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_0_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_0_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_0_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_0_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_0_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_0_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_1_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_1_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_1_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_1_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_1_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_1_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_1_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_2_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_2_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_2_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_2_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_2_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_2_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_2_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_3_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_3_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_3_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_3_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_3_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_3_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_3_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_4_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_4_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_4_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_4_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_4_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_4_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_4_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_5_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_5_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_5_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_5_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_5_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_5_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_5_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_6_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_6_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_6_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_6_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_6_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_6_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_6_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_7_cfg_l, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [1:0]  io_pmp_7_cfg_a, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_7_cfg_x, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_7_cfg_w, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_pmp_7_cfg_r, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [29:0] io_pmp_7_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_pmp_7_mask, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  input  [31:0] io_inst_0, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_trace_0_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_trace_0_iaddr, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output [31:0] io_trace_0_insn, // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
  output        io_trace_0_exception // @[:freechips.rocketchip.system.TinyConfig.fir@117979.4]
);
  reg  reg_mstatus_spp; // @[CSR.scala 238:24:freechips.rocketchip.system.TinyConfig.fir@118054.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 238:24:freechips.rocketchip.system.TinyConfig.fir@118054.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 238:24:freechips.rocketchip.system.TinyConfig.fir@118054.4]
  reg [31:0] _RAND_2;
  reg  reg_dcsr_ebreakm; // @[CSR.scala 246:21:freechips.rocketchip.system.TinyConfig.fir@118097.4]
  reg [31:0] _RAND_3;
  reg [2:0] reg_dcsr_cause; // @[CSR.scala 246:21:freechips.rocketchip.system.TinyConfig.fir@118097.4]
  reg [31:0] _RAND_4;
  reg  reg_dcsr_step; // @[CSR.scala 246:21:freechips.rocketchip.system.TinyConfig.fir@118097.4]
  reg [31:0] _RAND_5;
  reg  reg_debug; // @[CSR.scala 287:22:freechips.rocketchip.system.TinyConfig.fir@118153.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_dpc; // @[CSR.scala 288:20:freechips.rocketchip.system.TinyConfig.fir@118154.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_dscratch; // @[CSR.scala 289:25:freechips.rocketchip.system.TinyConfig.fir@118155.4]
  reg [31:0] _RAND_8;
  reg  reg_singleStepped; // @[CSR.scala 290:30:freechips.rocketchip.system.TinyConfig.fir@118156.4]
  reg [31:0] _RAND_9;
  reg  reg_bp_0_control_dmode; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_10;
  reg  reg_bp_0_control_action; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_11;
  reg [1:0] reg_bp_0_control_tmatch; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_12;
  reg  reg_bp_0_control_x; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_13;
  reg  reg_bp_0_control_w; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_14;
  reg  reg_bp_0_control_r; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_15;
  reg [31:0] reg_bp_0_address; // @[CSR.scala 293:19:freechips.rocketchip.system.TinyConfig.fir@118158.4]
  reg [31:0] _RAND_16;
  reg  reg_pmp_0_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_17;
  reg [1:0] reg_pmp_0_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_18;
  reg  reg_pmp_0_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_19;
  reg  reg_pmp_0_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_20;
  reg  reg_pmp_0_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_21;
  reg [29:0] reg_pmp_0_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_22;
  reg  reg_pmp_1_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_23;
  reg [1:0] reg_pmp_1_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_24;
  reg  reg_pmp_1_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_25;
  reg  reg_pmp_1_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_26;
  reg  reg_pmp_1_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_27;
  reg [29:0] reg_pmp_1_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_28;
  reg  reg_pmp_2_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_29;
  reg [1:0] reg_pmp_2_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_30;
  reg  reg_pmp_2_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_31;
  reg  reg_pmp_2_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_32;
  reg  reg_pmp_2_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_33;
  reg [29:0] reg_pmp_2_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_34;
  reg  reg_pmp_3_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_35;
  reg [1:0] reg_pmp_3_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_36;
  reg  reg_pmp_3_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_37;
  reg  reg_pmp_3_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_38;
  reg  reg_pmp_3_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_39;
  reg [29:0] reg_pmp_3_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_40;
  reg  reg_pmp_4_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_41;
  reg [1:0] reg_pmp_4_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_42;
  reg  reg_pmp_4_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_43;
  reg  reg_pmp_4_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_44;
  reg  reg_pmp_4_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_45;
  reg [29:0] reg_pmp_4_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_46;
  reg  reg_pmp_5_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_47;
  reg [1:0] reg_pmp_5_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_48;
  reg  reg_pmp_5_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_49;
  reg  reg_pmp_5_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_50;
  reg  reg_pmp_5_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_51;
  reg [29:0] reg_pmp_5_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_52;
  reg  reg_pmp_6_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_53;
  reg [1:0] reg_pmp_6_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_54;
  reg  reg_pmp_6_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_55;
  reg  reg_pmp_6_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_56;
  reg  reg_pmp_6_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_57;
  reg [29:0] reg_pmp_6_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_58;
  reg  reg_pmp_7_cfg_l; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_59;
  reg [1:0] reg_pmp_7_cfg_a; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_60;
  reg  reg_pmp_7_cfg_x; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_61;
  reg  reg_pmp_7_cfg_w; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_62;
  reg  reg_pmp_7_cfg_r; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_63;
  reg [29:0] reg_pmp_7_addr; // @[CSR.scala 294:20:freechips.rocketchip.system.TinyConfig.fir@118159.4]
  reg [31:0] _RAND_64;
  reg [31:0] reg_mie; // @[CSR.scala 296:20:freechips.rocketchip.system.TinyConfig.fir@118160.4]
  reg [31:0] _RAND_65;
  reg [31:0] reg_mepc; // @[CSR.scala 306:21:freechips.rocketchip.system.TinyConfig.fir@118168.4]
  reg [31:0] _RAND_66;
  reg [31:0] reg_mcause; // @[CSR.scala 307:23:freechips.rocketchip.system.TinyConfig.fir@118169.4]
  reg [31:0] _RAND_67;
  reg [31:0] reg_mtval; // @[CSR.scala 308:22:freechips.rocketchip.system.TinyConfig.fir@118170.4]
  reg [31:0] _RAND_68;
  reg [31:0] reg_mscratch; // @[CSR.scala 309:25:freechips.rocketchip.system.TinyConfig.fir@118171.4]
  reg [31:0] _RAND_69;
  reg [31:0] reg_mtvec; // @[CSR.scala 312:27:freechips.rocketchip.system.TinyConfig.fir@118172.4]
  reg [31:0] _RAND_70;
  reg  reg_wfi; // @[CSR.scala 332:50:freechips.rocketchip.system.TinyConfig.fir@118185.4]
  reg [31:0] _RAND_71;
  reg [5:0] _T_83; // @[Counters.scala 46:37:freechips.rocketchip.system.TinyConfig.fir@118188.4]
  reg [31:0] _RAND_72;
  wire [5:0] _GEN_415; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118189.4]
  wire [6:0] _T_84; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118189.4]
  reg [57:0] _T_85; // @[Counters.scala 51:27:freechips.rocketchip.system.TinyConfig.fir@118191.4]
  reg [63:0] _RAND_73;
  wire  _T_86; // @[Counters.scala 52:20:freechips.rocketchip.system.TinyConfig.fir@118192.4]
  wire [57:0] _T_88; // @[Counters.scala 52:43:freechips.rocketchip.system.TinyConfig.fir@118195.6]
  wire [63:0] _T_89; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118198.4]
  wire  _T_90; // @[CSR.scala 338:103:freechips.rocketchip.system.TinyConfig.fir@118199.4]
  reg [5:0] _T_91; // @[Counters.scala 46:37:freechips.rocketchip.system.TinyConfig.fir@118200.4]
  reg [31:0] _RAND_74;
  wire [5:0] _GEN_416; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118201.4]
  wire [6:0] _T_92; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118201.4]
  reg [57:0] _T_93; // @[Counters.scala 51:27:freechips.rocketchip.system.TinyConfig.fir@118203.4]
  reg [63:0] _RAND_75;
  wire  _T_94; // @[Counters.scala 52:20:freechips.rocketchip.system.TinyConfig.fir@118204.4]
  wire [57:0] _T_96; // @[Counters.scala 52:43:freechips.rocketchip.system.TinyConfig.fir@118207.6]
  wire [63:0] _T_97; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118210.4]
  wire [15:0] _T_112; // @[CSR.scala 351:22:freechips.rocketchip.system.TinyConfig.fir@118232.4]
  wire [15:0] read_mip; // @[CSR.scala 351:29:freechips.rocketchip.system.TinyConfig.fir@118233.4]
  wire [31:0] _GEN_417; // @[CSR.scala 354:56:freechips.rocketchip.system.TinyConfig.fir@118234.4]
  wire [31:0] pending_interrupts; // @[CSR.scala 354:56:freechips.rocketchip.system.TinyConfig.fir@118234.4]
  wire [14:0] d_interrupts; // @[CSR.scala 355:42:freechips.rocketchip.system.TinyConfig.fir@118236.4]
  wire [31:0] _T_116; // @[CSR.scala 356:73:freechips.rocketchip.system.TinyConfig.fir@118239.4]
  wire [31:0] _T_118; // @[CSR.scala 356:71:freechips.rocketchip.system.TinyConfig.fir@118241.4]
  wire [31:0] m_interrupts; // @[CSR.scala 356:25:freechips.rocketchip.system.TinyConfig.fir@118242.4]
  wire  _T_124; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118249.4]
  wire  _T_125; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118250.4]
  wire  _T_126; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118251.4]
  wire  _T_127; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118252.4]
  wire  _T_128; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118253.4]
  wire  _T_129; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118254.4]
  wire  _T_130; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118255.4]
  wire  _T_131; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118256.4]
  wire  _T_132; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118257.4]
  wire  _T_133; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118258.4]
  wire  _T_134; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118259.4]
  wire  _T_135; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118260.4]
  wire  _T_136; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118261.4]
  wire  _T_137; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118262.4]
  wire  _T_138; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118263.4]
  wire  _T_139; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118264.4]
  wire  _T_140; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118265.4]
  wire  _T_141; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118266.4]
  wire  _T_142; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118267.4]
  wire  _T_143; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118268.4]
  wire  _T_144; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118269.4]
  wire  _T_145; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118270.4]
  wire  _T_146; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118271.4]
  wire  _T_147; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118272.4]
  wire  _T_148; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118273.4]
  wire  _T_162; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118287.4]
  wire  _T_163; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118288.4]
  wire  _T_164; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118289.4]
  wire  _T_165; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118290.4]
  wire  _T_166; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118291.4]
  wire  _T_167; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118292.4]
  wire  _T_168; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118293.4]
  wire  _T_169; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118294.4]
  wire  _T_170; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118295.4]
  wire  _T_171; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118296.4]
  wire  _T_172; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118297.4]
  wire  _T_173; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118298.4]
  wire  _T_174; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118299.4]
  wire  _T_175; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118300.4]
  wire  _T_176; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118301.4]
  wire  _T_177; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118302.4]
  wire  _T_178; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118303.4]
  wire  _T_179; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118304.4]
  wire  _T_180; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118305.4]
  wire  _T_181; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118306.4]
  wire  _T_182; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118307.4]
  wire  _T_183; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118308.4]
  wire  _T_184; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118309.4]
  wire  anyInterrupt; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118310.4]
  wire [3:0] _T_249; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118375.4]
  wire [3:0] _T_250; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118376.4]
  wire [3:0] _T_251; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118377.4]
  wire [3:0] _T_252; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118378.4]
  wire [3:0] _T_253; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118379.4]
  wire [3:0] _T_254; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118380.4]
  wire [3:0] _T_255; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118381.4]
  wire [3:0] _T_256; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118382.4]
  wire [3:0] _T_257; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118383.4]
  wire [3:0] _T_258; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118384.4]
  wire [3:0] _T_259; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118385.4]
  wire [3:0] _T_260; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118386.4]
  wire [3:0] _T_261; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118387.4]
  wire [3:0] _T_262; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118388.4]
  wire [3:0] _T_263; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118389.4]
  wire [3:0] _T_264; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118390.4]
  wire [3:0] _T_265; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118391.4]
  wire [3:0] _T_266; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118392.4]
  wire [3:0] _T_267; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118393.4]
  wire [3:0] _T_268; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118394.4]
  wire [3:0] _T_269; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118395.4]
  wire [3:0] _T_270; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118396.4]
  wire [3:0] _T_271; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118397.4]
  wire [3:0] whichInterrupt; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118398.4]
  wire [31:0] _GEN_418; // @[CSR.scala 360:43:freechips.rocketchip.system.TinyConfig.fir@118399.4]
  wire  _T_273; // @[CSR.scala 361:36:freechips.rocketchip.system.TinyConfig.fir@118401.4]
  wire  _T_274; // @[CSR.scala 361:33:freechips.rocketchip.system.TinyConfig.fir@118402.4]
  wire  _T_275; // @[CSR.scala 361:51:freechips.rocketchip.system.TinyConfig.fir@118403.4]
  wire  _T_276; // @[CSR.scala 361:88:freechips.rocketchip.system.TinyConfig.fir@118404.4]
  wire  _T_277; // @[CSR.scala 361:76:freechips.rocketchip.system.TinyConfig.fir@118405.4]
  wire  _T_280; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118413.4]
  wire [30:0] _T_281; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118414.4]
  wire [30:0] _T_284; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118417.4]
  wire [30:0] _T_285; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118418.4]
  wire [30:0] _T_286; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118419.4]
  wire [32:0] _T_287; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118420.4]
  wire  _T_289; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118425.4]
  wire [30:0] _T_290; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118426.4]
  wire [30:0] _T_293; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118429.4]
  wire [30:0] _T_294; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118430.4]
  wire [30:0] _T_295; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118431.4]
  wire [32:0] _T_296; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118432.4]
  wire  _T_298; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118437.4]
  wire [30:0] _T_299; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118438.4]
  wire [30:0] _T_302; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118441.4]
  wire [30:0] _T_303; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118442.4]
  wire [30:0] _T_304; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118443.4]
  wire [32:0] _T_305; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118444.4]
  wire  _T_307; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118449.4]
  wire [30:0] _T_308; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118450.4]
  wire [30:0] _T_311; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118453.4]
  wire [30:0] _T_312; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118454.4]
  wire [30:0] _T_313; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118455.4]
  wire [32:0] _T_314; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118456.4]
  wire  _T_316; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118461.4]
  wire [30:0] _T_317; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118462.4]
  wire [30:0] _T_320; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118465.4]
  wire [30:0] _T_321; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118466.4]
  wire [30:0] _T_322; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118467.4]
  wire [32:0] _T_323; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118468.4]
  wire  _T_325; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118473.4]
  wire [30:0] _T_326; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118474.4]
  wire [30:0] _T_329; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118477.4]
  wire [30:0] _T_330; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118478.4]
  wire [30:0] _T_331; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118479.4]
  wire [32:0] _T_332; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118480.4]
  wire  _T_334; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118485.4]
  wire [30:0] _T_335; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118486.4]
  wire [30:0] _T_338; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118489.4]
  wire [30:0] _T_339; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118490.4]
  wire [30:0] _T_340; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118491.4]
  wire [32:0] _T_341; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118492.4]
  wire  _T_343; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118497.4]
  wire [30:0] _T_344; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118498.4]
  wire [30:0] _T_347; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118501.4]
  wire [30:0] _T_348; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118502.4]
  wire [30:0] _T_349; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118503.4]
  wire [32:0] _T_350; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118504.4]
  reg [31:0] reg_misa; // @[CSR.scala 378:21:freechips.rocketchip.system.TinyConfig.fir@118514.4]
  reg [31:0] _RAND_76;
  wire [6:0] _T_356; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118520.4]
  wire [18:0] _T_364; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118528.4]
  wire [14:0] _T_370; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118534.4]
  wire [101:0] _T_379; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118543.4]
  wire [31:0] read_mstatus; // @[CSR.scala 379:40:freechips.rocketchip.system.TinyConfig.fir@118544.4]
  wire  _T_380; // @[CSR.scala 936:41:freechips.rocketchip.system.TinyConfig.fir@118545.4]
  wire [6:0] _T_381; // @[CSR.scala 936:39:freechips.rocketchip.system.TinyConfig.fir@118546.4]
  wire [31:0] _T_383; // @[package.scala 131:41:freechips.rocketchip.system.TinyConfig.fir@118548.4]
  wire [31:0] _T_384; // @[package.scala 131:37:freechips.rocketchip.system.TinyConfig.fir@118549.4]
  wire [31:0] read_mtvec; // @[package.scala 131:35:freechips.rocketchip.system.TinyConfig.fir@118550.4]
  wire [6:0] _T_395; // @[CSR.scala 385:48:freechips.rocketchip.system.TinyConfig.fir@118562.4]
  wire [31:0] _T_403; // @[CSR.scala 385:48:freechips.rocketchip.system.TinyConfig.fir@118570.4]
  wire [31:0] _T_404; // @[CSR.scala 935:28:freechips.rocketchip.system.TinyConfig.fir@118571.4]
  wire  _T_405; // @[CSR.scala 935:45:freechips.rocketchip.system.TinyConfig.fir@118572.4]
  wire [1:0] _T_406; // @[CSR.scala 935:36:freechips.rocketchip.system.TinyConfig.fir@118573.4]
  wire [31:0] _GEN_419; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118574.4]
  wire [31:0] _T_407; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118574.4]
  wire [31:0] _T_408; // @[CSR.scala 935:26:freechips.rocketchip.system.TinyConfig.fir@118575.4]
  wire [31:0] _T_421; // @[CSR.scala 399:27:freechips.rocketchip.system.TinyConfig.fir@118588.4]
  wire [31:0] _T_422; // @[CSR.scala 935:28:freechips.rocketchip.system.TinyConfig.fir@118589.4]
  wire [31:0] _T_425; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118592.4]
  wire [31:0] _T_426; // @[CSR.scala 935:26:freechips.rocketchip.system.TinyConfig.fir@118593.4]
  wire [31:0] _T_457; // @[CSR.scala 436:50:freechips.rocketchip.system.TinyConfig.fir@118624.4]
  wire [31:0] _T_458; // @[CSR.scala 437:54:freechips.rocketchip.system.TinyConfig.fir@118625.4]
  wire [7:0] _T_473; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118651.4]
  wire [7:0] _T_483; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118661.4]
  wire [15:0] _T_489; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118667.4]
  wire [31:0] _T_491; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118669.4]
  wire [7:0] _T_496; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118674.4]
  wire [7:0] _T_506; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118684.4]
  wire [15:0] _T_512; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118690.4]
  wire [31:0] _T_514; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118692.4]
  wire  _T_562; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118744.4]
  wire  _T_563; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118745.4]
  wire  _T_564; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118746.4]
  wire  _T_565; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118747.4]
  wire  _T_566; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118748.4]
  wire  _T_567; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118749.4]
  wire  _T_568; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118750.4]
  wire  _T_569; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118751.4]
  wire  _T_570; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118752.4]
  wire  _T_571; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118753.4]
  wire  _T_572; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118754.4]
  wire  _T_574; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118756.4]
  wire  _T_575; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118757.4]
  wire  _T_576; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118758.4]
  wire  _T_577; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118759.4]
  wire  _T_578; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118760.4]
  wire  _T_666; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118848.4]
  wire  _T_667; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118849.4]
  wire  _T_668; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118850.4]
  wire  _T_669; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118851.4]
  wire  _T_672; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118854.4]
  wire  _T_673; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118855.4]
  wire  _T_674; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118856.4]
  wire  _T_675; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118857.4]
  wire  _T_676; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118858.4]
  wire  _T_677; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118859.4]
  wire  _T_678; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118860.4]
  wire  _T_679; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118861.4]
  wire  _T_689; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118871.4]
  wire  _T_691; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118873.4]
  wire  _T_692; // @[CSR.scala 913:13:freechips.rocketchip.system.TinyConfig.fir@118874.4]
  wire [31:0] _T_693; // @[CSR.scala 913:9:freechips.rocketchip.system.TinyConfig.fir@118875.4]
  wire [31:0] _T_694; // @[CSR.scala 913:34:freechips.rocketchip.system.TinyConfig.fir@118876.4]
  wire [1:0] _T_695; // @[CSR.scala 913:53:freechips.rocketchip.system.TinyConfig.fir@118877.4]
  wire  _T_696; // @[CSR.scala 913:59:freechips.rocketchip.system.TinyConfig.fir@118878.4]
  wire [31:0] _T_697; // @[CSR.scala 913:49:freechips.rocketchip.system.TinyConfig.fir@118879.4]
  wire [31:0] _T_698; // @[CSR.scala 913:45:freechips.rocketchip.system.TinyConfig.fir@118880.4]
  wire [31:0] wdata; // @[CSR.scala 913:43:freechips.rocketchip.system.TinyConfig.fir@118881.4]
  wire  system_insn; // @[CSR.scala 500:31:freechips.rocketchip.system.TinyConfig.fir@118882.4]
  wire [31:0] _T_699; // @[CSR.scala 512:28:freechips.rocketchip.system.TinyConfig.fir@118883.4]
  wire [31:0] _T_700; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118884.4]
  wire  _T_701; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118885.4]
  wire [31:0] _T_703; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118887.4]
  wire  _T_704; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118888.4]
  wire [31:0] _T_706; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118890.4]
  wire  _T_707; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118891.4]
  wire [31:0] _T_709; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118893.4]
  wire  _T_710; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118894.4]
  wire [31:0] _T_712; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118896.4]
  wire  _T_713; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118897.4]
  wire  insn_call; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118900.4]
  wire  insn_break; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118902.4]
  wire  insn_ret; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118904.4]
  wire  insn_cease; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118906.4]
  wire  insn_wfi; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118908.4]
  wire  _T_764; // @[CSR.scala 524:39:freechips.rocketchip.system.TinyConfig.fir@118954.4]
  wire  _T_765; // @[CSR.scala 524:57:freechips.rocketchip.system.TinyConfig.fir@118955.4]
  wire  _T_766; // @[CSR.scala 524:48:freechips.rocketchip.system.TinyConfig.fir@118956.4]
  wire  _T_779; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118972.4]
  wire  _T_780; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118973.4]
  wire  _T_781; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118974.4]
  wire  _T_782; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118975.4]
  wire  _T_783; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118976.4]
  wire  _T_784; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118977.4]
  wire  _T_785; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118978.4]
  wire  _T_786; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118979.4]
  wire  _T_787; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118980.4]
  wire  _T_788; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118981.4]
  wire  _T_789; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118982.4]
  wire  _T_790; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118983.4]
  wire  _T_791; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118984.4]
  wire  _T_792; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118985.4]
  wire  _T_793; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118986.4]
  wire  _T_794; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118987.4]
  wire  _T_795; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118988.4]
  wire  _T_796; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118989.4]
  wire  _T_797; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118990.4]
  wire  _T_798; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118991.4]
  wire  _T_799; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118992.4]
  wire  _T_800; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118993.4]
  wire  _T_801; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118994.4]
  wire  _T_802; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118995.4]
  wire  _T_803; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118996.4]
  wire  _T_804; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118997.4]
  wire  _T_805; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118998.4]
  wire  _T_806; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118999.4]
  wire  _T_807; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119000.4]
  wire  _T_808; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119001.4]
  wire  _T_809; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119002.4]
  wire  _T_810; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119003.4]
  wire  _T_811; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119004.4]
  wire  _T_812; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119005.4]
  wire  _T_813; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119006.4]
  wire  _T_814; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119007.4]
  wire  _T_815; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119008.4]
  wire  _T_816; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119009.4]
  wire  _T_817; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119010.4]
  wire  _T_818; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119011.4]
  wire  _T_819; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119012.4]
  wire  _T_820; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119013.4]
  wire  _T_821; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119014.4]
  wire  _T_822; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119015.4]
  wire  _T_823; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119016.4]
  wire  _T_824; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119017.4]
  wire  _T_825; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119018.4]
  wire  _T_826; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119019.4]
  wire  _T_827; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119020.4]
  wire  _T_828; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119021.4]
  wire  _T_829; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119022.4]
  wire  _T_830; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119023.4]
  wire  _T_831; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119024.4]
  wire  _T_832; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119025.4]
  wire  _T_833; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119026.4]
  wire  _T_834; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119027.4]
  wire  _T_835; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119028.4]
  wire  _T_836; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119029.4]
  wire  _T_837; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119030.4]
  wire  _T_838; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119031.4]
  wire  _T_839; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119032.4]
  wire  _T_840; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119033.4]
  wire  _T_841; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119034.4]
  wire  _T_842; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119035.4]
  wire  _T_843; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119036.4]
  wire  _T_844; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119037.4]
  wire  _T_845; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119038.4]
  wire  _T_846; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119039.4]
  wire  _T_847; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119040.4]
  wire  _T_848; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119041.4]
  wire  _T_849; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119042.4]
  wire  _T_850; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119043.4]
  wire  _T_851; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119044.4]
  wire  _T_852; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119045.4]
  wire  _T_853; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119046.4]
  wire  _T_854; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119047.4]
  wire  _T_855; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119048.4]
  wire  _T_856; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119049.4]
  wire  _T_857; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119050.4]
  wire  _T_858; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119051.4]
  wire  _T_859; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119052.4]
  wire  _T_860; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119053.4]
  wire  _T_861; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119054.4]
  wire  _T_862; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119055.4]
  wire  _T_863; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119056.4]
  wire  _T_864; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119057.4]
  wire  _T_865; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119058.4]
  wire  _T_866; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119059.4]
  wire  _T_867; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119060.4]
  wire  _T_868; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119061.4]
  wire  _T_869; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119062.4]
  wire  _T_870; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119063.4]
  wire  _T_871; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119064.4]
  wire  _T_872; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119065.4]
  wire  _T_873; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119066.4]
  wire  _T_874; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119067.4]
  wire  _T_875; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119068.4]
  wire  _T_876; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119069.4]
  wire  _T_877; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119070.4]
  wire  _T_878; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119071.4]
  wire  _T_879; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119072.4]
  wire  _T_880; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119073.4]
  wire  _T_881; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119074.4]
  wire  _T_882; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119075.4]
  wire  _T_883; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119076.4]
  wire  _T_884; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119077.4]
  wire  _T_885; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119078.4]
  wire  _T_886; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119079.4]
  wire  _T_887; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119080.4]
  wire  _T_888; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119081.4]
  wire  _T_889; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119082.4]
  wire  _T_890; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119083.4]
  wire  _T_891; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119084.4]
  wire  _T_892; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119085.4]
  wire  _T_893; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119086.4]
  wire  _T_894; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119087.4]
  wire  _T_895; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119088.4]
  wire  _T_896; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119089.4]
  wire  _T_897; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119090.4]
  wire  _T_898; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119091.4]
  wire  _T_899; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119092.4]
  wire  _T_900; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119093.4]
  wire  _T_901; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119094.4]
  wire  _T_902; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119095.4]
  wire  _T_903; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119096.4]
  wire  _T_904; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119097.4]
  wire  _T_905; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119098.4]
  wire  _T_906; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119099.4]
  wire  _T_907; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119100.4]
  wire  _T_908; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119101.4]
  wire  _T_909; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119102.4]
  wire  _T_910; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119103.4]
  wire  _T_911; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119104.4]
  wire  _T_912; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119105.4]
  wire  _T_913; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119106.4]
  wire  _T_914; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119107.4]
  wire  _T_915; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119108.4]
  wire  _T_916; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119109.4]
  wire  _T_917; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119110.4]
  wire  _T_918; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119111.4]
  wire  _T_919; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119112.4]
  wire  _T_920; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119113.4]
  wire  _T_921; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119114.4]
  wire  _T_922; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119115.4]
  wire  _T_923; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119116.4]
  wire  _T_924; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119117.4]
  wire  _T_925; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119118.4]
  wire  _T_926; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119119.4]
  wire  _T_927; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119120.4]
  wire  _T_928; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119121.4]
  wire  _T_929; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119122.4]
  wire  _T_930; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119123.4]
  wire  _T_931; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119124.4]
  wire  _T_932; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119125.4]
  wire  _T_933; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119126.4]
  wire  _T_934; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119127.4]
  wire  _T_935; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119128.4]
  wire  _T_936; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119129.4]
  wire  _T_937; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119130.4]
  wire  _T_938; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119131.4]
  wire  _T_939; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119132.4]
  wire  _T_940; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119133.4]
  wire  _T_941; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119134.4]
  wire  _T_942; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119135.4]
  wire  _T_943; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119136.4]
  wire  _T_944; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119137.4]
  wire  _T_945; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119138.4]
  wire  _T_946; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119139.4]
  wire  _T_947; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119140.4]
  wire  _T_948; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119141.4]
  wire  _T_949; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119142.4]
  wire  _T_950; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119143.4]
  wire  _T_951; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119144.4]
  wire  _T_952; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119145.4]
  wire  _T_953; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119146.4]
  wire  _T_954; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119147.4]
  wire  _T_955; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119148.4]
  wire  _T_956; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119149.4]
  wire  _T_957; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119150.4]
  wire  _T_958; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119151.4]
  wire  _T_959; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119152.4]
  wire  _T_960; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119153.4]
  wire  _T_961; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119154.4]
  wire  _T_962; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119155.4]
  wire  _T_963; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119156.4]
  wire  _T_964; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119157.4]
  wire  _T_965; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119158.4]
  wire  _T_966; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119159.4]
  wire  _T_967; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119160.4]
  wire  _T_968; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119161.4]
  wire  _T_969; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119162.4]
  wire  _T_970; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119163.4]
  wire  _T_971; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119164.4]
  wire  _T_972; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119165.4]
  wire  _T_973; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119166.4]
  wire  _T_974; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119167.4]
  wire  _T_975; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119168.4]
  wire  _T_976; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119169.4]
  wire  _T_977; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119170.4]
  wire  _T_978; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119171.4]
  wire  _T_979; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119172.4]
  wire  _T_980; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119173.4]
  wire  _T_981; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119174.4]
  wire  _T_982; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119175.4]
  wire  _T_983; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119176.4]
  wire  _T_984; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119177.4]
  wire  _T_985; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119178.4]
  wire  _T_986; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119179.4]
  wire  _T_987; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119180.4]
  wire  _T_988; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119181.4]
  wire  _T_989; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119182.4]
  wire  _T_990; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119183.4]
  wire  _T_991; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119184.4]
  wire  _T_992; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119185.4]
  wire  _T_993; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119186.4]
  wire  _T_994; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119187.4]
  wire  _T_995; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119188.4]
  wire  _T_996; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119189.4]
  wire  _T_997; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119190.4]
  wire  _T_998; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119191.4]
  wire  _T_999; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119192.4]
  wire  _T_1000; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119193.4]
  wire  _T_1001; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119194.4]
  wire  _T_1002; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119195.4]
  wire  _T_1003; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119196.4]
  wire  _T_1004; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119197.4]
  wire  _T_1005; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119198.4]
  wire  _T_1006; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119199.4]
  wire  _T_1007; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119200.4]
  wire  _T_1008; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119201.4]
  wire  _T_1009; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119202.4]
  wire  _T_1010; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119203.4]
  wire  _T_1011; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119204.4]
  wire  _T_1012; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119205.4]
  wire  _T_1013; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119206.4]
  wire  _T_1014; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119207.4]
  wire  _T_1015; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119208.4]
  wire  _T_1016; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119209.4]
  wire  _T_1017; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119210.4]
  wire  _T_1018; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119211.4]
  wire  _T_1019; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119212.4]
  wire  _T_1020; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119213.4]
  wire  _T_1021; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119214.4]
  wire  _T_1022; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119215.4]
  wire  _T_1023; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119216.4]
  wire  _T_1024; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119217.4]
  wire  _T_1025; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119218.4]
  wire  _T_1026; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119219.4]
  wire  _T_1027; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119220.4]
  wire  _T_1028; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119221.4]
  wire  _T_1029; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119222.4]
  wire  _T_1030; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119223.4]
  wire  _T_1031; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119224.4]
  wire  _T_1032; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119225.4]
  wire  _T_1033; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119226.4]
  wire  _T_1034; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119227.4]
  wire  _T_1035; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119228.4]
  wire  _T_1036; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119229.4]
  wire  _T_1037; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119230.4]
  wire  _T_1038; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119231.4]
  wire  _T_1039; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119232.4]
  wire  _T_1040; // @[CSR.scala 528:7:freechips.rocketchip.system.TinyConfig.fir@119233.4]
  wire  _T_1059; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119252.4]
  wire  _T_1060; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119253.4]
  wire  _T_1062; // @[CSR.scala 531:52:freechips.rocketchip.system.TinyConfig.fir@119255.4]
  wire  _T_1063; // @[CSR.scala 531:49:freechips.rocketchip.system.TinyConfig.fir@119256.4]
  wire  _T_1064; // @[CSR.scala 530:148:freechips.rocketchip.system.TinyConfig.fir@119257.4]
  wire  _T_1065; // @[CSR.scala 532:21:freechips.rocketchip.system.TinyConfig.fir@119258.4]
  wire [1:0] _T_1067; // @[CSR.scala 533:39:freechips.rocketchip.system.TinyConfig.fir@119261.4]
  wire  _T_1069; // @[CSR.scala 534:40:freechips.rocketchip.system.TinyConfig.fir@119264.4]
  wire  _T_1070; // @[CSR.scala 534:71:freechips.rocketchip.system.TinyConfig.fir@119265.4]
  wire  _T_1071; // @[CSR.scala 534:57:freechips.rocketchip.system.TinyConfig.fir@119266.4]
  wire  _T_1072; // @[CSR.scala 534:99:freechips.rocketchip.system.TinyConfig.fir@119267.4]
  wire  _T_1073; // @[CSR.scala 534:130:freechips.rocketchip.system.TinyConfig.fir@119268.4]
  wire  _T_1074; // @[CSR.scala 534:116:freechips.rocketchip.system.TinyConfig.fir@119269.4]
  wire  _T_1075; // @[CSR.scala 534:85:freechips.rocketchip.system.TinyConfig.fir@119270.4]
  wire [31:0] _T_1090; // @[CSR.scala 543:14:freechips.rocketchip.system.TinyConfig.fir@119287.4]
  wire [31:0] cause; // @[CSR.scala 542:8:freechips.rocketchip.system.TinyConfig.fir@119288.4]
  wire [7:0] cause_lsbs; // @[CSR.scala 544:25:freechips.rocketchip.system.TinyConfig.fir@119289.4]
  wire  _T_1091; // @[CSR.scala 545:30:freechips.rocketchip.system.TinyConfig.fir@119290.4]
  wire  _T_1092; // @[CSR.scala 545:53:freechips.rocketchip.system.TinyConfig.fir@119291.4]
  wire  causeIsDebugInt; // @[CSR.scala 545:39:freechips.rocketchip.system.TinyConfig.fir@119292.4]
  wire  _T_1094; // @[CSR.scala 546:29:freechips.rocketchip.system.TinyConfig.fir@119294.4]
  wire  causeIsDebugTrigger; // @[CSR.scala 546:44:freechips.rocketchip.system.TinyConfig.fir@119296.4]
  wire  _T_1098; // @[CSR.scala 547:42:freechips.rocketchip.system.TinyConfig.fir@119299.4]
  wire [3:0] _T_1101; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@119302.4]
  wire  _GEN_421; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119303.4]
  wire [3:0] _T_1102; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119303.4]
  wire  _T_1103; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119304.4]
  wire  causeIsDebugBreak; // @[CSR.scala 547:56:freechips.rocketchip.system.TinyConfig.fir@119305.4]
  wire  _T_1104; // @[CSR.scala 548:60:freechips.rocketchip.system.TinyConfig.fir@119306.4]
  wire  _T_1105; // @[CSR.scala 548:79:freechips.rocketchip.system.TinyConfig.fir@119307.4]
  wire  _T_1106; // @[CSR.scala 548:102:freechips.rocketchip.system.TinyConfig.fir@119308.4]
  wire  trapToDebug; // @[CSR.scala 548:123:freechips.rocketchip.system.TinyConfig.fir@119309.4]
  wire [11:0] _T_1108; // @[CSR.scala 549:37:freechips.rocketchip.system.TinyConfig.fir@119311.4]
  wire [11:0] debugTVec; // @[CSR.scala 549:22:freechips.rocketchip.system.TinyConfig.fir@119312.4]
  wire [4:0] _T_1118; // @[CSR.scala 558:32:freechips.rocketchip.system.TinyConfig.fir@119323.4]
  wire [6:0] _T_1119; // @[CSR.scala 558:59:freechips.rocketchip.system.TinyConfig.fir@119324.4]
  wire [24:0] _T_1120; // @[CSR.scala 559:33:freechips.rocketchip.system.TinyConfig.fir@119325.4]
  wire [31:0] _T_1121; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@119326.4]
  wire  _T_1122; // @[CSR.scala 560:24:freechips.rocketchip.system.TinyConfig.fir@119327.4]
  wire  _T_1124; // @[CSR.scala 560:28:freechips.rocketchip.system.TinyConfig.fir@119329.4]
  wire [2:0] _T_1125; // @[CSR.scala 560:70:freechips.rocketchip.system.TinyConfig.fir@119330.4]
  wire  _T_1126; // @[CSR.scala 560:94:freechips.rocketchip.system.TinyConfig.fir@119331.4]
  wire  _T_1127; // @[CSR.scala 560:55:freechips.rocketchip.system.TinyConfig.fir@119332.4]
  wire [29:0] _T_1128; // @[CSR.scala 561:38:freechips.rocketchip.system.TinyConfig.fir@119333.4]
  wire [31:0] _T_1129; // @[CSR.scala 561:56:freechips.rocketchip.system.TinyConfig.fir@119334.4]
  wire [31:0] notDebugTVec; // @[CSR.scala 561:8:freechips.rocketchip.system.TinyConfig.fir@119335.4]
  wire [31:0] tvec; // @[CSR.scala 563:17:freechips.rocketchip.system.TinyConfig.fir@119336.4]
  wire  _T_1130; // @[CSR.scala 566:24:freechips.rocketchip.system.TinyConfig.fir@119339.4]
  wire  _T_1134; // @[CSR.scala 569:32:freechips.rocketchip.system.TinyConfig.fir@119346.4]
  wire  _T_1135; // @[CSR.scala 569:53:freechips.rocketchip.system.TinyConfig.fir@119347.4]
  wire  exception; // @[CSR.scala 578:43:freechips.rocketchip.system.TinyConfig.fir@119362.4]
  wire [1:0] _T_1142; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119363.4]
  wire [1:0] _T_1144; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119365.4]
  wire [2:0] _T_1146; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119367.4]
  wire  _T_1148; // @[CSR.scala 579:79:freechips.rocketchip.system.TinyConfig.fir@119369.4]
  wire  _T_1150; // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119371.4]
  wire  _T_1151; // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119372.4]
  wire  _T_1153; // @[CSR.scala 581:18:freechips.rocketchip.system.TinyConfig.fir@119378.4]
  wire  _T_1155; // @[CSR.scala 581:36:freechips.rocketchip.system.TinyConfig.fir@119380.4]
  wire  _T_1156; // @[CSR.scala 582:28:freechips.rocketchip.system.TinyConfig.fir@119384.4]
  wire  _T_1157; // @[CSR.scala 582:32:freechips.rocketchip.system.TinyConfig.fir@119385.4]
  wire  _T_1158; // @[CSR.scala 582:55:freechips.rocketchip.system.TinyConfig.fir@119386.4]
  wire  _T_1160; // @[CSR.scala 584:22:freechips.rocketchip.system.TinyConfig.fir@119391.4]
  wire  _T_1168; // @[CSR.scala 587:10:freechips.rocketchip.system.TinyConfig.fir@119409.4]
  wire  _T_1169; // @[CSR.scala 587:42:freechips.rocketchip.system.TinyConfig.fir@119410.4]
  wire  _T_1170; // @[CSR.scala 587:29:freechips.rocketchip.system.TinyConfig.fir@119411.4]
  wire  _T_1172; // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119413.4]
  wire  _T_1173; // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119414.4]
  wire [31:0] _T_1174; // @[CSR.scala 934:28:freechips.rocketchip.system.TinyConfig.fir@119419.4]
  wire [31:0] _T_1175; // @[CSR.scala 934:31:freechips.rocketchip.system.TinyConfig.fir@119420.4]
  wire [31:0] epc; // @[CSR.scala 934:26:freechips.rocketchip.system.TinyConfig.fir@119421.4]
  wire [1:0] _T_1177; // @[CSR.scala 598:86:freechips.rocketchip.system.TinyConfig.fir@119431.10]
  wire [1:0] _T_1178; // @[CSR.scala 598:56:freechips.rocketchip.system.TinyConfig.fir@119432.10]
  wire [1:0] _GEN_48; // @[CSR.scala 602:27:freechips.rocketchip.system.TinyConfig.fir@119440.8]
  wire [1:0] _GEN_67; // @[CSR.scala 594:24:freechips.rocketchip.system.TinyConfig.fir@119426.6]
  wire [1:0] _GEN_85; // @[CSR.scala 593:20:freechips.rocketchip.system.TinyConfig.fir@119425.4]
  wire  _T_1468; // @[CSR.scala 649:47:freechips.rocketchip.system.TinyConfig.fir@119758.8]
  wire [31:0] _GEN_95; // @[CSR.scala 649:53:freechips.rocketchip.system.TinyConfig.fir@119760.8]
  reg  _T_1481; // @[Reg.scala 27:20:freechips.rocketchip.system.TinyConfig.fir@119786.4]
  reg [31:0] _RAND_77;
  wire [31:0] _T_1483; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119804.4]
  wire [31:0] _T_1484; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119805.4]
  wire [31:0] _T_1485; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119806.4]
  wire [31:0] _T_1486; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119807.4]
  wire [31:0] _T_1487; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119808.4]
  wire [15:0] _T_1488; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119809.4]
  wire [31:0] _T_1489; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119810.4]
  wire [31:0] _T_1490; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119811.4]
  wire [31:0] _T_1491; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119812.4]
  wire [31:0] _T_1492; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119813.4]
  wire [31:0] _T_1493; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119814.4]
  wire [31:0] _T_1495; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119816.4]
  wire [31:0] _T_1496; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119817.4]
  wire [31:0] _T_1497; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119818.4]
  wire [63:0] _T_1498; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119819.4]
  wire [63:0] _T_1499; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119820.4]
  wire [31:0] _T_1587; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119908.4]
  wire [31:0] _T_1588; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119909.4]
  wire [31:0] _T_1589; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119910.4]
  wire [31:0] _T_1590; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119911.4]
  wire [29:0] _T_1593; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119914.4]
  wire [29:0] _T_1594; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119915.4]
  wire [29:0] _T_1595; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119916.4]
  wire [29:0] _T_1596; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119917.4]
  wire [29:0] _T_1597; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119918.4]
  wire [29:0] _T_1598; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119919.4]
  wire [29:0] _T_1599; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119920.4]
  wire [29:0] _T_1600; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119921.4]
  wire [31:0] _T_1610; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119931.4]
  wire [31:0] _T_1612; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119933.4]
  wire [31:0] _T_1614; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119935.4]
  wire [31:0] _T_1615; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119936.4]
  wire [31:0] _T_1616; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119937.4]
  wire [31:0] _T_1617; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119938.4]
  wire [31:0] _GEN_424; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119939.4]
  wire [31:0] _T_1618; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119939.4]
  wire [31:0] _T_1619; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119940.4]
  wire [31:0] _T_1620; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119941.4]
  wire [31:0] _T_1621; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119942.4]
  wire [31:0] _T_1622; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119943.4]
  wire [31:0] _T_1623; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119944.4]
  wire [31:0] _T_1625; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119946.4]
  wire [31:0] _T_1626; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119947.4]
  wire [31:0] _T_1627; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119948.4]
  wire [63:0] _GEN_425; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119949.4]
  wire [63:0] _T_1628; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119949.4]
  wire [63:0] _T_1629; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119950.4]
  wire [63:0] _GEN_426; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120038.4]
  wire [63:0] _T_1717; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120038.4]
  wire [63:0] _GEN_427; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120039.4]
  wire [63:0] _T_1718; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120039.4]
  wire [63:0] _GEN_428; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120040.4]
  wire [63:0] _T_1719; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120040.4]
  wire [63:0] _GEN_429; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120041.4]
  wire [63:0] _T_1720; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120041.4]
  wire [63:0] _GEN_430; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120044.4]
  wire [63:0] _T_1723; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120044.4]
  wire [63:0] _GEN_431; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120045.4]
  wire [63:0] _T_1724; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120045.4]
  wire [63:0] _GEN_432; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120046.4]
  wire [63:0] _T_1725; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120046.4]
  wire [63:0] _GEN_433; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120047.4]
  wire [63:0] _T_1726; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120047.4]
  wire [63:0] _GEN_434; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120048.4]
  wire [63:0] _T_1727; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120048.4]
  wire [63:0] _GEN_435; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120049.4]
  wire [63:0] _T_1728; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120049.4]
  wire [63:0] _GEN_436; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120050.4]
  wire [63:0] _T_1729; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120050.4]
  wire [63:0] _GEN_437; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120051.4]
  wire [63:0] _T_1730; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120051.4]
  wire [63:0] _GEN_438; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120061.4]
  wire [63:0] _T_1740; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120061.4]
  wire [63:0] _GEN_439; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120063.4]
  wire [63:0] _T_1742; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120063.4]
  wire  _T_1746; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120070.6]
  wire  _T_1747; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120071.6]
  wire  _T_1748; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120072.6]
  wire  _T_3320; // @[package.scala 15:62:freechips.rocketchip.system.TinyConfig.fir@122175.4]
  wire  csr_wen; // @[package.scala 15:62:freechips.rocketchip.system.TinyConfig.fir@122176.4]
  wire [101:0] _T_3334; // @[:freechips.rocketchip.system.TinyConfig.fir@122194.8 :freechips.rocketchip.system.TinyConfig.fir@122196.8]
  wire  _T_3338; // @[CSR.scala 701:47:freechips.rocketchip.system.TinyConfig.fir@122203.8]
  wire  _T_3342; // @[CSR.scala 701:47:freechips.rocketchip.system.TinyConfig.fir@122211.8]
  wire  _T_3365; // @[CSR.scala 725:20:freechips.rocketchip.system.TinyConfig.fir@122261.8]
  wire  _T_3366; // @[CSR.scala 727:39:freechips.rocketchip.system.TinyConfig.fir@122262.8]
  wire  _T_3367; // @[CSR.scala 727:33:freechips.rocketchip.system.TinyConfig.fir@122263.8]
  wire  _T_3369; // @[CSR.scala 727:51:freechips.rocketchip.system.TinyConfig.fir@122265.8]
  wire  _T_3370; // @[CSR.scala 727:43:freechips.rocketchip.system.TinyConfig.fir@122266.8]
  wire [31:0] _T_3371; // @[CSR.scala 729:25:freechips.rocketchip.system.TinyConfig.fir@122268.10]
  wire  _T_3372; // @[CSR.scala 729:35:freechips.rocketchip.system.TinyConfig.fir@122269.10]
  wire [3:0] _T_3373; // @[CSR.scala 729:38:freechips.rocketchip.system.TinyConfig.fir@122270.10]
  wire [31:0] _GEN_440; // @[CSR.scala 729:32:freechips.rocketchip.system.TinyConfig.fir@122271.10]
  wire [31:0] _T_3374; // @[CSR.scala 729:32:freechips.rocketchip.system.TinyConfig.fir@122271.10]
  wire [31:0] _T_3375; // @[CSR.scala 729:23:freechips.rocketchip.system.TinyConfig.fir@122272.10]
  wire [31:0] _T_3376; // @[CSR.scala 729:55:freechips.rocketchip.system.TinyConfig.fir@122273.10]
  wire [31:0] _T_3378; // @[CSR.scala 729:73:freechips.rocketchip.system.TinyConfig.fir@122275.10]
  wire [31:0] _T_3379; // @[CSR.scala 729:62:freechips.rocketchip.system.TinyConfig.fir@122276.10]
  wire [31:0] _T_3421; // @[CSR.scala 744:59:freechips.rocketchip.system.TinyConfig.fir@122343.8]
  wire [31:0] _T_3423; // @[CSR.scala 934:31:freechips.rocketchip.system.TinyConfig.fir@122348.8]
  wire [31:0] _T_3424; // @[CSR.scala 934:26:freechips.rocketchip.system.TinyConfig.fir@122349.8]
  wire [31:0] _T_3425; // @[CSR.scala 749:62:freechips.rocketchip.system.TinyConfig.fir@122359.8]
  wire [31:0] _T_3427; // @[CSR.scala 928:47:freechips.rocketchip.system.TinyConfig.fir@122367.8]
  wire [63:0] _T_3428; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122368.8]
  wire [57:0] _T_3429; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122370.8]
  wire [63:0] _GEN_130; // @[CSR.scala 928:31:freechips.rocketchip.system.TinyConfig.fir@122366.6]
  wire [31:0] _T_3431; // @[CSR.scala 929:74:freechips.rocketchip.system.TinyConfig.fir@122375.8]
  wire [63:0] _T_3432; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122376.8]
  wire [57:0] _T_3433; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122378.8]
  wire [63:0] _GEN_132; // @[CSR.scala 929:31:freechips.rocketchip.system.TinyConfig.fir@122373.6]
  wire [31:0] _T_3434; // @[CSR.scala 928:47:freechips.rocketchip.system.TinyConfig.fir@122382.8]
  wire [63:0] _T_3435; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122383.8]
  wire [57:0] _T_3436; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122385.8]
  wire [63:0] _GEN_134; // @[CSR.scala 928:31:freechips.rocketchip.system.TinyConfig.fir@122381.6]
  wire [31:0] _T_3438; // @[CSR.scala 929:74:freechips.rocketchip.system.TinyConfig.fir@122390.8]
  wire [63:0] _T_3439; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122391.8]
  wire [57:0] _T_3440; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122393.8]
  wire [63:0] _GEN_136; // @[CSR.scala 929:31:freechips.rocketchip.system.TinyConfig.fir@122388.6]
  wire  _T_3453; // @[CSR.scala 768:43:freechips.rocketchip.system.TinyConfig.fir@122422.8]
  wire  _T_3461; // @[CSR.scala 819:37:freechips.rocketchip.system.TinyConfig.fir@122446.6]
  wire  _T_3462; // @[CSR.scala 819:55:freechips.rocketchip.system.TinyConfig.fir@122447.6]
  wire  _T_3466; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122459.10]
  wire  _T_3467; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122461.10]
  wire [1:0] _T_3473; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122473.10]
  wire [31:0] _T_3496; // @[CSR.scala 913:9:freechips.rocketchip.system.TinyConfig.fir@122505.10]
  wire [31:0] _T_3497; // @[CSR.scala 913:34:freechips.rocketchip.system.TinyConfig.fir@122506.10]
  wire [31:0] _T_3502; // @[CSR.scala 913:43:freechips.rocketchip.system.TinyConfig.fir@122511.10]
  wire  _T_3515; // @[CSR.scala 828:96:freechips.rocketchip.system.TinyConfig.fir@122537.10]
  wire  _T_3518; // @[CSR.scala 828:96:freechips.rocketchip.system.TinyConfig.fir@122543.10]
  wire  _T_3520; // @[CSR.scala 829:38:freechips.rocketchip.system.TinyConfig.fir@122547.10]
  wire  _T_3604; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122693.6]
  wire  _T_3605; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122694.6]
  wire [7:0] _T_3608; // @[:freechips.rocketchip.system.TinyConfig.fir@122699.8 :freechips.rocketchip.system.TinyConfig.fir@122701.8]
  wire  _T_3609; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122702.8]
  wire  _T_3610; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122704.8]
  wire  _T_3611; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122706.8]
  wire [1:0] _T_3612; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122708.8]
  wire  _T_3614; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122712.8]
  wire  _T_3615; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122715.8]
  wire  _T_3616; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122718.6]
  wire  _T_3617; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122719.6]
  wire  _T_3619; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122721.6]
  wire  _T_3620; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122722.6]
  wire  _T_3621; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122723.6]
  wire  _T_3622; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122724.6]
  wire  _T_3623; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122725.6]
  wire [31:0] _GEN_215; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122726.6]
  wire  _T_3624; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122729.6]
  wire  _T_3625; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122730.6]
  wire [23:0] _T_3626; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122732.8]
  wire [7:0] _T_3628; // @[:freechips.rocketchip.system.TinyConfig.fir@122735.8 :freechips.rocketchip.system.TinyConfig.fir@122737.8]
  wire  _T_3629; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122738.8]
  wire  _T_3630; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122740.8]
  wire  _T_3631; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122742.8]
  wire [1:0] _T_3632; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122744.8]
  wire  _T_3634; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122748.8]
  wire  _T_3635; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122751.8]
  wire  _T_3636; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122754.6]
  wire  _T_3637; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122755.6]
  wire  _T_3639; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122757.6]
  wire  _T_3640; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122758.6]
  wire  _T_3641; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122759.6]
  wire  _T_3642; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122760.6]
  wire  _T_3643; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122761.6]
  wire [31:0] _GEN_222; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122762.6]
  wire  _T_3644; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122765.6]
  wire  _T_3645; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122766.6]
  wire [15:0] _T_3646; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122768.8]
  wire [7:0] _T_3648; // @[:freechips.rocketchip.system.TinyConfig.fir@122771.8 :freechips.rocketchip.system.TinyConfig.fir@122773.8]
  wire  _T_3649; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122774.8]
  wire  _T_3650; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122776.8]
  wire  _T_3651; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122778.8]
  wire [1:0] _T_3652; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122780.8]
  wire  _T_3654; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122784.8]
  wire  _T_3655; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122787.8]
  wire  _T_3656; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122790.6]
  wire  _T_3657; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122791.6]
  wire  _T_3659; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122793.6]
  wire  _T_3660; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122794.6]
  wire  _T_3661; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122795.6]
  wire  _T_3662; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122796.6]
  wire  _T_3663; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122797.6]
  wire [31:0] _GEN_229; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122798.6]
  wire  _T_3664; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122801.6]
  wire  _T_3665; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122802.6]
  wire [7:0] _T_3666; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122804.8]
  wire  _T_3669; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122810.8]
  wire  _T_3670; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122812.8]
  wire  _T_3671; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122814.8]
  wire [1:0] _T_3672; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122816.8]
  wire  _T_3674; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122820.8]
  wire  _T_3675; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122823.8]
  wire  _T_3676; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122826.6]
  wire  _T_3677; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122827.6]
  wire  _T_3679; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122829.6]
  wire  _T_3680; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122830.6]
  wire  _T_3681; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122831.6]
  wire  _T_3682; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122832.6]
  wire  _T_3683; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122833.6]
  wire [31:0] _GEN_236; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122834.6]
  wire  _T_3684; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122837.6]
  wire  _T_3685; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122838.6]
  wire  _T_3696; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122862.6]
  wire  _T_3697; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122863.6]
  wire  _T_3699; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122865.6]
  wire  _T_3700; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122866.6]
  wire  _T_3701; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122867.6]
  wire  _T_3702; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122868.6]
  wire  _T_3703; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122869.6]
  wire [31:0] _GEN_243; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122870.6]
  wire  _T_3704; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122873.6]
  wire  _T_3705; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122874.6]
  wire  _T_3716; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122898.6]
  wire  _T_3717; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122899.6]
  wire  _T_3719; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122901.6]
  wire  _T_3720; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122902.6]
  wire  _T_3721; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122903.6]
  wire  _T_3722; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122904.6]
  wire  _T_3723; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122905.6]
  wire [31:0] _GEN_250; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122906.6]
  wire  _T_3724; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122909.6]
  wire  _T_3725; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122910.6]
  wire  _T_3736; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122934.6]
  wire  _T_3737; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122935.6]
  wire  _T_3739; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122937.6]
  wire  _T_3740; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122938.6]
  wire  _T_3741; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122939.6]
  wire  _T_3742; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122940.6]
  wire  _T_3743; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122941.6]
  wire [31:0] _GEN_257; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122942.6]
  wire  _T_3744; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122945.6]
  wire  _T_3745; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122946.6]
  wire  _T_3761; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122975.6]
  wire  _T_3762; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122976.6]
  wire  _T_3763; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122977.6]
  wire [31:0] _GEN_264; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122978.6]
  wire [63:0] _GEN_282; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [63:0] _GEN_284; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_329; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_336; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_343; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_350; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_357; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_364; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_371; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire [31:0] _GEN_378; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  wire  _T_3810; // @[CSR.scala 892:26:freechips.rocketchip.system.TinyConfig.fir@123141.4]
  assign _GEN_415 = {{5'd0}, io_retire}; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118189.4]
  assign _T_84 = _T_83 + _GEN_415; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118189.4]
  assign _T_86 = _T_84[6]; // @[Counters.scala 52:20:freechips.rocketchip.system.TinyConfig.fir@118192.4]
  assign _T_88 = _T_85 + 58'h1; // @[Counters.scala 52:43:freechips.rocketchip.system.TinyConfig.fir@118195.6]
  assign _T_89 = {_T_85,_T_83}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118198.4]
  assign _T_90 = io_csr_stall == 1'h0; // @[CSR.scala 338:103:freechips.rocketchip.system.TinyConfig.fir@118199.4]
  assign _GEN_416 = {{5'd0}, _T_90}; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118201.4]
  assign _T_92 = _T_91 + _GEN_416; // @[Counters.scala 47:33:freechips.rocketchip.system.TinyConfig.fir@118201.4]
  assign _T_94 = _T_92[6]; // @[Counters.scala 52:20:freechips.rocketchip.system.TinyConfig.fir@118204.4]
  assign _T_96 = _T_93 + 58'h1; // @[Counters.scala 52:43:freechips.rocketchip.system.TinyConfig.fir@118207.6]
  assign _T_97 = {_T_93,_T_91}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118210.4]
  assign _T_112 = {4'h0,io_interrupts_meip,1'h0,2'h0,io_interrupts_mtip,1'h0,2'h0,io_interrupts_msip,1'h0,2'h0}; // @[CSR.scala 351:22:freechips.rocketchip.system.TinyConfig.fir@118232.4]
  assign read_mip = _T_112 & 16'h888; // @[CSR.scala 351:29:freechips.rocketchip.system.TinyConfig.fir@118233.4]
  assign _GEN_417 = {{16'd0}, read_mip}; // @[CSR.scala 354:56:freechips.rocketchip.system.TinyConfig.fir@118234.4]
  assign pending_interrupts = _GEN_417 & reg_mie; // @[CSR.scala 354:56:freechips.rocketchip.system.TinyConfig.fir@118234.4]
  assign d_interrupts = {io_interrupts_debug, 14'h0}; // @[CSR.scala 355:42:freechips.rocketchip.system.TinyConfig.fir@118236.4]
  assign _T_116 = ~ pending_interrupts; // @[CSR.scala 356:73:freechips.rocketchip.system.TinyConfig.fir@118239.4]
  assign _T_118 = ~ _T_116; // @[CSR.scala 356:71:freechips.rocketchip.system.TinyConfig.fir@118241.4]
  assign m_interrupts = reg_mstatus_mie ? _T_118 : 32'h0; // @[CSR.scala 356:25:freechips.rocketchip.system.TinyConfig.fir@118242.4]
  assign _T_124 = d_interrupts[14]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118249.4]
  assign _T_125 = d_interrupts[13]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118250.4]
  assign _T_126 = d_interrupts[12]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118251.4]
  assign _T_127 = d_interrupts[11]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118252.4]
  assign _T_128 = d_interrupts[3]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118253.4]
  assign _T_129 = d_interrupts[7]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118254.4]
  assign _T_130 = d_interrupts[9]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118255.4]
  assign _T_131 = d_interrupts[1]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118256.4]
  assign _T_132 = d_interrupts[5]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118257.4]
  assign _T_133 = d_interrupts[8]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118258.4]
  assign _T_134 = d_interrupts[0]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118259.4]
  assign _T_135 = d_interrupts[4]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118260.4]
  assign _T_136 = m_interrupts[15]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118261.4]
  assign _T_137 = m_interrupts[14]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118262.4]
  assign _T_138 = m_interrupts[13]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118263.4]
  assign _T_139 = m_interrupts[12]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118264.4]
  assign _T_140 = m_interrupts[11]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118265.4]
  assign _T_141 = m_interrupts[3]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118266.4]
  assign _T_142 = m_interrupts[7]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118267.4]
  assign _T_143 = m_interrupts[9]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118268.4]
  assign _T_144 = m_interrupts[1]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118269.4]
  assign _T_145 = m_interrupts[5]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118270.4]
  assign _T_146 = m_interrupts[8]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118271.4]
  assign _T_147 = m_interrupts[0]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118272.4]
  assign _T_148 = m_interrupts[4]; // @[CSR.scala 907:76:freechips.rocketchip.system.TinyConfig.fir@118273.4]
  assign _T_162 = _T_124 | _T_125; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118287.4]
  assign _T_163 = _T_162 | _T_126; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118288.4]
  assign _T_164 = _T_163 | _T_127; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118289.4]
  assign _T_165 = _T_164 | _T_128; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118290.4]
  assign _T_166 = _T_165 | _T_129; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118291.4]
  assign _T_167 = _T_166 | _T_130; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118292.4]
  assign _T_168 = _T_167 | _T_131; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118293.4]
  assign _T_169 = _T_168 | _T_132; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118294.4]
  assign _T_170 = _T_169 | _T_133; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118295.4]
  assign _T_171 = _T_170 | _T_134; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118296.4]
  assign _T_172 = _T_171 | _T_135; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118297.4]
  assign _T_173 = _T_172 | _T_136; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118298.4]
  assign _T_174 = _T_173 | _T_137; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118299.4]
  assign _T_175 = _T_174 | _T_138; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118300.4]
  assign _T_176 = _T_175 | _T_139; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118301.4]
  assign _T_177 = _T_176 | _T_140; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118302.4]
  assign _T_178 = _T_177 | _T_141; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118303.4]
  assign _T_179 = _T_178 | _T_142; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118304.4]
  assign _T_180 = _T_179 | _T_143; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118305.4]
  assign _T_181 = _T_180 | _T_144; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118306.4]
  assign _T_182 = _T_181 | _T_145; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118307.4]
  assign _T_183 = _T_182 | _T_146; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118308.4]
  assign _T_184 = _T_183 | _T_147; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118309.4]
  assign anyInterrupt = _T_184 | _T_148; // @[CSR.scala 907:90:freechips.rocketchip.system.TinyConfig.fir@118310.4]
  assign _T_249 = _T_147 ? 4'h0 : 4'h4; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118375.4]
  assign _T_250 = _T_146 ? 4'h8 : _T_249; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118376.4]
  assign _T_251 = _T_145 ? 4'h5 : _T_250; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118377.4]
  assign _T_252 = _T_144 ? 4'h1 : _T_251; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118378.4]
  assign _T_253 = _T_143 ? 4'h9 : _T_252; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118379.4]
  assign _T_254 = _T_142 ? 4'h7 : _T_253; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118380.4]
  assign _T_255 = _T_141 ? 4'h3 : _T_254; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118381.4]
  assign _T_256 = _T_140 ? 4'hb : _T_255; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118382.4]
  assign _T_257 = _T_139 ? 4'hc : _T_256; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118383.4]
  assign _T_258 = _T_138 ? 4'hd : _T_257; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118384.4]
  assign _T_259 = _T_137 ? 4'he : _T_258; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118385.4]
  assign _T_260 = _T_136 ? 4'hf : _T_259; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118386.4]
  assign _T_261 = _T_135 ? 4'h4 : _T_260; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118387.4]
  assign _T_262 = _T_134 ? 4'h0 : _T_261; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118388.4]
  assign _T_263 = _T_133 ? 4'h8 : _T_262; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118389.4]
  assign _T_264 = _T_132 ? 4'h5 : _T_263; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118390.4]
  assign _T_265 = _T_131 ? 4'h1 : _T_264; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118391.4]
  assign _T_266 = _T_130 ? 4'h9 : _T_265; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118392.4]
  assign _T_267 = _T_129 ? 4'h7 : _T_266; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118393.4]
  assign _T_268 = _T_128 ? 4'h3 : _T_267; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118394.4]
  assign _T_269 = _T_127 ? 4'hb : _T_268; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118395.4]
  assign _T_270 = _T_126 ? 4'hc : _T_269; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118396.4]
  assign _T_271 = _T_125 ? 4'hd : _T_270; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118397.4]
  assign whichInterrupt = _T_124 ? 4'he : _T_271; // @[Mux.scala 48:69:freechips.rocketchip.system.TinyConfig.fir@118398.4]
  assign _GEN_418 = {{28'd0}, whichInterrupt}; // @[CSR.scala 360:43:freechips.rocketchip.system.TinyConfig.fir@118399.4]
  assign _T_273 = io_singleStep == 1'h0; // @[CSR.scala 361:36:freechips.rocketchip.system.TinyConfig.fir@118401.4]
  assign _T_274 = anyInterrupt & _T_273; // @[CSR.scala 361:33:freechips.rocketchip.system.TinyConfig.fir@118402.4]
  assign _T_275 = _T_274 | reg_singleStepped; // @[CSR.scala 361:51:freechips.rocketchip.system.TinyConfig.fir@118403.4]
  assign _T_276 = reg_debug | io_status_cease; // @[CSR.scala 361:88:freechips.rocketchip.system.TinyConfig.fir@118404.4]
  assign _T_277 = _T_276 == 1'h0; // @[CSR.scala 361:76:freechips.rocketchip.system.TinyConfig.fir@118405.4]
  assign _T_280 = reg_pmp_0_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118413.4]
  assign _T_281 = {reg_pmp_0_addr,_T_280}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118414.4]
  assign _T_284 = _T_281 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118417.4]
  assign _T_285 = ~ _T_284; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118418.4]
  assign _T_286 = _T_281 & _T_285; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118419.4]
  assign _T_287 = {_T_286,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118420.4]
  assign _T_289 = reg_pmp_1_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118425.4]
  assign _T_290 = {reg_pmp_1_addr,_T_289}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118426.4]
  assign _T_293 = _T_290 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118429.4]
  assign _T_294 = ~ _T_293; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118430.4]
  assign _T_295 = _T_290 & _T_294; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118431.4]
  assign _T_296 = {_T_295,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118432.4]
  assign _T_298 = reg_pmp_2_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118437.4]
  assign _T_299 = {reg_pmp_2_addr,_T_298}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118438.4]
  assign _T_302 = _T_299 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118441.4]
  assign _T_303 = ~ _T_302; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118442.4]
  assign _T_304 = _T_299 & _T_303; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118443.4]
  assign _T_305 = {_T_304,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118444.4]
  assign _T_307 = reg_pmp_3_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118449.4]
  assign _T_308 = {reg_pmp_3_addr,_T_307}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118450.4]
  assign _T_311 = _T_308 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118453.4]
  assign _T_312 = ~ _T_311; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118454.4]
  assign _T_313 = _T_308 & _T_312; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118455.4]
  assign _T_314 = {_T_313,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118456.4]
  assign _T_316 = reg_pmp_4_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118461.4]
  assign _T_317 = {reg_pmp_4_addr,_T_316}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118462.4]
  assign _T_320 = _T_317 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118465.4]
  assign _T_321 = ~ _T_320; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118466.4]
  assign _T_322 = _T_317 & _T_321; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118467.4]
  assign _T_323 = {_T_322,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118468.4]
  assign _T_325 = reg_pmp_5_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118473.4]
  assign _T_326 = {reg_pmp_5_addr,_T_325}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118474.4]
  assign _T_329 = _T_326 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118477.4]
  assign _T_330 = ~ _T_329; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118478.4]
  assign _T_331 = _T_326 & _T_330; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118479.4]
  assign _T_332 = {_T_331,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118480.4]
  assign _T_334 = reg_pmp_6_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118485.4]
  assign _T_335 = {reg_pmp_6_addr,_T_334}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118486.4]
  assign _T_338 = _T_335 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118489.4]
  assign _T_339 = ~ _T_338; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118490.4]
  assign _T_340 = _T_335 & _T_339; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118491.4]
  assign _T_341 = {_T_340,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118492.4]
  assign _T_343 = reg_pmp_7_cfg_a[0]; // @[PMP.scala 57:31:freechips.rocketchip.system.TinyConfig.fir@118497.4]
  assign _T_344 = {reg_pmp_7_addr,_T_343}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118498.4]
  assign _T_347 = _T_344 + 31'h1; // @[PMP.scala 58:23:freechips.rocketchip.system.TinyConfig.fir@118501.4]
  assign _T_348 = ~ _T_347; // @[PMP.scala 58:16:freechips.rocketchip.system.TinyConfig.fir@118502.4]
  assign _T_349 = _T_344 & _T_348; // @[PMP.scala 58:14:freechips.rocketchip.system.TinyConfig.fir@118503.4]
  assign _T_350 = {_T_349,2'h3}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118504.4]
  assign _T_356 = {io_status_hpie,io_status_spie,io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie}; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118520.4]
  assign _T_364 = {io_status_sum,io_status_mprv,io_status_xs,io_status_fs,io_status_mpp,io_status_hpp,io_status_spp,io_status_mpie,_T_356}; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118528.4]
  assign _T_370 = {io_status_uxl,io_status_sd_rv32,io_status_zero1,io_status_tsr,io_status_tw,io_status_tvm,io_status_mxr}; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118534.4]
  assign _T_379 = {io_status_debug,io_status_cease,io_status_isa,io_status_dprv,io_status_prv,io_status_sd,io_status_zero2,io_status_sxl,_T_370,_T_364}; // @[CSR.scala 379:38:freechips.rocketchip.system.TinyConfig.fir@118543.4]
  assign read_mstatus = _T_379[31:0]; // @[CSR.scala 379:40:freechips.rocketchip.system.TinyConfig.fir@118544.4]
  assign _T_380 = reg_mtvec[0]; // @[CSR.scala 936:41:freechips.rocketchip.system.TinyConfig.fir@118545.4]
  assign _T_381 = _T_380 ? 7'h7e : 7'h2; // @[CSR.scala 936:39:freechips.rocketchip.system.TinyConfig.fir@118546.4]
  assign _T_383 = {{25'd0}, _T_381}; // @[package.scala 131:41:freechips.rocketchip.system.TinyConfig.fir@118548.4]
  assign _T_384 = ~ _T_383; // @[package.scala 131:37:freechips.rocketchip.system.TinyConfig.fir@118549.4]
  assign read_mtvec = reg_mtvec & _T_384; // @[package.scala 131:35:freechips.rocketchip.system.TinyConfig.fir@118550.4]
  assign _T_395 = {4'h8,reg_bp_0_control_x,reg_bp_0_control_w,reg_bp_0_control_r}; // @[CSR.scala 385:48:freechips.rocketchip.system.TinyConfig.fir@118562.4]
  assign _T_403 = {4'h2,reg_bp_0_control_dmode,14'h400,reg_bp_0_control_action,1'h0,2'h0,reg_bp_0_control_tmatch,_T_395}; // @[CSR.scala 385:48:freechips.rocketchip.system.TinyConfig.fir@118570.4]
  assign _T_404 = ~ reg_mepc; // @[CSR.scala 935:28:freechips.rocketchip.system.TinyConfig.fir@118571.4]
  assign _T_405 = reg_misa[2]; // @[CSR.scala 935:45:freechips.rocketchip.system.TinyConfig.fir@118572.4]
  assign _T_406 = _T_405 ? 2'h1 : 2'h3; // @[CSR.scala 935:36:freechips.rocketchip.system.TinyConfig.fir@118573.4]
  assign _GEN_419 = {{30'd0}, _T_406}; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118574.4]
  assign _T_407 = _T_404 | _GEN_419; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118574.4]
  assign _T_408 = ~ _T_407; // @[CSR.scala 935:26:freechips.rocketchip.system.TinyConfig.fir@118575.4]
  assign _T_421 = {4'h4,12'h0,reg_dcsr_ebreakm,3'h0,2'h0,1'h0,reg_dcsr_cause,3'h0,reg_dcsr_step,2'h3}; // @[CSR.scala 399:27:freechips.rocketchip.system.TinyConfig.fir@118588.4]
  assign _T_422 = ~ reg_dpc; // @[CSR.scala 935:28:freechips.rocketchip.system.TinyConfig.fir@118589.4]
  assign _T_425 = _T_422 | _GEN_419; // @[CSR.scala 935:31:freechips.rocketchip.system.TinyConfig.fir@118592.4]
  assign _T_426 = ~ _T_425; // @[CSR.scala 935:26:freechips.rocketchip.system.TinyConfig.fir@118593.4]
  assign _T_457 = _T_97[63:32]; // @[CSR.scala 436:50:freechips.rocketchip.system.TinyConfig.fir@118624.4]
  assign _T_458 = _T_89[63:32]; // @[CSR.scala 437:54:freechips.rocketchip.system.TinyConfig.fir@118625.4]
  assign _T_473 = {reg_pmp_0_cfg_l,2'h0,reg_pmp_0_cfg_a,reg_pmp_0_cfg_x,reg_pmp_0_cfg_w,reg_pmp_0_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118651.4]
  assign _T_483 = {reg_pmp_2_cfg_l,2'h0,reg_pmp_2_cfg_a,reg_pmp_2_cfg_x,reg_pmp_2_cfg_w,reg_pmp_2_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118661.4]
  assign _T_489 = {reg_pmp_1_cfg_l,2'h0,reg_pmp_1_cfg_a,reg_pmp_1_cfg_x,reg_pmp_1_cfg_w,reg_pmp_1_cfg_r,_T_473}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118667.4]
  assign _T_491 = {reg_pmp_3_cfg_l,2'h0,reg_pmp_3_cfg_a,reg_pmp_3_cfg_x,reg_pmp_3_cfg_w,reg_pmp_3_cfg_r,_T_483,_T_489}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118669.4]
  assign _T_496 = {reg_pmp_4_cfg_l,2'h0,reg_pmp_4_cfg_a,reg_pmp_4_cfg_x,reg_pmp_4_cfg_w,reg_pmp_4_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118674.4]
  assign _T_506 = {reg_pmp_6_cfg_l,2'h0,reg_pmp_6_cfg_a,reg_pmp_6_cfg_x,reg_pmp_6_cfg_w,reg_pmp_6_cfg_r}; // @[package.scala 36:38:freechips.rocketchip.system.TinyConfig.fir@118684.4]
  assign _T_512 = {reg_pmp_5_cfg_l,2'h0,reg_pmp_5_cfg_a,reg_pmp_5_cfg_x,reg_pmp_5_cfg_w,reg_pmp_5_cfg_r,_T_496}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118690.4]
  assign _T_514 = {reg_pmp_7_cfg_l,2'h0,reg_pmp_7_cfg_a,reg_pmp_7_cfg_x,reg_pmp_7_cfg_w,reg_pmp_7_cfg_r,_T_506,_T_512}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@118692.4]
  assign _T_562 = io_rw_addr == 12'h7a1; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118744.4]
  assign _T_563 = io_rw_addr == 12'h7a2; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118745.4]
  assign _T_564 = io_rw_addr == 12'h301; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118746.4]
  assign _T_565 = io_rw_addr == 12'h300; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118747.4]
  assign _T_566 = io_rw_addr == 12'h305; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118748.4]
  assign _T_567 = io_rw_addr == 12'h344; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118749.4]
  assign _T_568 = io_rw_addr == 12'h304; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118750.4]
  assign _T_569 = io_rw_addr == 12'h340; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118751.4]
  assign _T_570 = io_rw_addr == 12'h341; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118752.4]
  assign _T_571 = io_rw_addr == 12'h343; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118753.4]
  assign _T_572 = io_rw_addr == 12'h342; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118754.4]
  assign _T_574 = io_rw_addr == 12'h7b0; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118756.4]
  assign _T_575 = io_rw_addr == 12'h7b1; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118757.4]
  assign _T_576 = io_rw_addr == 12'h7b2; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118758.4]
  assign _T_577 = io_rw_addr == 12'hb00; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118759.4]
  assign _T_578 = io_rw_addr == 12'hb02; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118760.4]
  assign _T_666 = io_rw_addr == 12'hb80; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118848.4]
  assign _T_667 = io_rw_addr == 12'hb82; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118849.4]
  assign _T_668 = io_rw_addr == 12'h3a0; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118850.4]
  assign _T_669 = io_rw_addr == 12'h3a1; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118851.4]
  assign _T_672 = io_rw_addr == 12'h3b0; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118854.4]
  assign _T_673 = io_rw_addr == 12'h3b1; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118855.4]
  assign _T_674 = io_rw_addr == 12'h3b2; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118856.4]
  assign _T_675 = io_rw_addr == 12'h3b3; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118857.4]
  assign _T_676 = io_rw_addr == 12'h3b4; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118858.4]
  assign _T_677 = io_rw_addr == 12'h3b5; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118859.4]
  assign _T_678 = io_rw_addr == 12'h3b6; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118860.4]
  assign _T_679 = io_rw_addr == 12'h3b7; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118861.4]
  assign _T_689 = io_rw_addr == 12'hf12; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118871.4]
  assign _T_691 = io_rw_addr == 12'hf13; // @[CSR.scala 497:73:freechips.rocketchip.system.TinyConfig.fir@118873.4]
  assign _T_692 = io_rw_cmd[1]; // @[CSR.scala 913:13:freechips.rocketchip.system.TinyConfig.fir@118874.4]
  assign _T_693 = _T_692 ? io_rw_rdata : 32'h0; // @[CSR.scala 913:9:freechips.rocketchip.system.TinyConfig.fir@118875.4]
  assign _T_694 = _T_693 | io_rw_wdata; // @[CSR.scala 913:34:freechips.rocketchip.system.TinyConfig.fir@118876.4]
  assign _T_695 = io_rw_cmd[1:0]; // @[CSR.scala 913:53:freechips.rocketchip.system.TinyConfig.fir@118877.4]
  assign _T_696 = _T_695 == 2'h3; // @[CSR.scala 913:59:freechips.rocketchip.system.TinyConfig.fir@118878.4]
  assign _T_697 = _T_696 ? io_rw_wdata : 32'h0; // @[CSR.scala 913:49:freechips.rocketchip.system.TinyConfig.fir@118879.4]
  assign _T_698 = ~ _T_697; // @[CSR.scala 913:45:freechips.rocketchip.system.TinyConfig.fir@118880.4]
  assign wdata = _T_694 & _T_698; // @[CSR.scala 913:43:freechips.rocketchip.system.TinyConfig.fir@118881.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 500:31:freechips.rocketchip.system.TinyConfig.fir@118882.4]
  assign _T_699 = {io_rw_addr, 20'h0}; // @[CSR.scala 512:28:freechips.rocketchip.system.TinyConfig.fir@118883.4]
  assign _T_700 = _T_699 & 32'h20100000; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118884.4]
  assign _T_701 = _T_700 == 32'h0; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118885.4]
  assign _T_703 = _T_699 & 32'h10100000; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118887.4]
  assign _T_704 = _T_703 == 32'h100000; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118888.4]
  assign _T_706 = _T_699 & 32'h20400000; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118890.4]
  assign _T_707 = _T_706 == 32'h20000000; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118891.4]
  assign _T_709 = _T_699 & 32'h20200000; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118893.4]
  assign _T_710 = _T_709 == 32'h20000000; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118894.4]
  assign _T_712 = _T_699 & 32'h30000000; // @[Decode.scala 14:65:freechips.rocketchip.system.TinyConfig.fir@118896.4]
  assign _T_713 = _T_712 == 32'h10000000; // @[Decode.scala 14:121:freechips.rocketchip.system.TinyConfig.fir@118897.4]
  assign insn_call = system_insn & _T_701; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118900.4]
  assign insn_break = system_insn & _T_704; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118902.4]
  assign insn_ret = system_insn & _T_707; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118904.4]
  assign insn_cease = system_insn & _T_710; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118906.4]
  assign insn_wfi = system_insn & _T_713; // @[CSR.scala 512:95:freechips.rocketchip.system.TinyConfig.fir@118908.4]
  assign _T_764 = io_status_fs == 2'h0; // @[CSR.scala 524:39:freechips.rocketchip.system.TinyConfig.fir@118954.4]
  assign _T_765 = reg_misa[5]; // @[CSR.scala 524:57:freechips.rocketchip.system.TinyConfig.fir@118955.4]
  assign _T_766 = _T_765 == 1'h0; // @[CSR.scala 524:48:freechips.rocketchip.system.TinyConfig.fir@118956.4]
  assign _T_779 = io_decode_0_csr == 12'h7a0; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118972.4]
  assign _T_780 = io_decode_0_csr == 12'h7a1; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118973.4]
  assign _T_781 = io_decode_0_csr == 12'h7a2; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118974.4]
  assign _T_782 = io_decode_0_csr == 12'h301; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118975.4]
  assign _T_783 = io_decode_0_csr == 12'h300; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118976.4]
  assign _T_784 = io_decode_0_csr == 12'h305; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118977.4]
  assign _T_785 = io_decode_0_csr == 12'h344; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118978.4]
  assign _T_786 = io_decode_0_csr == 12'h304; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118979.4]
  assign _T_787 = io_decode_0_csr == 12'h340; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118980.4]
  assign _T_788 = io_decode_0_csr == 12'h341; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118981.4]
  assign _T_789 = io_decode_0_csr == 12'h343; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118982.4]
  assign _T_790 = io_decode_0_csr == 12'h342; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118983.4]
  assign _T_791 = io_decode_0_csr == 12'hf14; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118984.4]
  assign _T_792 = io_decode_0_csr == 12'h7b0; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118985.4]
  assign _T_793 = io_decode_0_csr == 12'h7b1; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118986.4]
  assign _T_794 = io_decode_0_csr == 12'h7b2; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118987.4]
  assign _T_795 = io_decode_0_csr == 12'hb00; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118988.4]
  assign _T_796 = io_decode_0_csr == 12'hb02; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118989.4]
  assign _T_797 = io_decode_0_csr == 12'h323; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118990.4]
  assign _T_798 = io_decode_0_csr == 12'hb03; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118991.4]
  assign _T_799 = io_decode_0_csr == 12'hb83; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118992.4]
  assign _T_800 = io_decode_0_csr == 12'h324; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118993.4]
  assign _T_801 = io_decode_0_csr == 12'hb04; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118994.4]
  assign _T_802 = io_decode_0_csr == 12'hb84; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118995.4]
  assign _T_803 = io_decode_0_csr == 12'h325; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118996.4]
  assign _T_804 = io_decode_0_csr == 12'hb05; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118997.4]
  assign _T_805 = io_decode_0_csr == 12'hb85; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118998.4]
  assign _T_806 = io_decode_0_csr == 12'h326; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@118999.4]
  assign _T_807 = io_decode_0_csr == 12'hb06; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119000.4]
  assign _T_808 = io_decode_0_csr == 12'hb86; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119001.4]
  assign _T_809 = io_decode_0_csr == 12'h327; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119002.4]
  assign _T_810 = io_decode_0_csr == 12'hb07; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119003.4]
  assign _T_811 = io_decode_0_csr == 12'hb87; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119004.4]
  assign _T_812 = io_decode_0_csr == 12'h328; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119005.4]
  assign _T_813 = io_decode_0_csr == 12'hb08; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119006.4]
  assign _T_814 = io_decode_0_csr == 12'hb88; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119007.4]
  assign _T_815 = io_decode_0_csr == 12'h329; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119008.4]
  assign _T_816 = io_decode_0_csr == 12'hb09; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119009.4]
  assign _T_817 = io_decode_0_csr == 12'hb89; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119010.4]
  assign _T_818 = io_decode_0_csr == 12'h32a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119011.4]
  assign _T_819 = io_decode_0_csr == 12'hb0a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119012.4]
  assign _T_820 = io_decode_0_csr == 12'hb8a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119013.4]
  assign _T_821 = io_decode_0_csr == 12'h32b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119014.4]
  assign _T_822 = io_decode_0_csr == 12'hb0b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119015.4]
  assign _T_823 = io_decode_0_csr == 12'hb8b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119016.4]
  assign _T_824 = io_decode_0_csr == 12'h32c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119017.4]
  assign _T_825 = io_decode_0_csr == 12'hb0c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119018.4]
  assign _T_826 = io_decode_0_csr == 12'hb8c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119019.4]
  assign _T_827 = io_decode_0_csr == 12'h32d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119020.4]
  assign _T_828 = io_decode_0_csr == 12'hb0d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119021.4]
  assign _T_829 = io_decode_0_csr == 12'hb8d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119022.4]
  assign _T_830 = io_decode_0_csr == 12'h32e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119023.4]
  assign _T_831 = io_decode_0_csr == 12'hb0e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119024.4]
  assign _T_832 = io_decode_0_csr == 12'hb8e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119025.4]
  assign _T_833 = io_decode_0_csr == 12'h32f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119026.4]
  assign _T_834 = io_decode_0_csr == 12'hb0f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119027.4]
  assign _T_835 = io_decode_0_csr == 12'hb8f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119028.4]
  assign _T_836 = io_decode_0_csr == 12'h330; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119029.4]
  assign _T_837 = io_decode_0_csr == 12'hb10; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119030.4]
  assign _T_838 = io_decode_0_csr == 12'hb90; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119031.4]
  assign _T_839 = io_decode_0_csr == 12'h331; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119032.4]
  assign _T_840 = io_decode_0_csr == 12'hb11; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119033.4]
  assign _T_841 = io_decode_0_csr == 12'hb91; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119034.4]
  assign _T_842 = io_decode_0_csr == 12'h332; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119035.4]
  assign _T_843 = io_decode_0_csr == 12'hb12; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119036.4]
  assign _T_844 = io_decode_0_csr == 12'hb92; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119037.4]
  assign _T_845 = io_decode_0_csr == 12'h333; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119038.4]
  assign _T_846 = io_decode_0_csr == 12'hb13; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119039.4]
  assign _T_847 = io_decode_0_csr == 12'hb93; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119040.4]
  assign _T_848 = io_decode_0_csr == 12'h334; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119041.4]
  assign _T_849 = io_decode_0_csr == 12'hb14; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119042.4]
  assign _T_850 = io_decode_0_csr == 12'hb94; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119043.4]
  assign _T_851 = io_decode_0_csr == 12'h335; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119044.4]
  assign _T_852 = io_decode_0_csr == 12'hb15; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119045.4]
  assign _T_853 = io_decode_0_csr == 12'hb95; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119046.4]
  assign _T_854 = io_decode_0_csr == 12'h336; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119047.4]
  assign _T_855 = io_decode_0_csr == 12'hb16; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119048.4]
  assign _T_856 = io_decode_0_csr == 12'hb96; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119049.4]
  assign _T_857 = io_decode_0_csr == 12'h337; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119050.4]
  assign _T_858 = io_decode_0_csr == 12'hb17; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119051.4]
  assign _T_859 = io_decode_0_csr == 12'hb97; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119052.4]
  assign _T_860 = io_decode_0_csr == 12'h338; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119053.4]
  assign _T_861 = io_decode_0_csr == 12'hb18; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119054.4]
  assign _T_862 = io_decode_0_csr == 12'hb98; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119055.4]
  assign _T_863 = io_decode_0_csr == 12'h339; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119056.4]
  assign _T_864 = io_decode_0_csr == 12'hb19; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119057.4]
  assign _T_865 = io_decode_0_csr == 12'hb99; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119058.4]
  assign _T_866 = io_decode_0_csr == 12'h33a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119059.4]
  assign _T_867 = io_decode_0_csr == 12'hb1a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119060.4]
  assign _T_868 = io_decode_0_csr == 12'hb9a; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119061.4]
  assign _T_869 = io_decode_0_csr == 12'h33b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119062.4]
  assign _T_870 = io_decode_0_csr == 12'hb1b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119063.4]
  assign _T_871 = io_decode_0_csr == 12'hb9b; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119064.4]
  assign _T_872 = io_decode_0_csr == 12'h33c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119065.4]
  assign _T_873 = io_decode_0_csr == 12'hb1c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119066.4]
  assign _T_874 = io_decode_0_csr == 12'hb9c; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119067.4]
  assign _T_875 = io_decode_0_csr == 12'h33d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119068.4]
  assign _T_876 = io_decode_0_csr == 12'hb1d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119069.4]
  assign _T_877 = io_decode_0_csr == 12'hb9d; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119070.4]
  assign _T_878 = io_decode_0_csr == 12'h33e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119071.4]
  assign _T_879 = io_decode_0_csr == 12'hb1e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119072.4]
  assign _T_880 = io_decode_0_csr == 12'hb9e; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119073.4]
  assign _T_881 = io_decode_0_csr == 12'h33f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119074.4]
  assign _T_882 = io_decode_0_csr == 12'hb1f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119075.4]
  assign _T_883 = io_decode_0_csr == 12'hb9f; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119076.4]
  assign _T_884 = io_decode_0_csr == 12'hb80; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119077.4]
  assign _T_885 = io_decode_0_csr == 12'hb82; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119078.4]
  assign _T_886 = io_decode_0_csr == 12'h3a0; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119079.4]
  assign _T_887 = io_decode_0_csr == 12'h3a1; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119080.4]
  assign _T_888 = io_decode_0_csr == 12'h3a2; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119081.4]
  assign _T_889 = io_decode_0_csr == 12'h3a3; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119082.4]
  assign _T_890 = io_decode_0_csr == 12'h3b0; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119083.4]
  assign _T_891 = io_decode_0_csr == 12'h3b1; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119084.4]
  assign _T_892 = io_decode_0_csr == 12'h3b2; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119085.4]
  assign _T_893 = io_decode_0_csr == 12'h3b3; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119086.4]
  assign _T_894 = io_decode_0_csr == 12'h3b4; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119087.4]
  assign _T_895 = io_decode_0_csr == 12'h3b5; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119088.4]
  assign _T_896 = io_decode_0_csr == 12'h3b6; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119089.4]
  assign _T_897 = io_decode_0_csr == 12'h3b7; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119090.4]
  assign _T_898 = io_decode_0_csr == 12'h3b8; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119091.4]
  assign _T_899 = io_decode_0_csr == 12'h3b9; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119092.4]
  assign _T_900 = io_decode_0_csr == 12'h3ba; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119093.4]
  assign _T_901 = io_decode_0_csr == 12'h3bb; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119094.4]
  assign _T_902 = io_decode_0_csr == 12'h3bc; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119095.4]
  assign _T_903 = io_decode_0_csr == 12'h3bd; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119096.4]
  assign _T_904 = io_decode_0_csr == 12'h3be; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119097.4]
  assign _T_905 = io_decode_0_csr == 12'h3bf; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119098.4]
  assign _T_906 = io_decode_0_csr == 12'h7c1; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119099.4]
  assign _T_907 = io_decode_0_csr == 12'hf12; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119100.4]
  assign _T_908 = io_decode_0_csr == 12'hf11; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119101.4]
  assign _T_909 = io_decode_0_csr == 12'hf13; // @[CSR.scala 517:99:freechips.rocketchip.system.TinyConfig.fir@119102.4]
  assign _T_910 = _T_779 | _T_780; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119103.4]
  assign _T_911 = _T_910 | _T_781; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119104.4]
  assign _T_912 = _T_911 | _T_782; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119105.4]
  assign _T_913 = _T_912 | _T_783; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119106.4]
  assign _T_914 = _T_913 | _T_784; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119107.4]
  assign _T_915 = _T_914 | _T_785; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119108.4]
  assign _T_916 = _T_915 | _T_786; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119109.4]
  assign _T_917 = _T_916 | _T_787; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119110.4]
  assign _T_918 = _T_917 | _T_788; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119111.4]
  assign _T_919 = _T_918 | _T_789; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119112.4]
  assign _T_920 = _T_919 | _T_790; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119113.4]
  assign _T_921 = _T_920 | _T_791; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119114.4]
  assign _T_922 = _T_921 | _T_792; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119115.4]
  assign _T_923 = _T_922 | _T_793; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119116.4]
  assign _T_924 = _T_923 | _T_794; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119117.4]
  assign _T_925 = _T_924 | _T_795; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119118.4]
  assign _T_926 = _T_925 | _T_796; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119119.4]
  assign _T_927 = _T_926 | _T_797; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119120.4]
  assign _T_928 = _T_927 | _T_798; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119121.4]
  assign _T_929 = _T_928 | _T_799; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119122.4]
  assign _T_930 = _T_929 | _T_800; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119123.4]
  assign _T_931 = _T_930 | _T_801; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119124.4]
  assign _T_932 = _T_931 | _T_802; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119125.4]
  assign _T_933 = _T_932 | _T_803; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119126.4]
  assign _T_934 = _T_933 | _T_804; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119127.4]
  assign _T_935 = _T_934 | _T_805; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119128.4]
  assign _T_936 = _T_935 | _T_806; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119129.4]
  assign _T_937 = _T_936 | _T_807; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119130.4]
  assign _T_938 = _T_937 | _T_808; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119131.4]
  assign _T_939 = _T_938 | _T_809; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119132.4]
  assign _T_940 = _T_939 | _T_810; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119133.4]
  assign _T_941 = _T_940 | _T_811; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119134.4]
  assign _T_942 = _T_941 | _T_812; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119135.4]
  assign _T_943 = _T_942 | _T_813; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119136.4]
  assign _T_944 = _T_943 | _T_814; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119137.4]
  assign _T_945 = _T_944 | _T_815; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119138.4]
  assign _T_946 = _T_945 | _T_816; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119139.4]
  assign _T_947 = _T_946 | _T_817; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119140.4]
  assign _T_948 = _T_947 | _T_818; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119141.4]
  assign _T_949 = _T_948 | _T_819; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119142.4]
  assign _T_950 = _T_949 | _T_820; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119143.4]
  assign _T_951 = _T_950 | _T_821; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119144.4]
  assign _T_952 = _T_951 | _T_822; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119145.4]
  assign _T_953 = _T_952 | _T_823; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119146.4]
  assign _T_954 = _T_953 | _T_824; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119147.4]
  assign _T_955 = _T_954 | _T_825; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119148.4]
  assign _T_956 = _T_955 | _T_826; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119149.4]
  assign _T_957 = _T_956 | _T_827; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119150.4]
  assign _T_958 = _T_957 | _T_828; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119151.4]
  assign _T_959 = _T_958 | _T_829; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119152.4]
  assign _T_960 = _T_959 | _T_830; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119153.4]
  assign _T_961 = _T_960 | _T_831; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119154.4]
  assign _T_962 = _T_961 | _T_832; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119155.4]
  assign _T_963 = _T_962 | _T_833; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119156.4]
  assign _T_964 = _T_963 | _T_834; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119157.4]
  assign _T_965 = _T_964 | _T_835; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119158.4]
  assign _T_966 = _T_965 | _T_836; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119159.4]
  assign _T_967 = _T_966 | _T_837; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119160.4]
  assign _T_968 = _T_967 | _T_838; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119161.4]
  assign _T_969 = _T_968 | _T_839; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119162.4]
  assign _T_970 = _T_969 | _T_840; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119163.4]
  assign _T_971 = _T_970 | _T_841; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119164.4]
  assign _T_972 = _T_971 | _T_842; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119165.4]
  assign _T_973 = _T_972 | _T_843; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119166.4]
  assign _T_974 = _T_973 | _T_844; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119167.4]
  assign _T_975 = _T_974 | _T_845; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119168.4]
  assign _T_976 = _T_975 | _T_846; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119169.4]
  assign _T_977 = _T_976 | _T_847; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119170.4]
  assign _T_978 = _T_977 | _T_848; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119171.4]
  assign _T_979 = _T_978 | _T_849; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119172.4]
  assign _T_980 = _T_979 | _T_850; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119173.4]
  assign _T_981 = _T_980 | _T_851; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119174.4]
  assign _T_982 = _T_981 | _T_852; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119175.4]
  assign _T_983 = _T_982 | _T_853; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119176.4]
  assign _T_984 = _T_983 | _T_854; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119177.4]
  assign _T_985 = _T_984 | _T_855; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119178.4]
  assign _T_986 = _T_985 | _T_856; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119179.4]
  assign _T_987 = _T_986 | _T_857; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119180.4]
  assign _T_988 = _T_987 | _T_858; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119181.4]
  assign _T_989 = _T_988 | _T_859; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119182.4]
  assign _T_990 = _T_989 | _T_860; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119183.4]
  assign _T_991 = _T_990 | _T_861; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119184.4]
  assign _T_992 = _T_991 | _T_862; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119185.4]
  assign _T_993 = _T_992 | _T_863; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119186.4]
  assign _T_994 = _T_993 | _T_864; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119187.4]
  assign _T_995 = _T_994 | _T_865; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119188.4]
  assign _T_996 = _T_995 | _T_866; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119189.4]
  assign _T_997 = _T_996 | _T_867; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119190.4]
  assign _T_998 = _T_997 | _T_868; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119191.4]
  assign _T_999 = _T_998 | _T_869; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119192.4]
  assign _T_1000 = _T_999 | _T_870; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119193.4]
  assign _T_1001 = _T_1000 | _T_871; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119194.4]
  assign _T_1002 = _T_1001 | _T_872; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119195.4]
  assign _T_1003 = _T_1002 | _T_873; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119196.4]
  assign _T_1004 = _T_1003 | _T_874; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119197.4]
  assign _T_1005 = _T_1004 | _T_875; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119198.4]
  assign _T_1006 = _T_1005 | _T_876; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119199.4]
  assign _T_1007 = _T_1006 | _T_877; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119200.4]
  assign _T_1008 = _T_1007 | _T_878; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119201.4]
  assign _T_1009 = _T_1008 | _T_879; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119202.4]
  assign _T_1010 = _T_1009 | _T_880; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119203.4]
  assign _T_1011 = _T_1010 | _T_881; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119204.4]
  assign _T_1012 = _T_1011 | _T_882; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119205.4]
  assign _T_1013 = _T_1012 | _T_883; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119206.4]
  assign _T_1014 = _T_1013 | _T_884; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119207.4]
  assign _T_1015 = _T_1014 | _T_885; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119208.4]
  assign _T_1016 = _T_1015 | _T_886; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119209.4]
  assign _T_1017 = _T_1016 | _T_887; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119210.4]
  assign _T_1018 = _T_1017 | _T_888; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119211.4]
  assign _T_1019 = _T_1018 | _T_889; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119212.4]
  assign _T_1020 = _T_1019 | _T_890; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119213.4]
  assign _T_1021 = _T_1020 | _T_891; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119214.4]
  assign _T_1022 = _T_1021 | _T_892; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119215.4]
  assign _T_1023 = _T_1022 | _T_893; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119216.4]
  assign _T_1024 = _T_1023 | _T_894; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119217.4]
  assign _T_1025 = _T_1024 | _T_895; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119218.4]
  assign _T_1026 = _T_1025 | _T_896; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119219.4]
  assign _T_1027 = _T_1026 | _T_897; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119220.4]
  assign _T_1028 = _T_1027 | _T_898; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119221.4]
  assign _T_1029 = _T_1028 | _T_899; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119222.4]
  assign _T_1030 = _T_1029 | _T_900; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119223.4]
  assign _T_1031 = _T_1030 | _T_901; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119224.4]
  assign _T_1032 = _T_1031 | _T_902; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119225.4]
  assign _T_1033 = _T_1032 | _T_903; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119226.4]
  assign _T_1034 = _T_1033 | _T_904; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119227.4]
  assign _T_1035 = _T_1034 | _T_905; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119228.4]
  assign _T_1036 = _T_1035 | _T_906; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119229.4]
  assign _T_1037 = _T_1036 | _T_907; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119230.4]
  assign _T_1038 = _T_1037 | _T_908; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119231.4]
  assign _T_1039 = _T_1038 | _T_909; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119232.4]
  assign _T_1040 = _T_1039 == 1'h0; // @[CSR.scala 528:7:freechips.rocketchip.system.TinyConfig.fir@119233.4]
  assign _T_1059 = _T_792 | _T_793; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119252.4]
  assign _T_1060 = _T_1059 | _T_794; // @[CSR.scala 517:115:freechips.rocketchip.system.TinyConfig.fir@119253.4]
  assign _T_1062 = reg_debug == 1'h0; // @[CSR.scala 531:52:freechips.rocketchip.system.TinyConfig.fir@119255.4]
  assign _T_1063 = _T_1060 & _T_1062; // @[CSR.scala 531:49:freechips.rocketchip.system.TinyConfig.fir@119256.4]
  assign _T_1064 = _T_1040 | _T_1063; // @[CSR.scala 530:148:freechips.rocketchip.system.TinyConfig.fir@119257.4]
  assign _T_1065 = io_decode_0_fp_csr & io_decode_0_fp_illegal; // @[CSR.scala 532:21:freechips.rocketchip.system.TinyConfig.fir@119258.4]
  assign _T_1067 = io_decode_0_csr[11:10]; // @[CSR.scala 533:39:freechips.rocketchip.system.TinyConfig.fir@119261.4]
  assign _T_1069 = io_decode_0_csr >= 12'h340; // @[CSR.scala 534:40:freechips.rocketchip.system.TinyConfig.fir@119264.4]
  assign _T_1070 = io_decode_0_csr <= 12'h343; // @[CSR.scala 534:71:freechips.rocketchip.system.TinyConfig.fir@119265.4]
  assign _T_1071 = _T_1069 & _T_1070; // @[CSR.scala 534:57:freechips.rocketchip.system.TinyConfig.fir@119266.4]
  assign _T_1072 = io_decode_0_csr >= 12'h140; // @[CSR.scala 534:99:freechips.rocketchip.system.TinyConfig.fir@119267.4]
  assign _T_1073 = io_decode_0_csr <= 12'h143; // @[CSR.scala 534:130:freechips.rocketchip.system.TinyConfig.fir@119268.4]
  assign _T_1074 = _T_1072 & _T_1073; // @[CSR.scala 534:116:freechips.rocketchip.system.TinyConfig.fir@119269.4]
  assign _T_1075 = _T_1071 | _T_1074; // @[CSR.scala 534:85:freechips.rocketchip.system.TinyConfig.fir@119270.4]
  assign _T_1090 = insn_break ? 32'h3 : io_cause; // @[CSR.scala 543:14:freechips.rocketchip.system.TinyConfig.fir@119287.4]
  assign cause = insn_call ? 32'hb : _T_1090; // @[CSR.scala 542:8:freechips.rocketchip.system.TinyConfig.fir@119288.4]
  assign cause_lsbs = cause[7:0]; // @[CSR.scala 544:25:freechips.rocketchip.system.TinyConfig.fir@119289.4]
  assign _T_1091 = cause[31]; // @[CSR.scala 545:30:freechips.rocketchip.system.TinyConfig.fir@119290.4]
  assign _T_1092 = cause_lsbs == 8'he; // @[CSR.scala 545:53:freechips.rocketchip.system.TinyConfig.fir@119291.4]
  assign causeIsDebugInt = _T_1091 & _T_1092; // @[CSR.scala 545:39:freechips.rocketchip.system.TinyConfig.fir@119292.4]
  assign _T_1094 = _T_1091 == 1'h0; // @[CSR.scala 546:29:freechips.rocketchip.system.TinyConfig.fir@119294.4]
  assign causeIsDebugTrigger = _T_1094 & _T_1092; // @[CSR.scala 546:44:freechips.rocketchip.system.TinyConfig.fir@119296.4]
  assign _T_1098 = _T_1094 & insn_break; // @[CSR.scala 547:42:freechips.rocketchip.system.TinyConfig.fir@119299.4]
  assign _T_1101 = {reg_dcsr_ebreakm,1'h0,2'h0}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@119302.4]
  assign _GEN_421 = _T_1101[3:3]; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119303.4]
  assign _T_1102 = {{3'd0}, _GEN_421}; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119303.4]
  assign _T_1103 = _T_1102[0]; // @[CSR.scala 547:134:freechips.rocketchip.system.TinyConfig.fir@119304.4]
  assign causeIsDebugBreak = _T_1098 & _T_1103; // @[CSR.scala 547:56:freechips.rocketchip.system.TinyConfig.fir@119305.4]
  assign _T_1104 = reg_singleStepped | causeIsDebugInt; // @[CSR.scala 548:60:freechips.rocketchip.system.TinyConfig.fir@119306.4]
  assign _T_1105 = _T_1104 | causeIsDebugTrigger; // @[CSR.scala 548:79:freechips.rocketchip.system.TinyConfig.fir@119307.4]
  assign _T_1106 = _T_1105 | causeIsDebugBreak; // @[CSR.scala 548:102:freechips.rocketchip.system.TinyConfig.fir@119308.4]
  assign trapToDebug = _T_1106 | reg_debug; // @[CSR.scala 548:123:freechips.rocketchip.system.TinyConfig.fir@119309.4]
  assign _T_1108 = insn_break ? 12'h800 : 12'h808; // @[CSR.scala 549:37:freechips.rocketchip.system.TinyConfig.fir@119311.4]
  assign debugTVec = reg_debug ? _T_1108 : 12'h800; // @[CSR.scala 549:22:freechips.rocketchip.system.TinyConfig.fir@119312.4]
  assign _T_1118 = cause[4:0]; // @[CSR.scala 558:32:freechips.rocketchip.system.TinyConfig.fir@119323.4]
  assign _T_1119 = {_T_1118, 2'h0}; // @[CSR.scala 558:59:freechips.rocketchip.system.TinyConfig.fir@119324.4]
  assign _T_1120 = read_mtvec[31:7]; // @[CSR.scala 559:33:freechips.rocketchip.system.TinyConfig.fir@119325.4]
  assign _T_1121 = {_T_1120,_T_1119}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@119326.4]
  assign _T_1122 = read_mtvec[0]; // @[CSR.scala 560:24:freechips.rocketchip.system.TinyConfig.fir@119327.4]
  assign _T_1124 = _T_1122 & _T_1091; // @[CSR.scala 560:28:freechips.rocketchip.system.TinyConfig.fir@119329.4]
  assign _T_1125 = cause_lsbs[7:5]; // @[CSR.scala 560:70:freechips.rocketchip.system.TinyConfig.fir@119330.4]
  assign _T_1126 = _T_1125 == 3'h0; // @[CSR.scala 560:94:freechips.rocketchip.system.TinyConfig.fir@119331.4]
  assign _T_1127 = _T_1124 & _T_1126; // @[CSR.scala 560:55:freechips.rocketchip.system.TinyConfig.fir@119332.4]
  assign _T_1128 = read_mtvec[31:2]; // @[CSR.scala 561:38:freechips.rocketchip.system.TinyConfig.fir@119333.4]
  assign _T_1129 = {_T_1128, 2'h0}; // @[CSR.scala 561:56:freechips.rocketchip.system.TinyConfig.fir@119334.4]
  assign notDebugTVec = _T_1127 ? _T_1121 : _T_1129; // @[CSR.scala 561:8:freechips.rocketchip.system.TinyConfig.fir@119335.4]
  assign tvec = trapToDebug ? {{20'd0}, debugTVec} : notDebugTVec; // @[CSR.scala 563:17:freechips.rocketchip.system.TinyConfig.fir@119336.4]
  assign _T_1130 = insn_call | insn_break; // @[CSR.scala 566:24:freechips.rocketchip.system.TinyConfig.fir@119339.4]
  assign _T_1134 = io_status_fs == 2'h3; // @[CSR.scala 569:32:freechips.rocketchip.system.TinyConfig.fir@119346.4]
  assign _T_1135 = io_status_xs == 2'h3; // @[CSR.scala 569:53:freechips.rocketchip.system.TinyConfig.fir@119347.4]
  assign exception = _T_1130 | io_exception; // @[CSR.scala 578:43:freechips.rocketchip.system.TinyConfig.fir@119362.4]
  assign _T_1142 = insn_ret + insn_call; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119363.4]
  assign _T_1144 = insn_break + io_exception; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119365.4]
  assign _T_1146 = _T_1142 + _T_1144; // @[Bitwise.scala 48:55:freechips.rocketchip.system.TinyConfig.fir@119367.4]
  assign _T_1148 = _T_1146 <= 3'h1; // @[CSR.scala 579:79:freechips.rocketchip.system.TinyConfig.fir@119369.4]
  assign _T_1150 = _T_1148 | reset; // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119371.4]
  assign _T_1151 = _T_1150 == 1'h0; // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119372.4]
  assign _T_1153 = insn_wfi & _T_273; // @[CSR.scala 581:18:freechips.rocketchip.system.TinyConfig.fir@119378.4]
  assign _T_1155 = _T_1153 & _T_1062; // @[CSR.scala 581:36:freechips.rocketchip.system.TinyConfig.fir@119380.4]
  assign _T_1156 = pending_interrupts != 32'h0; // @[CSR.scala 582:28:freechips.rocketchip.system.TinyConfig.fir@119384.4]
  assign _T_1157 = _T_1156 | io_interrupts_debug; // @[CSR.scala 582:32:freechips.rocketchip.system.TinyConfig.fir@119385.4]
  assign _T_1158 = _T_1157 | exception; // @[CSR.scala 582:55:freechips.rocketchip.system.TinyConfig.fir@119386.4]
  assign _T_1160 = io_retire | exception; // @[CSR.scala 584:22:freechips.rocketchip.system.TinyConfig.fir@119391.4]
  assign _T_1168 = reg_singleStepped == 1'h0; // @[CSR.scala 587:10:freechips.rocketchip.system.TinyConfig.fir@119409.4]
  assign _T_1169 = io_retire == 1'h0; // @[CSR.scala 587:42:freechips.rocketchip.system.TinyConfig.fir@119410.4]
  assign _T_1170 = _T_1168 | _T_1169; // @[CSR.scala 587:29:freechips.rocketchip.system.TinyConfig.fir@119411.4]
  assign _T_1172 = _T_1170 | reset; // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119413.4]
  assign _T_1173 = _T_1172 == 1'h0; // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119414.4]
  assign _T_1174 = ~ io_pc; // @[CSR.scala 934:28:freechips.rocketchip.system.TinyConfig.fir@119419.4]
  assign _T_1175 = _T_1174 | 32'h1; // @[CSR.scala 934:31:freechips.rocketchip.system.TinyConfig.fir@119420.4]
  assign epc = ~ _T_1175; // @[CSR.scala 934:26:freechips.rocketchip.system.TinyConfig.fir@119421.4]
  assign _T_1177 = causeIsDebugTrigger ? 2'h2 : 2'h1; // @[CSR.scala 598:86:freechips.rocketchip.system.TinyConfig.fir@119431.10]
  assign _T_1178 = causeIsDebugInt ? 2'h3 : _T_1177; // @[CSR.scala 598:56:freechips.rocketchip.system.TinyConfig.fir@119432.10]
  assign _GEN_48 = {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 602:27:freechips.rocketchip.system.TinyConfig.fir@119440.8]
  assign _GEN_67 = trapToDebug ? {{1'd0}, reg_mstatus_spp} : _GEN_48; // @[CSR.scala 594:24:freechips.rocketchip.system.TinyConfig.fir@119426.6]
  assign _GEN_85 = exception ? _GEN_67 : {{1'd0}, reg_mstatus_spp}; // @[CSR.scala 593:20:freechips.rocketchip.system.TinyConfig.fir@119425.4]
  assign _T_1468 = io_rw_addr[10]; // @[CSR.scala 649:47:freechips.rocketchip.system.TinyConfig.fir@119758.8]
  assign _GEN_95 = _T_1468 ? _T_426 : _T_408; // @[CSR.scala 649:53:freechips.rocketchip.system.TinyConfig.fir@119760.8]
  assign _T_1483 = _T_562 ? _T_403 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119804.4]
  assign _T_1484 = _T_563 ? reg_bp_0_address : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119805.4]
  assign _T_1485 = _T_564 ? reg_misa : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119806.4]
  assign _T_1486 = _T_565 ? read_mstatus : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119807.4]
  assign _T_1487 = _T_566 ? read_mtvec : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119808.4]
  assign _T_1488 = _T_567 ? read_mip : 16'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119809.4]
  assign _T_1489 = _T_568 ? reg_mie : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119810.4]
  assign _T_1490 = _T_569 ? reg_mscratch : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119811.4]
  assign _T_1491 = _T_570 ? _T_408 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119812.4]
  assign _T_1492 = _T_571 ? reg_mtval : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119813.4]
  assign _T_1493 = _T_572 ? reg_mcause : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119814.4]
  assign _T_1495 = _T_574 ? _T_421 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119816.4]
  assign _T_1496 = _T_575 ? _T_426 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119817.4]
  assign _T_1497 = _T_576 ? reg_dscratch : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119818.4]
  assign _T_1498 = _T_577 ? _T_97 : 64'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119819.4]
  assign _T_1499 = _T_578 ? _T_89 : 64'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119820.4]
  assign _T_1587 = _T_666 ? _T_457 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119908.4]
  assign _T_1588 = _T_667 ? _T_458 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119909.4]
  assign _T_1589 = _T_668 ? _T_491 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119910.4]
  assign _T_1590 = _T_669 ? _T_514 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119911.4]
  assign _T_1593 = _T_672 ? reg_pmp_0_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119914.4]
  assign _T_1594 = _T_673 ? reg_pmp_1_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119915.4]
  assign _T_1595 = _T_674 ? reg_pmp_2_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119916.4]
  assign _T_1596 = _T_675 ? reg_pmp_3_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119917.4]
  assign _T_1597 = _T_676 ? reg_pmp_4_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119918.4]
  assign _T_1598 = _T_677 ? reg_pmp_5_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119919.4]
  assign _T_1599 = _T_678 ? reg_pmp_6_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119920.4]
  assign _T_1600 = _T_679 ? reg_pmp_7_addr : 30'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119921.4]
  assign _T_1610 = _T_689 ? 32'h1 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119931.4]
  assign _T_1612 = _T_691 ? 32'h20181004 : 32'h0; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119933.4]
  assign _T_1614 = _T_1483 | _T_1484; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119935.4]
  assign _T_1615 = _T_1614 | _T_1485; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119936.4]
  assign _T_1616 = _T_1615 | _T_1486; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119937.4]
  assign _T_1617 = _T_1616 | _T_1487; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119938.4]
  assign _GEN_424 = {{16'd0}, _T_1488}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119939.4]
  assign _T_1618 = _T_1617 | _GEN_424; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119939.4]
  assign _T_1619 = _T_1618 | _T_1489; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119940.4]
  assign _T_1620 = _T_1619 | _T_1490; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119941.4]
  assign _T_1621 = _T_1620 | _T_1491; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119942.4]
  assign _T_1622 = _T_1621 | _T_1492; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119943.4]
  assign _T_1623 = _T_1622 | _T_1493; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119944.4]
  assign _T_1625 = _T_1623 | _T_1495; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119946.4]
  assign _T_1626 = _T_1625 | _T_1496; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119947.4]
  assign _T_1627 = _T_1626 | _T_1497; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119948.4]
  assign _GEN_425 = {{32'd0}, _T_1627}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119949.4]
  assign _T_1628 = _GEN_425 | _T_1498; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119949.4]
  assign _T_1629 = _T_1628 | _T_1499; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@119950.4]
  assign _GEN_426 = {{32'd0}, _T_1587}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120038.4]
  assign _T_1717 = _T_1629 | _GEN_426; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120038.4]
  assign _GEN_427 = {{32'd0}, _T_1588}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120039.4]
  assign _T_1718 = _T_1717 | _GEN_427; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120039.4]
  assign _GEN_428 = {{32'd0}, _T_1589}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120040.4]
  assign _T_1719 = _T_1718 | _GEN_428; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120040.4]
  assign _GEN_429 = {{32'd0}, _T_1590}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120041.4]
  assign _T_1720 = _T_1719 | _GEN_429; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120041.4]
  assign _GEN_430 = {{34'd0}, _T_1593}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120044.4]
  assign _T_1723 = _T_1720 | _GEN_430; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120044.4]
  assign _GEN_431 = {{34'd0}, _T_1594}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120045.4]
  assign _T_1724 = _T_1723 | _GEN_431; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120045.4]
  assign _GEN_432 = {{34'd0}, _T_1595}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120046.4]
  assign _T_1725 = _T_1724 | _GEN_432; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120046.4]
  assign _GEN_433 = {{34'd0}, _T_1596}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120047.4]
  assign _T_1726 = _T_1725 | _GEN_433; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120047.4]
  assign _GEN_434 = {{34'd0}, _T_1597}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120048.4]
  assign _T_1727 = _T_1726 | _GEN_434; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120048.4]
  assign _GEN_435 = {{34'd0}, _T_1598}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120049.4]
  assign _T_1728 = _T_1727 | _GEN_435; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120049.4]
  assign _GEN_436 = {{34'd0}, _T_1599}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120050.4]
  assign _T_1729 = _T_1728 | _GEN_436; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120050.4]
  assign _GEN_437 = {{34'd0}, _T_1600}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120051.4]
  assign _T_1730 = _T_1729 | _GEN_437; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120051.4]
  assign _GEN_438 = {{32'd0}, _T_1610}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120061.4]
  assign _T_1740 = _T_1730 | _GEN_438; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120061.4]
  assign _GEN_439 = {{32'd0}, _T_1612}; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120063.4]
  assign _T_1742 = _T_1740 | _GEN_439; // @[Mux.scala 28:72:freechips.rocketchip.system.TinyConfig.fir@120063.4]
  assign _T_1746 = io_rw_cmd == 3'h5; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120070.6]
  assign _T_1747 = io_rw_cmd == 3'h6; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120071.6]
  assign _T_1748 = io_rw_cmd == 3'h7; // @[package.scala 15:47:freechips.rocketchip.system.TinyConfig.fir@120072.6]
  assign _T_3320 = _T_1747 | _T_1748; // @[package.scala 15:62:freechips.rocketchip.system.TinyConfig.fir@122175.4]
  assign csr_wen = _T_3320 | _T_1746; // @[package.scala 15:62:freechips.rocketchip.system.TinyConfig.fir@122176.4]
  assign _T_3334 = {{70'd0}, wdata}; // @[:freechips.rocketchip.system.TinyConfig.fir@122194.8 :freechips.rocketchip.system.TinyConfig.fir@122196.8]
  assign _T_3338 = _T_3334[3]; // @[CSR.scala 701:47:freechips.rocketchip.system.TinyConfig.fir@122203.8]
  assign _T_3342 = _T_3334[7]; // @[CSR.scala 701:47:freechips.rocketchip.system.TinyConfig.fir@122211.8]
  assign _T_3365 = wdata[5]; // @[CSR.scala 725:20:freechips.rocketchip.system.TinyConfig.fir@122261.8]
  assign _T_3366 = io_pc[1]; // @[CSR.scala 727:39:freechips.rocketchip.system.TinyConfig.fir@122262.8]
  assign _T_3367 = _T_3366 == 1'h0; // @[CSR.scala 727:33:freechips.rocketchip.system.TinyConfig.fir@122263.8]
  assign _T_3369 = wdata[2]; // @[CSR.scala 727:51:freechips.rocketchip.system.TinyConfig.fir@122265.8]
  assign _T_3370 = _T_3367 | _T_3369; // @[CSR.scala 727:43:freechips.rocketchip.system.TinyConfig.fir@122266.8]
  assign _T_3371 = ~ wdata; // @[CSR.scala 729:25:freechips.rocketchip.system.TinyConfig.fir@122268.10]
  assign _T_3372 = _T_3365 == 1'h0; // @[CSR.scala 729:35:freechips.rocketchip.system.TinyConfig.fir@122269.10]
  assign _T_3373 = {_T_3372, 3'h0}; // @[CSR.scala 729:38:freechips.rocketchip.system.TinyConfig.fir@122270.10]
  assign _GEN_440 = {{28'd0}, _T_3373}; // @[CSR.scala 729:32:freechips.rocketchip.system.TinyConfig.fir@122271.10]
  assign _T_3374 = _T_3371 | _GEN_440; // @[CSR.scala 729:32:freechips.rocketchip.system.TinyConfig.fir@122271.10]
  assign _T_3375 = ~ _T_3374; // @[CSR.scala 729:23:freechips.rocketchip.system.TinyConfig.fir@122272.10]
  assign _T_3376 = _T_3375 & 32'h1005; // @[CSR.scala 729:55:freechips.rocketchip.system.TinyConfig.fir@122273.10]
  assign _T_3378 = reg_misa & 32'hffffeffa; // @[CSR.scala 729:73:freechips.rocketchip.system.TinyConfig.fir@122275.10]
  assign _T_3379 = _T_3376 | _T_3378; // @[CSR.scala 729:62:freechips.rocketchip.system.TinyConfig.fir@122276.10]
  assign _T_3421 = wdata & 32'h888; // @[CSR.scala 744:59:freechips.rocketchip.system.TinyConfig.fir@122343.8]
  assign _T_3423 = _T_3371 | 32'h1; // @[CSR.scala 934:31:freechips.rocketchip.system.TinyConfig.fir@122348.8]
  assign _T_3424 = ~ _T_3423; // @[CSR.scala 934:26:freechips.rocketchip.system.TinyConfig.fir@122349.8]
  assign _T_3425 = wdata & 32'h8000000f; // @[CSR.scala 749:62:freechips.rocketchip.system.TinyConfig.fir@122359.8]
  assign _T_3427 = _T_97[63:32]; // @[CSR.scala 928:47:freechips.rocketchip.system.TinyConfig.fir@122367.8]
  assign _T_3428 = {_T_3427,wdata}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122368.8]
  assign _T_3429 = _T_3428[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122370.8]
  assign _GEN_130 = _T_577 ? _T_3428 : {{57'd0}, _T_92}; // @[CSR.scala 928:31:freechips.rocketchip.system.TinyConfig.fir@122366.6]
  assign _T_3431 = _T_97[31:0]; // @[CSR.scala 929:74:freechips.rocketchip.system.TinyConfig.fir@122375.8]
  assign _T_3432 = {wdata,_T_3431}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122376.8]
  assign _T_3433 = _T_3432[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122378.8]
  assign _GEN_132 = _T_666 ? _T_3432 : _GEN_130; // @[CSR.scala 929:31:freechips.rocketchip.system.TinyConfig.fir@122373.6]
  assign _T_3434 = _T_89[63:32]; // @[CSR.scala 928:47:freechips.rocketchip.system.TinyConfig.fir@122382.8]
  assign _T_3435 = {_T_3434,wdata}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122383.8]
  assign _T_3436 = _T_3435[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122385.8]
  assign _GEN_134 = _T_578 ? _T_3435 : {{57'd0}, _T_84}; // @[CSR.scala 928:31:freechips.rocketchip.system.TinyConfig.fir@122381.6]
  assign _T_3438 = _T_89[31:0]; // @[CSR.scala 929:74:freechips.rocketchip.system.TinyConfig.fir@122390.8]
  assign _T_3439 = {wdata,_T_3438}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@122391.8]
  assign _T_3440 = _T_3439[63:6]; // @[Counters.scala 67:28:freechips.rocketchip.system.TinyConfig.fir@122393.8]
  assign _GEN_136 = _T_667 ? _T_3439 : _GEN_134; // @[CSR.scala 929:31:freechips.rocketchip.system.TinyConfig.fir@122388.6]
  assign _T_3453 = wdata[15]; // @[CSR.scala 768:43:freechips.rocketchip.system.TinyConfig.fir@122422.8]
  assign _T_3461 = reg_bp_0_control_dmode == 1'h0; // @[CSR.scala 819:37:freechips.rocketchip.system.TinyConfig.fir@122446.6]
  assign _T_3462 = _T_3461 | reg_debug; // @[CSR.scala 819:55:freechips.rocketchip.system.TinyConfig.fir@122447.6]
  assign _T_3466 = wdata[0]; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122459.10]
  assign _T_3467 = wdata[1]; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122461.10]
  assign _T_3473 = wdata[8:7]; // @[CSR.scala 822:41:freechips.rocketchip.system.TinyConfig.fir@122473.10]
  assign _T_3496 = _T_692 ? _T_403 : 32'h0; // @[CSR.scala 913:9:freechips.rocketchip.system.TinyConfig.fir@122505.10]
  assign _T_3497 = _T_3496 | io_rw_wdata; // @[CSR.scala 913:34:freechips.rocketchip.system.TinyConfig.fir@122506.10]
  assign _T_3502 = _T_3497 & _T_698; // @[CSR.scala 913:43:freechips.rocketchip.system.TinyConfig.fir@122511.10]
  assign _T_3515 = _T_3502[12]; // @[CSR.scala 828:96:freechips.rocketchip.system.TinyConfig.fir@122537.10]
  assign _T_3518 = _T_3502[27]; // @[CSR.scala 828:96:freechips.rocketchip.system.TinyConfig.fir@122543.10]
  assign _T_3520 = _T_3518 & reg_debug; // @[CSR.scala 829:38:freechips.rocketchip.system.TinyConfig.fir@122547.10]
  assign _T_3604 = reg_pmp_0_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122693.6]
  assign _T_3605 = _T_668 & _T_3604; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122694.6]
  assign _T_3608 = wdata[7:0]; // @[:freechips.rocketchip.system.TinyConfig.fir@122699.8 :freechips.rocketchip.system.TinyConfig.fir@122701.8]
  assign _T_3609 = _T_3608[0]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122702.8]
  assign _T_3610 = _T_3608[1]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122704.8]
  assign _T_3611 = _T_3608[2]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122706.8]
  assign _T_3612 = _T_3608[4:3]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122708.8]
  assign _T_3614 = _T_3608[7]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122712.8]
  assign _T_3615 = _T_3610 & _T_3609; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122715.8]
  assign _T_3616 = reg_pmp_1_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122718.6]
  assign _T_3617 = _T_3616 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122719.6]
  assign _T_3619 = _T_3617 & _T_289; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122721.6]
  assign _T_3620 = reg_pmp_1_cfg_l & _T_3619; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122722.6]
  assign _T_3621 = reg_pmp_0_cfg_l | _T_3620; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122723.6]
  assign _T_3622 = _T_3621 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122724.6]
  assign _T_3623 = _T_672 & _T_3622; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122725.6]
  assign _GEN_215 = _T_3623 ? wdata : {{2'd0}, reg_pmp_0_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122726.6]
  assign _T_3624 = reg_pmp_1_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122729.6]
  assign _T_3625 = _T_668 & _T_3624; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122730.6]
  assign _T_3626 = wdata[31:8]; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122732.8]
  assign _T_3628 = _T_3626[7:0]; // @[:freechips.rocketchip.system.TinyConfig.fir@122735.8 :freechips.rocketchip.system.TinyConfig.fir@122737.8]
  assign _T_3629 = _T_3628[0]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122738.8]
  assign _T_3630 = _T_3628[1]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122740.8]
  assign _T_3631 = _T_3628[2]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122742.8]
  assign _T_3632 = _T_3628[4:3]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122744.8]
  assign _T_3634 = _T_3628[7]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122748.8]
  assign _T_3635 = _T_3630 & _T_3629; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122751.8]
  assign _T_3636 = reg_pmp_2_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122754.6]
  assign _T_3637 = _T_3636 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122755.6]
  assign _T_3639 = _T_3637 & _T_298; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122757.6]
  assign _T_3640 = reg_pmp_2_cfg_l & _T_3639; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122758.6]
  assign _T_3641 = reg_pmp_1_cfg_l | _T_3640; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122759.6]
  assign _T_3642 = _T_3641 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122760.6]
  assign _T_3643 = _T_673 & _T_3642; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122761.6]
  assign _GEN_222 = _T_3643 ? wdata : {{2'd0}, reg_pmp_1_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122762.6]
  assign _T_3644 = reg_pmp_2_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122765.6]
  assign _T_3645 = _T_668 & _T_3644; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122766.6]
  assign _T_3646 = wdata[31:16]; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122768.8]
  assign _T_3648 = _T_3646[7:0]; // @[:freechips.rocketchip.system.TinyConfig.fir@122771.8 :freechips.rocketchip.system.TinyConfig.fir@122773.8]
  assign _T_3649 = _T_3648[0]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122774.8]
  assign _T_3650 = _T_3648[1]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122776.8]
  assign _T_3651 = _T_3648[2]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122778.8]
  assign _T_3652 = _T_3648[4:3]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122780.8]
  assign _T_3654 = _T_3648[7]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122784.8]
  assign _T_3655 = _T_3650 & _T_3649; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122787.8]
  assign _T_3656 = reg_pmp_3_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122790.6]
  assign _T_3657 = _T_3656 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122791.6]
  assign _T_3659 = _T_3657 & _T_307; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122793.6]
  assign _T_3660 = reg_pmp_3_cfg_l & _T_3659; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122794.6]
  assign _T_3661 = reg_pmp_2_cfg_l | _T_3660; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122795.6]
  assign _T_3662 = _T_3661 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122796.6]
  assign _T_3663 = _T_674 & _T_3662; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122797.6]
  assign _GEN_229 = _T_3663 ? wdata : {{2'd0}, reg_pmp_2_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122798.6]
  assign _T_3664 = reg_pmp_3_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122801.6]
  assign _T_3665 = _T_668 & _T_3664; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122802.6]
  assign _T_3666 = wdata[31:24]; // @[CSR.scala 840:53:freechips.rocketchip.system.TinyConfig.fir@122804.8]
  assign _T_3669 = _T_3666[0]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122810.8]
  assign _T_3670 = _T_3666[1]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122812.8]
  assign _T_3671 = _T_3666[2]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122814.8]
  assign _T_3672 = _T_3666[4:3]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122816.8]
  assign _T_3674 = _T_3666[7]; // @[CSR.scala 840:46:freechips.rocketchip.system.TinyConfig.fir@122820.8]
  assign _T_3675 = _T_3670 & _T_3669; // @[CSR.scala 843:31:freechips.rocketchip.system.TinyConfig.fir@122823.8]
  assign _T_3676 = reg_pmp_4_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122826.6]
  assign _T_3677 = _T_3676 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122827.6]
  assign _T_3679 = _T_3677 & _T_316; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122829.6]
  assign _T_3680 = reg_pmp_4_cfg_l & _T_3679; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122830.6]
  assign _T_3681 = reg_pmp_3_cfg_l | _T_3680; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122831.6]
  assign _T_3682 = _T_3681 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122832.6]
  assign _T_3683 = _T_675 & _T_3682; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122833.6]
  assign _GEN_236 = _T_3683 ? wdata : {{2'd0}, reg_pmp_3_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122834.6]
  assign _T_3684 = reg_pmp_4_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122837.6]
  assign _T_3685 = _T_669 & _T_3684; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122838.6]
  assign _T_3696 = reg_pmp_5_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122862.6]
  assign _T_3697 = _T_3696 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122863.6]
  assign _T_3699 = _T_3697 & _T_325; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122865.6]
  assign _T_3700 = reg_pmp_5_cfg_l & _T_3699; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122866.6]
  assign _T_3701 = reg_pmp_4_cfg_l | _T_3700; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122867.6]
  assign _T_3702 = _T_3701 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122868.6]
  assign _T_3703 = _T_676 & _T_3702; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122869.6]
  assign _GEN_243 = _T_3703 ? wdata : {{2'd0}, reg_pmp_4_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122870.6]
  assign _T_3704 = reg_pmp_5_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122873.6]
  assign _T_3705 = _T_669 & _T_3704; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122874.6]
  assign _T_3716 = reg_pmp_6_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122898.6]
  assign _T_3717 = _T_3716 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122899.6]
  assign _T_3719 = _T_3717 & _T_334; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122901.6]
  assign _T_3720 = reg_pmp_6_cfg_l & _T_3719; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122902.6]
  assign _T_3721 = reg_pmp_5_cfg_l | _T_3720; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122903.6]
  assign _T_3722 = _T_3721 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122904.6]
  assign _T_3723 = _T_677 & _T_3722; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122905.6]
  assign _GEN_250 = _T_3723 ? wdata : {{2'd0}, reg_pmp_5_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122906.6]
  assign _T_3724 = reg_pmp_6_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122909.6]
  assign _T_3725 = _T_669 & _T_3724; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122910.6]
  assign _T_3736 = reg_pmp_7_cfg_a[1]; // @[PMP.scala 45:20:freechips.rocketchip.system.TinyConfig.fir@122934.6]
  assign _T_3737 = _T_3736 == 1'h0; // @[PMP.scala 47:13:freechips.rocketchip.system.TinyConfig.fir@122935.6]
  assign _T_3739 = _T_3737 & _T_343; // @[PMP.scala 47:20:freechips.rocketchip.system.TinyConfig.fir@122937.6]
  assign _T_3740 = reg_pmp_7_cfg_l & _T_3739; // @[PMP.scala 49:62:freechips.rocketchip.system.TinyConfig.fir@122938.6]
  assign _T_3741 = reg_pmp_6_cfg_l | _T_3740; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122939.6]
  assign _T_3742 = _T_3741 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122940.6]
  assign _T_3743 = _T_678 & _T_3742; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122941.6]
  assign _GEN_257 = _T_3743 ? wdata : {{2'd0}, reg_pmp_6_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122942.6]
  assign _T_3744 = reg_pmp_7_cfg_l == 1'h0; // @[CSR.scala 839:60:freechips.rocketchip.system.TinyConfig.fir@122945.6]
  assign _T_3745 = _T_669 & _T_3744; // @[CSR.scala 839:57:freechips.rocketchip.system.TinyConfig.fir@122946.6]
  assign _T_3761 = reg_pmp_7_cfg_l | _T_3740; // @[PMP.scala 49:44:freechips.rocketchip.system.TinyConfig.fir@122975.6]
  assign _T_3762 = _T_3761 == 1'h0; // @[CSR.scala 848:48:freechips.rocketchip.system.TinyConfig.fir@122976.6]
  assign _T_3763 = _T_679 & _T_3762; // @[CSR.scala 848:45:freechips.rocketchip.system.TinyConfig.fir@122977.6]
  assign _GEN_264 = _T_3763 ? wdata : {{2'd0}, reg_pmp_7_addr}; // @[CSR.scala 848:71:freechips.rocketchip.system.TinyConfig.fir@122978.6]
  assign _GEN_282 = csr_wen ? _GEN_132 : {{57'd0}, _T_92}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_284 = csr_wen ? _GEN_136 : {{57'd0}, _T_84}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_329 = csr_wen ? _GEN_215 : {{2'd0}, reg_pmp_0_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_336 = csr_wen ? _GEN_222 : {{2'd0}, reg_pmp_1_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_343 = csr_wen ? _GEN_229 : {{2'd0}, reg_pmp_2_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_350 = csr_wen ? _GEN_236 : {{2'd0}, reg_pmp_3_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_357 = csr_wen ? _GEN_243 : {{2'd0}, reg_pmp_4_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_364 = csr_wen ? _GEN_250 : {{2'd0}, reg_pmp_5_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_371 = csr_wen ? _GEN_257 : {{2'd0}, reg_pmp_6_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _GEN_378 = csr_wen ? _GEN_264 : {{2'd0}, reg_pmp_7_addr}; // @[CSR.scala 699:18:freechips.rocketchip.system.TinyConfig.fir@122190.4]
  assign _T_3810 = io_retire > 1'h0; // @[CSR.scala 892:26:freechips.rocketchip.system.TinyConfig.fir@123141.4]
  assign io_rw_rdata = _T_1742[31:0]; // @[CSR.scala 672:15:freechips.rocketchip.system.TinyConfig.fir@120066.4]
  assign io_decode_0_fp_illegal = _T_764 | _T_766; // @[CSR.scala 524:23:freechips.rocketchip.system.TinyConfig.fir@118958.4]
  assign io_decode_0_fp_csr = 1'h0; // @[CSR.scala 525:19:freechips.rocketchip.system.TinyConfig.fir@118964.4]
  assign io_decode_0_read_illegal = _T_1064 | _T_1065; // @[CSR.scala 527:25:freechips.rocketchip.system.TinyConfig.fir@119260.4]
  assign io_decode_0_write_illegal = _T_1067 == 2'h3; // @[CSR.scala 533:26:freechips.rocketchip.system.TinyConfig.fir@119263.4]
  assign io_decode_0_write_flush = _T_1075 == 1'h0; // @[CSR.scala 534:24:freechips.rocketchip.system.TinyConfig.fir@119272.4]
  assign io_csr_stall = reg_wfi | io_status_cease; // @[CSR.scala 663:16:freechips.rocketchip.system.TinyConfig.fir@119785.4]
  assign io_eret = _T_1130 | insn_ret; // @[CSR.scala 566:11:freechips.rocketchip.system.TinyConfig.fir@119341.4]
  assign io_singleStep = reg_dcsr_step & _T_1062; // @[CSR.scala 567:17:freechips.rocketchip.system.TinyConfig.fir@119344.4]
  assign io_status_debug = reg_debug; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 570:19:freechips.rocketchip.system.TinyConfig.fir@119350.4]
  assign io_status_cease = _T_1481; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 664:19:freechips.rocketchip.system.TinyConfig.fir@119790.4]
  assign io_status_isa = reg_misa; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 571:17:freechips.rocketchip.system.TinyConfig.fir@119351.4]
  assign io_status_dprv = 2'h3; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 574:18:freechips.rocketchip.system.TinyConfig.fir@119359.4]
  assign io_status_prv = 2'h3; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_sd = _T_1134 | _T_1135; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 569:16:freechips.rocketchip.system.TinyConfig.fir@119349.4]
  assign io_status_zero2 = 27'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_sxl = 2'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 573:17:freechips.rocketchip.system.TinyConfig.fir@119353.4]
  assign io_status_uxl = 2'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 572:17:freechips.rocketchip.system.TinyConfig.fir@119352.4]
  assign io_status_sd_rv32 = io_status_sd; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4 CSR.scala 576:23:freechips.rocketchip.system.TinyConfig.fir@119360.4]
  assign io_status_zero1 = 8'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_tsr = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_tw = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_tvm = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_mxr = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_sum = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_xs = 2'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_fs = 2'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_hpp = 2'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_spp = reg_mstatus_spp; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_hpie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_spie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_upie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_hie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_sie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_status_uie = 1'h0; // @[CSR.scala 568:13:freechips.rocketchip.system.TinyConfig.fir@119345.4]
  assign io_evec = insn_ret ? _GEN_95 : tvec; // @[CSR.scala 564:11:freechips.rocketchip.system.TinyConfig.fir@119337.4 CSR.scala 648:15:freechips.rocketchip.system.TinyConfig.fir@119755.8 CSR.scala 652:15:freechips.rocketchip.system.TinyConfig.fir@119768.10 CSR.scala 658:15:freechips.rocketchip.system.TinyConfig.fir@119780.10]
  assign io_time = _T_97[31:0]; // @[CSR.scala 662:11:freechips.rocketchip.system.TinyConfig.fir@119783.4]
  assign io_interrupt = _T_275 & _T_277; // @[CSR.scala 361:16:freechips.rocketchip.system.TinyConfig.fir@118407.4]
  assign io_interrupt_cause = 32'h80000000 + _GEN_418; // @[CSR.scala 362:22:freechips.rocketchip.system.TinyConfig.fir@118408.4]
  assign io_bp_0_control_action = reg_bp_0_control_action; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_bp_0_control_tmatch = reg_bp_0_control_tmatch; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_bp_0_control_x = reg_bp_0_control_x; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_bp_0_control_w = reg_bp_0_control_w; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_bp_0_control_r = reg_bp_0_control_r; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_bp_0_address = reg_bp_0_address; // @[CSR.scala 363:9:freechips.rocketchip.system.TinyConfig.fir@118409.4]
  assign io_pmp_0_cfg_l = reg_pmp_0_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_cfg_a = reg_pmp_0_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_cfg_x = reg_pmp_0_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_cfg_w = reg_pmp_0_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_cfg_r = reg_pmp_0_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_addr = reg_pmp_0_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_0_mask = _T_287[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118506.4]
  assign io_pmp_1_cfg_l = reg_pmp_1_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_cfg_a = reg_pmp_1_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_cfg_x = reg_pmp_1_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_cfg_w = reg_pmp_1_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_cfg_r = reg_pmp_1_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_addr = reg_pmp_1_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_1_mask = _T_296[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118507.4]
  assign io_pmp_2_cfg_l = reg_pmp_2_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_cfg_a = reg_pmp_2_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_cfg_x = reg_pmp_2_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_cfg_w = reg_pmp_2_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_cfg_r = reg_pmp_2_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_addr = reg_pmp_2_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_2_mask = _T_305[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118508.4]
  assign io_pmp_3_cfg_l = reg_pmp_3_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_cfg_a = reg_pmp_3_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_cfg_x = reg_pmp_3_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_cfg_w = reg_pmp_3_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_cfg_r = reg_pmp_3_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_addr = reg_pmp_3_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_3_mask = _T_314[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118509.4]
  assign io_pmp_4_cfg_l = reg_pmp_4_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_cfg_a = reg_pmp_4_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_cfg_x = reg_pmp_4_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_cfg_w = reg_pmp_4_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_cfg_r = reg_pmp_4_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_addr = reg_pmp_4_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_4_mask = _T_323[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118510.4]
  assign io_pmp_5_cfg_l = reg_pmp_5_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_cfg_a = reg_pmp_5_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_cfg_x = reg_pmp_5_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_cfg_w = reg_pmp_5_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_cfg_r = reg_pmp_5_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_addr = reg_pmp_5_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_5_mask = _T_332[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118511.4]
  assign io_pmp_6_cfg_l = reg_pmp_6_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_cfg_a = reg_pmp_6_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_cfg_x = reg_pmp_6_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_cfg_w = reg_pmp_6_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_cfg_r = reg_pmp_6_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_addr = reg_pmp_6_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_6_mask = _T_341[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118512.4]
  assign io_pmp_7_cfg_l = reg_pmp_7_cfg_l; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_cfg_a = reg_pmp_7_cfg_a; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_cfg_x = reg_pmp_7_cfg_x; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_cfg_w = reg_pmp_7_cfg_w; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_cfg_r = reg_pmp_7_cfg_r; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_addr = reg_pmp_7_addr; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_pmp_7_mask = _T_350[31:0]; // @[CSR.scala 364:10:freechips.rocketchip.system.TinyConfig.fir@118513.4]
  assign io_trace_0_valid = _T_3810 | io_trace_0_exception; // @[CSR.scala 892:13:freechips.rocketchip.system.TinyConfig.fir@123143.4]
  assign io_trace_0_iaddr = io_pc; // @[CSR.scala 894:13:freechips.rocketchip.system.TinyConfig.fir@123145.4]
  assign io_trace_0_insn = io_inst_0; // @[CSR.scala 893:12:freechips.rocketchip.system.TinyConfig.fir@123144.4]
  assign io_trace_0_exception = _T_1130 | io_exception; // @[CSR.scala 891:17:freechips.rocketchip.system.TinyConfig.fir@123140.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_spp = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_dcsr_cause = _RAND_4[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_debug = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_dpc = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_dscratch = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_singleStepped = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_bp_0_control_dmode = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_bp_0_control_action = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_bp_0_control_tmatch = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_bp_0_control_x = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_bp_0_control_w = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_bp_0_control_r = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_bp_0_address = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  reg_pmp_0_cfg_l = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  reg_pmp_0_cfg_a = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  reg_pmp_0_cfg_x = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  reg_pmp_0_cfg_w = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  reg_pmp_0_cfg_r = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  reg_pmp_0_addr = _RAND_22[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  reg_pmp_1_cfg_l = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  reg_pmp_1_cfg_a = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  reg_pmp_1_cfg_x = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  reg_pmp_1_cfg_w = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  reg_pmp_1_cfg_r = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  reg_pmp_1_addr = _RAND_28[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  reg_pmp_2_cfg_l = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  reg_pmp_2_cfg_a = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  reg_pmp_2_cfg_x = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  reg_pmp_2_cfg_w = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  reg_pmp_2_cfg_r = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  reg_pmp_2_addr = _RAND_34[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  reg_pmp_3_cfg_l = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  reg_pmp_3_cfg_a = _RAND_36[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  reg_pmp_3_cfg_x = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  reg_pmp_3_cfg_w = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  reg_pmp_3_cfg_r = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  reg_pmp_3_addr = _RAND_40[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  reg_pmp_4_cfg_l = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  reg_pmp_4_cfg_a = _RAND_42[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  reg_pmp_4_cfg_x = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  reg_pmp_4_cfg_w = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  reg_pmp_4_cfg_r = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  reg_pmp_4_addr = _RAND_46[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  reg_pmp_5_cfg_l = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_pmp_5_cfg_a = _RAND_48[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  reg_pmp_5_cfg_x = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  reg_pmp_5_cfg_w = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  reg_pmp_5_cfg_r = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  reg_pmp_5_addr = _RAND_52[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  reg_pmp_6_cfg_l = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  reg_pmp_6_cfg_a = _RAND_54[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  reg_pmp_6_cfg_x = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  reg_pmp_6_cfg_w = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  reg_pmp_6_cfg_r = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  reg_pmp_6_addr = _RAND_58[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  reg_pmp_7_cfg_l = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  reg_pmp_7_cfg_a = _RAND_60[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  reg_pmp_7_cfg_x = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  reg_pmp_7_cfg_w = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  reg_pmp_7_cfg_r = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  reg_pmp_7_addr = _RAND_64[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  reg_mie = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  reg_mepc = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  reg_mcause = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  reg_mtval = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  reg_mscratch = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  reg_mtvec = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  reg_wfi = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_83 = _RAND_72[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {2{`RANDOM}};
  _T_85 = _RAND_73[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_91 = _RAND_74[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {2{`RANDOM}};
  _T_93 = _RAND_75[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  reg_misa = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1481 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_spp <= 1'h0;
    end else begin
      reg_mstatus_spp <= _GEN_85[0];
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_565) begin
          reg_mstatus_mpie <= _T_3342;
        end else begin
          if (insn_ret) begin
            if (_T_1468) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  reg_mstatus_mpie <= reg_mstatus_mie;
                end
              end
            end else begin
              reg_mstatus_mpie <= 1'h1;
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_1468) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mpie <= reg_mstatus_mie;
              end
            end
          end else begin
            reg_mstatus_mpie <= 1'h1;
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mpie <= reg_mstatus_mie;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_565) begin
          reg_mstatus_mie <= _T_3338;
        end else begin
          if (insn_ret) begin
            if (_T_1468) begin
              if (exception) begin
                if (!(trapToDebug)) begin
                  reg_mstatus_mie <= 1'h0;
                end
              end
            end else begin
              reg_mstatus_mie <= reg_mstatus_mpie;
            end
          end else begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end
        end
      end else begin
        if (insn_ret) begin
          if (_T_1468) begin
            if (exception) begin
              if (!(trapToDebug)) begin
                reg_mstatus_mie <= 1'h0;
              end
            end
          end else begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end else begin
          if (exception) begin
            if (!(trapToDebug)) begin
              reg_mstatus_mie <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_574) begin
          reg_dcsr_ebreakm <= _T_3453;
        end
      end
    end
    if (reset) begin
      reg_dcsr_cause <= 3'h0;
    end else begin
      if (exception) begin
        if (trapToDebug) begin
          if (_T_1062) begin
            if (reg_singleStepped) begin
              reg_dcsr_cause <= 3'h4;
            end else begin
              reg_dcsr_cause <= {{1'd0}, _T_1178};
            end
          end
        end
      end
    end
    if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_574) begin
          reg_dcsr_step <= _T_3369;
        end
      end
    end
    if (reset) begin
      reg_debug <= 1'h0;
    end else begin
      if (insn_ret) begin
        if (_T_1468) begin
          reg_debug <= 1'h0;
        end else begin
          if (exception) begin
            if (trapToDebug) begin
              if (_T_1062) begin
                reg_debug <= 1'h1;
              end
            end
          end
        end
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_1062) begin
              reg_debug <= 1'h1;
            end
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_575) begin
        reg_dpc <= _T_3424;
      end else begin
        if (exception) begin
          if (trapToDebug) begin
            if (_T_1062) begin
              reg_dpc <= epc;
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (trapToDebug) begin
          if (_T_1062) begin
            reg_dpc <= epc;
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_576) begin
        reg_dscratch <= wdata;
      end
    end
    if (_T_273) begin
      reg_singleStepped <= 1'h0;
    end else begin
      if (_T_1160) begin
        reg_singleStepped <= 1'h1;
      end
    end
    if (reset) begin
      reg_bp_0_control_dmode <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3462) begin
          if (_T_562) begin
            reg_bp_0_control_dmode <= _T_3520;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_action <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3462) begin
          if (_T_562) begin
            if (_T_3520) begin
              reg_bp_0_control_action <= _T_3515;
            end else begin
              reg_bp_0_control_action <= 1'h0;
            end
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_3462) begin
        if (_T_562) begin
          reg_bp_0_control_tmatch <= _T_3473;
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_x <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3462) begin
          if (_T_562) begin
            reg_bp_0_control_x <= _T_3369;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_w <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3462) begin
          if (_T_562) begin
            reg_bp_0_control_w <= _T_3467;
          end
        end
      end
    end
    if (reset) begin
      reg_bp_0_control_r <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3462) begin
          if (_T_562) begin
            reg_bp_0_control_r <= _T_3466;
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_3462) begin
        if (_T_563) begin
          reg_bp_0_address <= wdata;
        end
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3605) begin
          reg_pmp_0_cfg_l <= _T_3614;
        end
      end
    end
    if (reset) begin
      reg_pmp_0_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3605) begin
          reg_pmp_0_cfg_a <= _T_3612;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3605) begin
        reg_pmp_0_cfg_x <= _T_3611;
      end
    end
    if (csr_wen) begin
      if (_T_3605) begin
        reg_pmp_0_cfg_w <= _T_3615;
      end
    end
    if (csr_wen) begin
      if (_T_3605) begin
        reg_pmp_0_cfg_r <= _T_3609;
      end
    end
    reg_pmp_0_addr <= _GEN_329[29:0];
    if (reset) begin
      reg_pmp_1_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3625) begin
          reg_pmp_1_cfg_l <= _T_3634;
        end
      end
    end
    if (reset) begin
      reg_pmp_1_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3625) begin
          reg_pmp_1_cfg_a <= _T_3632;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3625) begin
        reg_pmp_1_cfg_x <= _T_3631;
      end
    end
    if (csr_wen) begin
      if (_T_3625) begin
        reg_pmp_1_cfg_w <= _T_3635;
      end
    end
    if (csr_wen) begin
      if (_T_3625) begin
        reg_pmp_1_cfg_r <= _T_3629;
      end
    end
    reg_pmp_1_addr <= _GEN_336[29:0];
    if (reset) begin
      reg_pmp_2_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3645) begin
          reg_pmp_2_cfg_l <= _T_3654;
        end
      end
    end
    if (reset) begin
      reg_pmp_2_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3645) begin
          reg_pmp_2_cfg_a <= _T_3652;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3645) begin
        reg_pmp_2_cfg_x <= _T_3651;
      end
    end
    if (csr_wen) begin
      if (_T_3645) begin
        reg_pmp_2_cfg_w <= _T_3655;
      end
    end
    if (csr_wen) begin
      if (_T_3645) begin
        reg_pmp_2_cfg_r <= _T_3649;
      end
    end
    reg_pmp_2_addr <= _GEN_343[29:0];
    if (reset) begin
      reg_pmp_3_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3665) begin
          reg_pmp_3_cfg_l <= _T_3674;
        end
      end
    end
    if (reset) begin
      reg_pmp_3_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3665) begin
          reg_pmp_3_cfg_a <= _T_3672;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3665) begin
        reg_pmp_3_cfg_x <= _T_3671;
      end
    end
    if (csr_wen) begin
      if (_T_3665) begin
        reg_pmp_3_cfg_w <= _T_3675;
      end
    end
    if (csr_wen) begin
      if (_T_3665) begin
        reg_pmp_3_cfg_r <= _T_3669;
      end
    end
    reg_pmp_3_addr <= _GEN_350[29:0];
    if (reset) begin
      reg_pmp_4_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3685) begin
          reg_pmp_4_cfg_l <= _T_3614;
        end
      end
    end
    if (reset) begin
      reg_pmp_4_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3685) begin
          reg_pmp_4_cfg_a <= _T_3612;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3685) begin
        reg_pmp_4_cfg_x <= _T_3611;
      end
    end
    if (csr_wen) begin
      if (_T_3685) begin
        reg_pmp_4_cfg_w <= _T_3615;
      end
    end
    if (csr_wen) begin
      if (_T_3685) begin
        reg_pmp_4_cfg_r <= _T_3609;
      end
    end
    reg_pmp_4_addr <= _GEN_357[29:0];
    if (reset) begin
      reg_pmp_5_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3705) begin
          reg_pmp_5_cfg_l <= _T_3634;
        end
      end
    end
    if (reset) begin
      reg_pmp_5_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3705) begin
          reg_pmp_5_cfg_a <= _T_3632;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3705) begin
        reg_pmp_5_cfg_x <= _T_3631;
      end
    end
    if (csr_wen) begin
      if (_T_3705) begin
        reg_pmp_5_cfg_w <= _T_3635;
      end
    end
    if (csr_wen) begin
      if (_T_3705) begin
        reg_pmp_5_cfg_r <= _T_3629;
      end
    end
    reg_pmp_5_addr <= _GEN_364[29:0];
    if (reset) begin
      reg_pmp_6_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3725) begin
          reg_pmp_6_cfg_l <= _T_3654;
        end
      end
    end
    if (reset) begin
      reg_pmp_6_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3725) begin
          reg_pmp_6_cfg_a <= _T_3652;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3725) begin
        reg_pmp_6_cfg_x <= _T_3651;
      end
    end
    if (csr_wen) begin
      if (_T_3725) begin
        reg_pmp_6_cfg_w <= _T_3655;
      end
    end
    if (csr_wen) begin
      if (_T_3725) begin
        reg_pmp_6_cfg_r <= _T_3649;
      end
    end
    reg_pmp_6_addr <= _GEN_371[29:0];
    if (reset) begin
      reg_pmp_7_cfg_l <= 1'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3745) begin
          reg_pmp_7_cfg_l <= _T_3674;
        end
      end
    end
    if (reset) begin
      reg_pmp_7_cfg_a <= 2'h0;
    end else begin
      if (csr_wen) begin
        if (_T_3745) begin
          reg_pmp_7_cfg_a <= _T_3672;
        end
      end
    end
    if (csr_wen) begin
      if (_T_3745) begin
        reg_pmp_7_cfg_x <= _T_3671;
      end
    end
    if (csr_wen) begin
      if (_T_3745) begin
        reg_pmp_7_cfg_w <= _T_3675;
      end
    end
    if (csr_wen) begin
      if (_T_3745) begin
        reg_pmp_7_cfg_r <= _T_3669;
      end
    end
    reg_pmp_7_addr <= _GEN_378[29:0];
    if (csr_wen) begin
      if (_T_568) begin
        reg_mie <= _T_3421;
      end
    end
    if (csr_wen) begin
      if (_T_570) begin
        reg_mepc <= _T_3424;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mepc <= epc;
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          reg_mepc <= epc;
        end
      end
    end
    if (csr_wen) begin
      if (_T_572) begin
        reg_mcause <= _T_3425;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            if (insn_call) begin
              reg_mcause <= 32'hb;
            end else begin
              if (insn_break) begin
                reg_mcause <= 32'h3;
              end else begin
                reg_mcause <= io_cause;
              end
            end
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          if (insn_call) begin
            reg_mcause <= 32'hb;
          end else begin
            if (insn_break) begin
              reg_mcause <= 32'h3;
            end else begin
              reg_mcause <= io_cause;
            end
          end
        end
      end
    end
    if (csr_wen) begin
      if (_T_571) begin
        reg_mtval <= wdata;
      end else begin
        if (exception) begin
          if (!(trapToDebug)) begin
            reg_mtval <= io_tval;
          end
        end
      end
    end else begin
      if (exception) begin
        if (!(trapToDebug)) begin
          reg_mtval <= io_tval;
        end
      end
    end
    if (csr_wen) begin
      if (_T_569) begin
        reg_mscratch <= wdata;
      end
    end
    if (reset) begin
      reg_mtvec <= 32'h0;
    end else begin
      if (csr_wen) begin
        if (_T_566) begin
          reg_mtvec <= wdata;
        end
      end
    end
    if (reset) begin
      _T_83 <= 6'h0;
    end else begin
      _T_83 <= _GEN_284[5:0];
    end
    if (reset) begin
      _T_85 <= 58'h0;
    end else begin
      if (csr_wen) begin
        if (_T_667) begin
          _T_85 <= _T_3440;
        end else begin
          if (_T_578) begin
            _T_85 <= _T_3436;
          end else begin
            if (_T_86) begin
              _T_85 <= _T_88;
            end
          end
        end
      end else begin
        if (_T_86) begin
          _T_85 <= _T_88;
        end
      end
    end
    if (reset) begin
      reg_misa <= 32'h40801105;
    end else begin
      if (csr_wen) begin
        if (_T_564) begin
          if (_T_3370) begin
            reg_misa <= _T_3379;
          end
        end
      end
    end
    if (reset) begin
      _T_1481 <= 1'h0;
    end else begin
      if (insn_cease) begin
        _T_1481 <= 1'h1;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1151) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:579 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119374.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1151) begin
          $fatal; // @[CSR.scala 579:9:freechips.rocketchip.system.TinyConfig.fir@119375.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1173) begin
          $fwrite(32'h80000002,"Assertion failed\n    at CSR.scala:587 assert(!reg_singleStepped || io.retire === UInt(0))\n"); // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119416.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_1173) begin
          $fatal; // @[CSR.scala 587:9:freechips.rocketchip.system.TinyConfig.fir@119417.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
  always @(posedge io_ungated_clock) begin
    if (reset) begin
      reg_wfi <= 1'h0;
    end else begin
      if (_T_1158) begin
        reg_wfi <= 1'h0;
      end else begin
        if (_T_1155) begin
          reg_wfi <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_91 <= 6'h0;
    end else begin
      _T_91 <= _GEN_282[5:0];
    end
    if (reset) begin
      _T_93 <= 58'h0;
    end else begin
      if (csr_wen) begin
        if (_T_666) begin
          _T_93 <= _T_3433;
        end else begin
          if (_T_577) begin
            _T_93 <= _T_3429;
          end else begin
            if (_T_94) begin
              _T_93 <= _T_96;
            end
          end
        end
      end else begin
        if (_T_94) begin
          _T_93 <= _T_96;
        end
      end
    end
  end
endmodule