module perf_counters
(
  clk_i,
  rst_ni,
  debug_mode_i,
  addr_i,
  we_i,
  data_i,
  data_o,
  commit_instr_i,
  commit_ack_i,
  l1_icache_miss_i,
  l1_dcache_miss_i,
  itlb_miss_i,
  dtlb_miss_i,
  sb_full_i,
  if_empty_i,
  ex_i,
  eret_i,
  resolved_branch_i
);

  input [4:0] addr_i;
  input [63:0] data_i;
  output [63:0] data_o;
  input [723:0] commit_instr_i;
  input [1:0] commit_ack_i;
  input [128:0] ex_i;
  input [133:0] resolved_branch_i;
  input clk_i;
  input rst_ni;
  input debug_mode_i;
  input we_i;
  input l1_icache_miss_i;
  input l1_dcache_miss_i;
  input itlb_miss_i;
  input dtlb_miss_i;
  input sb_full_i;
  input if_empty_i;
  input eret_i;
  wire [63:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,
  N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,
  N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,
  N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,
  N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,
  N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,
  N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,
  N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,
  N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,
  N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,
  N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,
  N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,
  N4118,N4119,N4120,N4121,N4122,N4123;
  wire [895:0] perf_counter_d;
  reg [895:0] perf_counter_q;

  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[895] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[895] <= perf_counter_d[895];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[894] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[894] <= perf_counter_d[894];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[893] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[893] <= perf_counter_d[893];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[892] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[892] <= perf_counter_d[892];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[891] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[891] <= perf_counter_d[891];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[890] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[890] <= perf_counter_d[890];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[889] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[889] <= perf_counter_d[889];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[888] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[888] <= perf_counter_d[888];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[887] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[887] <= perf_counter_d[887];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[886] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[886] <= perf_counter_d[886];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[885] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[885] <= perf_counter_d[885];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[884] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[884] <= perf_counter_d[884];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[883] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[883] <= perf_counter_d[883];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[882] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[882] <= perf_counter_d[882];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[881] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[881] <= perf_counter_d[881];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[880] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[880] <= perf_counter_d[880];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[879] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[879] <= perf_counter_d[879];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[878] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[878] <= perf_counter_d[878];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[877] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[877] <= perf_counter_d[877];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[876] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[876] <= perf_counter_d[876];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[875] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[875] <= perf_counter_d[875];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[874] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[874] <= perf_counter_d[874];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[873] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[873] <= perf_counter_d[873];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[872] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[872] <= perf_counter_d[872];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[871] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[871] <= perf_counter_d[871];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[870] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[870] <= perf_counter_d[870];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[869] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[869] <= perf_counter_d[869];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[868] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[868] <= perf_counter_d[868];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[867] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[867] <= perf_counter_d[867];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[866] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[866] <= perf_counter_d[866];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[865] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[865] <= perf_counter_d[865];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[864] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[864] <= perf_counter_d[864];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[863] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[863] <= perf_counter_d[863];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[862] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[862] <= perf_counter_d[862];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[861] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[861] <= perf_counter_d[861];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[860] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[860] <= perf_counter_d[860];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[859] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[859] <= perf_counter_d[859];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[858] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[858] <= perf_counter_d[858];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[857] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[857] <= perf_counter_d[857];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[856] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[856] <= perf_counter_d[856];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[855] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[855] <= perf_counter_d[855];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[854] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[854] <= perf_counter_d[854];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[853] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[853] <= perf_counter_d[853];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[852] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[852] <= perf_counter_d[852];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[851] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[851] <= perf_counter_d[851];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[850] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[850] <= perf_counter_d[850];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[849] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[849] <= perf_counter_d[849];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[848] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[848] <= perf_counter_d[848];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[847] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[847] <= perf_counter_d[847];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[846] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[846] <= perf_counter_d[846];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[845] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[845] <= perf_counter_d[845];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[844] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[844] <= perf_counter_d[844];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[843] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[843] <= perf_counter_d[843];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[842] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[842] <= perf_counter_d[842];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[841] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[841] <= perf_counter_d[841];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[840] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[840] <= perf_counter_d[840];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[839] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[839] <= perf_counter_d[839];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[838] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[838] <= perf_counter_d[838];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[837] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[837] <= perf_counter_d[837];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[836] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[836] <= perf_counter_d[836];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[835] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[835] <= perf_counter_d[835];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[834] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[834] <= perf_counter_d[834];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[833] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[833] <= perf_counter_d[833];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[832] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[832] <= perf_counter_d[832];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[831] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[831] <= perf_counter_d[831];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[830] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[830] <= perf_counter_d[830];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[829] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[829] <= perf_counter_d[829];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[828] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[828] <= perf_counter_d[828];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[827] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[827] <= perf_counter_d[827];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[826] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[826] <= perf_counter_d[826];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[825] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[825] <= perf_counter_d[825];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[824] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[824] <= perf_counter_d[824];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[823] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[823] <= perf_counter_d[823];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[822] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[822] <= perf_counter_d[822];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[821] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[821] <= perf_counter_d[821];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[820] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[820] <= perf_counter_d[820];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[819] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[819] <= perf_counter_d[819];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[818] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[818] <= perf_counter_d[818];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[817] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[817] <= perf_counter_d[817];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[816] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[816] <= perf_counter_d[816];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[815] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[815] <= perf_counter_d[815];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[814] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[814] <= perf_counter_d[814];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[813] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[813] <= perf_counter_d[813];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[812] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[812] <= perf_counter_d[812];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[811] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[811] <= perf_counter_d[811];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[810] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[810] <= perf_counter_d[810];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[809] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[809] <= perf_counter_d[809];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[808] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[808] <= perf_counter_d[808];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[807] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[807] <= perf_counter_d[807];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[806] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[806] <= perf_counter_d[806];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[805] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[805] <= perf_counter_d[805];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[804] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[804] <= perf_counter_d[804];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[803] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[803] <= perf_counter_d[803];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[802] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[802] <= perf_counter_d[802];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[801] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[801] <= perf_counter_d[801];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[800] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[800] <= perf_counter_d[800];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[799] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[799] <= perf_counter_d[799];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[798] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[798] <= perf_counter_d[798];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[797] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[797] <= perf_counter_d[797];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[796] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[796] <= perf_counter_d[796];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[795] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[795] <= perf_counter_d[795];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[794] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[794] <= perf_counter_d[794];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[793] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[793] <= perf_counter_d[793];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[792] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[792] <= perf_counter_d[792];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[791] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[791] <= perf_counter_d[791];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[790] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[790] <= perf_counter_d[790];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[789] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[789] <= perf_counter_d[789];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[788] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[788] <= perf_counter_d[788];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[787] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[787] <= perf_counter_d[787];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[786] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[786] <= perf_counter_d[786];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[785] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[785] <= perf_counter_d[785];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[784] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[784] <= perf_counter_d[784];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[783] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[783] <= perf_counter_d[783];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[782] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[782] <= perf_counter_d[782];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[781] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[781] <= perf_counter_d[781];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[780] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[780] <= perf_counter_d[780];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[779] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[779] <= perf_counter_d[779];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[778] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[778] <= perf_counter_d[778];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[777] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[777] <= perf_counter_d[777];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[776] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[776] <= perf_counter_d[776];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[775] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[775] <= perf_counter_d[775];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[774] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[774] <= perf_counter_d[774];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[773] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[773] <= perf_counter_d[773];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[772] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[772] <= perf_counter_d[772];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[771] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[771] <= perf_counter_d[771];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[770] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[770] <= perf_counter_d[770];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[769] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[769] <= perf_counter_d[769];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[768] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[768] <= perf_counter_d[768];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[767] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[767] <= perf_counter_d[767];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[766] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[766] <= perf_counter_d[766];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[765] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[765] <= perf_counter_d[765];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[764] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[764] <= perf_counter_d[764];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[763] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[763] <= perf_counter_d[763];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[762] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[762] <= perf_counter_d[762];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[761] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[761] <= perf_counter_d[761];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[760] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[760] <= perf_counter_d[760];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[759] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[759] <= perf_counter_d[759];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[758] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[758] <= perf_counter_d[758];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[757] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[757] <= perf_counter_d[757];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[756] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[756] <= perf_counter_d[756];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[755] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[755] <= perf_counter_d[755];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[754] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[754] <= perf_counter_d[754];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[753] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[753] <= perf_counter_d[753];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[752] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[752] <= perf_counter_d[752];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[751] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[751] <= perf_counter_d[751];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[750] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[750] <= perf_counter_d[750];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[749] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[749] <= perf_counter_d[749];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[748] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[748] <= perf_counter_d[748];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[747] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[747] <= perf_counter_d[747];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[746] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[746] <= perf_counter_d[746];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[745] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[745] <= perf_counter_d[745];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[744] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[744] <= perf_counter_d[744];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[743] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[743] <= perf_counter_d[743];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[742] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[742] <= perf_counter_d[742];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[741] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[741] <= perf_counter_d[741];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[740] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[740] <= perf_counter_d[740];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[739] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[739] <= perf_counter_d[739];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[738] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[738] <= perf_counter_d[738];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[737] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[737] <= perf_counter_d[737];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[736] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[736] <= perf_counter_d[736];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[735] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[735] <= perf_counter_d[735];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[734] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[734] <= perf_counter_d[734];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[733] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[733] <= perf_counter_d[733];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[732] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[732] <= perf_counter_d[732];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[731] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[731] <= perf_counter_d[731];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[730] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[730] <= perf_counter_d[730];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[729] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[729] <= perf_counter_d[729];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[728] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[728] <= perf_counter_d[728];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[727] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[727] <= perf_counter_d[727];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[726] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[726] <= perf_counter_d[726];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[725] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[725] <= perf_counter_d[725];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[724] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[724] <= perf_counter_d[724];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[723] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[723] <= perf_counter_d[723];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[722] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[722] <= perf_counter_d[722];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[721] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[721] <= perf_counter_d[721];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[720] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[720] <= perf_counter_d[720];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[719] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[719] <= perf_counter_d[719];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[718] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[718] <= perf_counter_d[718];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[717] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[717] <= perf_counter_d[717];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[716] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[716] <= perf_counter_d[716];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[715] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[715] <= perf_counter_d[715];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[714] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[714] <= perf_counter_d[714];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[713] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[713] <= perf_counter_d[713];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[712] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[712] <= perf_counter_d[712];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[711] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[711] <= perf_counter_d[711];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[710] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[710] <= perf_counter_d[710];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[709] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[709] <= perf_counter_d[709];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[708] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[708] <= perf_counter_d[708];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[707] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[707] <= perf_counter_d[707];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[706] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[706] <= perf_counter_d[706];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[705] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[705] <= perf_counter_d[705];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[704] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[704] <= perf_counter_d[704];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[703] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[703] <= perf_counter_d[703];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[702] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[702] <= perf_counter_d[702];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[701] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[701] <= perf_counter_d[701];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[700] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[700] <= perf_counter_d[700];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[699] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[699] <= perf_counter_d[699];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[698] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[698] <= perf_counter_d[698];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[697] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[697] <= perf_counter_d[697];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[696] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[696] <= perf_counter_d[696];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[695] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[695] <= perf_counter_d[695];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[694] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[694] <= perf_counter_d[694];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[693] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[693] <= perf_counter_d[693];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[692] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[692] <= perf_counter_d[692];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[691] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[691] <= perf_counter_d[691];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[690] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[690] <= perf_counter_d[690];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[689] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[689] <= perf_counter_d[689];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[688] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[688] <= perf_counter_d[688];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[687] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[687] <= perf_counter_d[687];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[686] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[686] <= perf_counter_d[686];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[685] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[685] <= perf_counter_d[685];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[684] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[684] <= perf_counter_d[684];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[683] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[683] <= perf_counter_d[683];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[682] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[682] <= perf_counter_d[682];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[681] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[681] <= perf_counter_d[681];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[680] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[680] <= perf_counter_d[680];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[679] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[679] <= perf_counter_d[679];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[678] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[678] <= perf_counter_d[678];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[677] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[677] <= perf_counter_d[677];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[676] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[676] <= perf_counter_d[676];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[675] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[675] <= perf_counter_d[675];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[674] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[674] <= perf_counter_d[674];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[673] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[673] <= perf_counter_d[673];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[672] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[672] <= perf_counter_d[672];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[671] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[671] <= perf_counter_d[671];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[670] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[670] <= perf_counter_d[670];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[669] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[669] <= perf_counter_d[669];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[668] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[668] <= perf_counter_d[668];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[667] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[667] <= perf_counter_d[667];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[666] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[666] <= perf_counter_d[666];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[665] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[665] <= perf_counter_d[665];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[664] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[664] <= perf_counter_d[664];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[663] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[663] <= perf_counter_d[663];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[662] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[662] <= perf_counter_d[662];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[661] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[661] <= perf_counter_d[661];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[660] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[660] <= perf_counter_d[660];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[659] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[659] <= perf_counter_d[659];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[658] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[658] <= perf_counter_d[658];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[657] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[657] <= perf_counter_d[657];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[656] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[656] <= perf_counter_d[656];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[655] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[655] <= perf_counter_d[655];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[654] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[654] <= perf_counter_d[654];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[653] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[653] <= perf_counter_d[653];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[652] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[652] <= perf_counter_d[652];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[651] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[651] <= perf_counter_d[651];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[650] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[650] <= perf_counter_d[650];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[649] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[649] <= perf_counter_d[649];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[648] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[648] <= perf_counter_d[648];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[647] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[647] <= perf_counter_d[647];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[646] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[646] <= perf_counter_d[646];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[645] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[645] <= perf_counter_d[645];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[644] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[644] <= perf_counter_d[644];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[643] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[643] <= perf_counter_d[643];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[642] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[642] <= perf_counter_d[642];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[641] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[641] <= perf_counter_d[641];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[640] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[640] <= perf_counter_d[640];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[639] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[639] <= perf_counter_d[639];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[638] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[638] <= perf_counter_d[638];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[637] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[637] <= perf_counter_d[637];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[636] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[636] <= perf_counter_d[636];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[635] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[635] <= perf_counter_d[635];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[634] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[634] <= perf_counter_d[634];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[633] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[633] <= perf_counter_d[633];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[632] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[632] <= perf_counter_d[632];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[631] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[631] <= perf_counter_d[631];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[630] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[630] <= perf_counter_d[630];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[629] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[629] <= perf_counter_d[629];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[628] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[628] <= perf_counter_d[628];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[627] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[627] <= perf_counter_d[627];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[626] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[626] <= perf_counter_d[626];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[625] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[625] <= perf_counter_d[625];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[624] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[624] <= perf_counter_d[624];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[623] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[623] <= perf_counter_d[623];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[622] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[622] <= perf_counter_d[622];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[621] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[621] <= perf_counter_d[621];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[620] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[620] <= perf_counter_d[620];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[619] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[619] <= perf_counter_d[619];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[618] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[618] <= perf_counter_d[618];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[617] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[617] <= perf_counter_d[617];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[616] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[616] <= perf_counter_d[616];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[615] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[615] <= perf_counter_d[615];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[614] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[614] <= perf_counter_d[614];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[613] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[613] <= perf_counter_d[613];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[612] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[612] <= perf_counter_d[612];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[611] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[611] <= perf_counter_d[611];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[610] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[610] <= perf_counter_d[610];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[609] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[609] <= perf_counter_d[609];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[608] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[608] <= perf_counter_d[608];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[607] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[607] <= perf_counter_d[607];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[606] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[606] <= perf_counter_d[606];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[605] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[605] <= perf_counter_d[605];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[604] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[604] <= perf_counter_d[604];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[603] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[603] <= perf_counter_d[603];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[602] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[602] <= perf_counter_d[602];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[601] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[601] <= perf_counter_d[601];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[600] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[600] <= perf_counter_d[600];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[599] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[599] <= perf_counter_d[599];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[598] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[598] <= perf_counter_d[598];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[597] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[597] <= perf_counter_d[597];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[596] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[596] <= perf_counter_d[596];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[595] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[595] <= perf_counter_d[595];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[594] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[594] <= perf_counter_d[594];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[593] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[593] <= perf_counter_d[593];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[592] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[592] <= perf_counter_d[592];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[591] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[591] <= perf_counter_d[591];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[590] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[590] <= perf_counter_d[590];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[589] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[589] <= perf_counter_d[589];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[588] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[588] <= perf_counter_d[588];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[587] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[587] <= perf_counter_d[587];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[586] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[586] <= perf_counter_d[586];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[585] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[585] <= perf_counter_d[585];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[584] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[584] <= perf_counter_d[584];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[583] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[583] <= perf_counter_d[583];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[582] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[582] <= perf_counter_d[582];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[581] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[581] <= perf_counter_d[581];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[580] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[580] <= perf_counter_d[580];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[579] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[579] <= perf_counter_d[579];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[578] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[578] <= perf_counter_d[578];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[577] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[577] <= perf_counter_d[577];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[576] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[576] <= perf_counter_d[576];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[575] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[575] <= perf_counter_d[575];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[574] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[574] <= perf_counter_d[574];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[573] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[573] <= perf_counter_d[573];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[572] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[572] <= perf_counter_d[572];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[571] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[571] <= perf_counter_d[571];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[570] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[570] <= perf_counter_d[570];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[569] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[569] <= perf_counter_d[569];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[568] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[568] <= perf_counter_d[568];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[567] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[567] <= perf_counter_d[567];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[566] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[566] <= perf_counter_d[566];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[565] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[565] <= perf_counter_d[565];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[564] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[564] <= perf_counter_d[564];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[563] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[563] <= perf_counter_d[563];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[562] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[562] <= perf_counter_d[562];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[561] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[561] <= perf_counter_d[561];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[560] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[560] <= perf_counter_d[560];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[559] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[559] <= perf_counter_d[559];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[558] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[558] <= perf_counter_d[558];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[557] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[557] <= perf_counter_d[557];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[556] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[556] <= perf_counter_d[556];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[555] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[555] <= perf_counter_d[555];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[554] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[554] <= perf_counter_d[554];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[553] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[553] <= perf_counter_d[553];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[552] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[552] <= perf_counter_d[552];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[551] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[551] <= perf_counter_d[551];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[550] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[550] <= perf_counter_d[550];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[549] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[549] <= perf_counter_d[549];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[548] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[548] <= perf_counter_d[548];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[547] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[547] <= perf_counter_d[547];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[546] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[546] <= perf_counter_d[546];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[545] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[545] <= perf_counter_d[545];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[544] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[544] <= perf_counter_d[544];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[543] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[543] <= perf_counter_d[543];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[542] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[542] <= perf_counter_d[542];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[541] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[541] <= perf_counter_d[541];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[540] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[540] <= perf_counter_d[540];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[539] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[539] <= perf_counter_d[539];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[538] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[538] <= perf_counter_d[538];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[537] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[537] <= perf_counter_d[537];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[536] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[536] <= perf_counter_d[536];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[535] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[535] <= perf_counter_d[535];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[534] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[534] <= perf_counter_d[534];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[533] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[533] <= perf_counter_d[533];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[532] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[532] <= perf_counter_d[532];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[531] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[531] <= perf_counter_d[531];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[530] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[530] <= perf_counter_d[530];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[529] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[529] <= perf_counter_d[529];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[528] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[528] <= perf_counter_d[528];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[527] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[527] <= perf_counter_d[527];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[526] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[526] <= perf_counter_d[526];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[525] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[525] <= perf_counter_d[525];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[524] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[524] <= perf_counter_d[524];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[523] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[523] <= perf_counter_d[523];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[522] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[522] <= perf_counter_d[522];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[521] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[521] <= perf_counter_d[521];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[520] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[520] <= perf_counter_d[520];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[519] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[519] <= perf_counter_d[519];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[518] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[518] <= perf_counter_d[518];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[517] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[517] <= perf_counter_d[517];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[516] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[516] <= perf_counter_d[516];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[515] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[515] <= perf_counter_d[515];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[514] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[514] <= perf_counter_d[514];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[513] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[513] <= perf_counter_d[513];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[512] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[512] <= perf_counter_d[512];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[511] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[511] <= perf_counter_d[511];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[510] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[510] <= perf_counter_d[510];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[509] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[509] <= perf_counter_d[509];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[508] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[508] <= perf_counter_d[508];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[507] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[507] <= perf_counter_d[507];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[506] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[506] <= perf_counter_d[506];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[505] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[505] <= perf_counter_d[505];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[504] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[504] <= perf_counter_d[504];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[503] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[503] <= perf_counter_d[503];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[502] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[502] <= perf_counter_d[502];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[501] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[501] <= perf_counter_d[501];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[500] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[500] <= perf_counter_d[500];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[499] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[499] <= perf_counter_d[499];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[498] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[498] <= perf_counter_d[498];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[497] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[497] <= perf_counter_d[497];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[496] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[496] <= perf_counter_d[496];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[495] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[495] <= perf_counter_d[495];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[494] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[494] <= perf_counter_d[494];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[493] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[493] <= perf_counter_d[493];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[492] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[492] <= perf_counter_d[492];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[491] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[491] <= perf_counter_d[491];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[490] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[490] <= perf_counter_d[490];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[489] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[489] <= perf_counter_d[489];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[488] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[488] <= perf_counter_d[488];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[487] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[487] <= perf_counter_d[487];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[486] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[486] <= perf_counter_d[486];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[485] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[485] <= perf_counter_d[485];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[484] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[484] <= perf_counter_d[484];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[483] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[483] <= perf_counter_d[483];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[482] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[482] <= perf_counter_d[482];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[481] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[481] <= perf_counter_d[481];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[480] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[480] <= perf_counter_d[480];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[479] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[479] <= perf_counter_d[479];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[478] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[478] <= perf_counter_d[478];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[477] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[477] <= perf_counter_d[477];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[476] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[476] <= perf_counter_d[476];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[475] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[475] <= perf_counter_d[475];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[474] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[474] <= perf_counter_d[474];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[473] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[473] <= perf_counter_d[473];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[472] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[472] <= perf_counter_d[472];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[471] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[471] <= perf_counter_d[471];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[470] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[470] <= perf_counter_d[470];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[469] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[469] <= perf_counter_d[469];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[468] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[468] <= perf_counter_d[468];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[467] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[467] <= perf_counter_d[467];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[466] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[466] <= perf_counter_d[466];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[465] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[465] <= perf_counter_d[465];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[464] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[464] <= perf_counter_d[464];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[463] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[463] <= perf_counter_d[463];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[462] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[462] <= perf_counter_d[462];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[461] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[461] <= perf_counter_d[461];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[460] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[460] <= perf_counter_d[460];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[459] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[459] <= perf_counter_d[459];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[458] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[458] <= perf_counter_d[458];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[457] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[457] <= perf_counter_d[457];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[456] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[456] <= perf_counter_d[456];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[455] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[455] <= perf_counter_d[455];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[454] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[454] <= perf_counter_d[454];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[453] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[453] <= perf_counter_d[453];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[452] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[452] <= perf_counter_d[452];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[451] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[451] <= perf_counter_d[451];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[450] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[450] <= perf_counter_d[450];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[449] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[449] <= perf_counter_d[449];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[448] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[448] <= perf_counter_d[448];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[447] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[447] <= perf_counter_d[447];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[446] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[446] <= perf_counter_d[446];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[445] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[445] <= perf_counter_d[445];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[444] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[444] <= perf_counter_d[444];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[443] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[443] <= perf_counter_d[443];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[442] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[442] <= perf_counter_d[442];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[441] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[441] <= perf_counter_d[441];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[440] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[440] <= perf_counter_d[440];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[439] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[439] <= perf_counter_d[439];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[438] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[438] <= perf_counter_d[438];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[437] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[437] <= perf_counter_d[437];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[436] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[436] <= perf_counter_d[436];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[435] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[435] <= perf_counter_d[435];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[434] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[434] <= perf_counter_d[434];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[433] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[433] <= perf_counter_d[433];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[432] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[432] <= perf_counter_d[432];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[431] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[431] <= perf_counter_d[431];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[430] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[430] <= perf_counter_d[430];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[429] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[429] <= perf_counter_d[429];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[428] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[428] <= perf_counter_d[428];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[427] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[427] <= perf_counter_d[427];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[426] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[426] <= perf_counter_d[426];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[425] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[425] <= perf_counter_d[425];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[424] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[424] <= perf_counter_d[424];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[423] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[423] <= perf_counter_d[423];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[422] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[422] <= perf_counter_d[422];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[421] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[421] <= perf_counter_d[421];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[420] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[420] <= perf_counter_d[420];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[419] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[419] <= perf_counter_d[419];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[418] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[418] <= perf_counter_d[418];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[417] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[417] <= perf_counter_d[417];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[416] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[416] <= perf_counter_d[416];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[415] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[415] <= perf_counter_d[415];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[414] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[414] <= perf_counter_d[414];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[413] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[413] <= perf_counter_d[413];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[412] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[412] <= perf_counter_d[412];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[411] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[411] <= perf_counter_d[411];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[410] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[410] <= perf_counter_d[410];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[409] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[409] <= perf_counter_d[409];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[408] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[408] <= perf_counter_d[408];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[407] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[407] <= perf_counter_d[407];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[406] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[406] <= perf_counter_d[406];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[405] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[405] <= perf_counter_d[405];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[404] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[404] <= perf_counter_d[404];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[403] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[403] <= perf_counter_d[403];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[402] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[402] <= perf_counter_d[402];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[401] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[401] <= perf_counter_d[401];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[400] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[400] <= perf_counter_d[400];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[399] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[399] <= perf_counter_d[399];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[398] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[398] <= perf_counter_d[398];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[397] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[397] <= perf_counter_d[397];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[396] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[396] <= perf_counter_d[396];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[395] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[395] <= perf_counter_d[395];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[394] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[394] <= perf_counter_d[394];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[393] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[393] <= perf_counter_d[393];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[392] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[392] <= perf_counter_d[392];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[391] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[391] <= perf_counter_d[391];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[390] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[390] <= perf_counter_d[390];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[389] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[389] <= perf_counter_d[389];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[388] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[388] <= perf_counter_d[388];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[387] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[387] <= perf_counter_d[387];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[386] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[386] <= perf_counter_d[386];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[385] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[385] <= perf_counter_d[385];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[384] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[384] <= perf_counter_d[384];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[383] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[383] <= perf_counter_d[383];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[382] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[382] <= perf_counter_d[382];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[381] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[381] <= perf_counter_d[381];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[380] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[380] <= perf_counter_d[380];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[379] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[379] <= perf_counter_d[379];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[378] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[378] <= perf_counter_d[378];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[377] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[377] <= perf_counter_d[377];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[376] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[376] <= perf_counter_d[376];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[375] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[375] <= perf_counter_d[375];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[374] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[374] <= perf_counter_d[374];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[373] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[373] <= perf_counter_d[373];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[372] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[372] <= perf_counter_d[372];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[371] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[371] <= perf_counter_d[371];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[370] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[370] <= perf_counter_d[370];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[369] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[369] <= perf_counter_d[369];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[368] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[368] <= perf_counter_d[368];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[367] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[367] <= perf_counter_d[367];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[366] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[366] <= perf_counter_d[366];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[365] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[365] <= perf_counter_d[365];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[364] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[364] <= perf_counter_d[364];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[363] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[363] <= perf_counter_d[363];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[362] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[362] <= perf_counter_d[362];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[361] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[361] <= perf_counter_d[361];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[360] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[360] <= perf_counter_d[360];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[359] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[359] <= perf_counter_d[359];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[358] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[358] <= perf_counter_d[358];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[357] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[357] <= perf_counter_d[357];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[356] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[356] <= perf_counter_d[356];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[355] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[355] <= perf_counter_d[355];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[354] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[354] <= perf_counter_d[354];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[353] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[353] <= perf_counter_d[353];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[352] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[352] <= perf_counter_d[352];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[351] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[351] <= perf_counter_d[351];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[350] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[350] <= perf_counter_d[350];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[349] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[349] <= perf_counter_d[349];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[348] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[348] <= perf_counter_d[348];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[347] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[347] <= perf_counter_d[347];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[346] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[346] <= perf_counter_d[346];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[345] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[345] <= perf_counter_d[345];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[344] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[344] <= perf_counter_d[344];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[343] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[343] <= perf_counter_d[343];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[342] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[342] <= perf_counter_d[342];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[341] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[341] <= perf_counter_d[341];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[340] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[340] <= perf_counter_d[340];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[339] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[339] <= perf_counter_d[339];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[338] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[338] <= perf_counter_d[338];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[337] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[337] <= perf_counter_d[337];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[336] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[336] <= perf_counter_d[336];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[335] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[335] <= perf_counter_d[335];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[334] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[334] <= perf_counter_d[334];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[333] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[333] <= perf_counter_d[333];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[332] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[332] <= perf_counter_d[332];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[331] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[331] <= perf_counter_d[331];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[330] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[330] <= perf_counter_d[330];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[329] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[329] <= perf_counter_d[329];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[328] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[328] <= perf_counter_d[328];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[327] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[327] <= perf_counter_d[327];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[326] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[326] <= perf_counter_d[326];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[325] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[325] <= perf_counter_d[325];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[324] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[324] <= perf_counter_d[324];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[323] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[323] <= perf_counter_d[323];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[322] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[322] <= perf_counter_d[322];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[321] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[321] <= perf_counter_d[321];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[320] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[320] <= perf_counter_d[320];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[319] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[319] <= perf_counter_d[319];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[318] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[318] <= perf_counter_d[318];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[317] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[317] <= perf_counter_d[317];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[316] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[316] <= perf_counter_d[316];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[315] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[315] <= perf_counter_d[315];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[314] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[314] <= perf_counter_d[314];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[313] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[313] <= perf_counter_d[313];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[312] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[312] <= perf_counter_d[312];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[311] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[311] <= perf_counter_d[311];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[310] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[310] <= perf_counter_d[310];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[309] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[309] <= perf_counter_d[309];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[308] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[308] <= perf_counter_d[308];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[307] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[307] <= perf_counter_d[307];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[306] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[306] <= perf_counter_d[306];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[305] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[305] <= perf_counter_d[305];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[304] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[304] <= perf_counter_d[304];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[303] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[303] <= perf_counter_d[303];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[302] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[302] <= perf_counter_d[302];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[301] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[301] <= perf_counter_d[301];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[300] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[300] <= perf_counter_d[300];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[299] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[299] <= perf_counter_d[299];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[298] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[298] <= perf_counter_d[298];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[297] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[297] <= perf_counter_d[297];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[296] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[296] <= perf_counter_d[296];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[295] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[295] <= perf_counter_d[295];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[294] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[294] <= perf_counter_d[294];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[293] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[293] <= perf_counter_d[293];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[292] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[292] <= perf_counter_d[292];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[291] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[291] <= perf_counter_d[291];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[290] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[290] <= perf_counter_d[290];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[289] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[289] <= perf_counter_d[289];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[288] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[288] <= perf_counter_d[288];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[287] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[287] <= perf_counter_d[287];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[286] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[286] <= perf_counter_d[286];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[285] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[285] <= perf_counter_d[285];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[284] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[284] <= perf_counter_d[284];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[283] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[283] <= perf_counter_d[283];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[282] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[282] <= perf_counter_d[282];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[281] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[281] <= perf_counter_d[281];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[280] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[280] <= perf_counter_d[280];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[279] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[279] <= perf_counter_d[279];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[278] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[278] <= perf_counter_d[278];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[277] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[277] <= perf_counter_d[277];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[276] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[276] <= perf_counter_d[276];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[275] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[275] <= perf_counter_d[275];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[274] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[274] <= perf_counter_d[274];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[273] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[273] <= perf_counter_d[273];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[272] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[272] <= perf_counter_d[272];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[271] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[271] <= perf_counter_d[271];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[270] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[270] <= perf_counter_d[270];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[269] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[269] <= perf_counter_d[269];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[268] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[268] <= perf_counter_d[268];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[267] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[267] <= perf_counter_d[267];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[266] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[266] <= perf_counter_d[266];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[265] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[265] <= perf_counter_d[265];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[264] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[264] <= perf_counter_d[264];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[263] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[263] <= perf_counter_d[263];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[262] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[262] <= perf_counter_d[262];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[261] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[261] <= perf_counter_d[261];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[260] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[260] <= perf_counter_d[260];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[259] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[259] <= perf_counter_d[259];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[258] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[258] <= perf_counter_d[258];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[257] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[257] <= perf_counter_d[257];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[256] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[256] <= perf_counter_d[256];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[255] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[255] <= perf_counter_d[255];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[254] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[254] <= perf_counter_d[254];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[253] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[253] <= perf_counter_d[253];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[252] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[252] <= perf_counter_d[252];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[251] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[251] <= perf_counter_d[251];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[250] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[250] <= perf_counter_d[250];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[249] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[249] <= perf_counter_d[249];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[248] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[248] <= perf_counter_d[248];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[247] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[247] <= perf_counter_d[247];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[246] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[246] <= perf_counter_d[246];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[245] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[245] <= perf_counter_d[245];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[244] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[244] <= perf_counter_d[244];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[243] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[243] <= perf_counter_d[243];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[242] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[242] <= perf_counter_d[242];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[241] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[241] <= perf_counter_d[241];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[240] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[240] <= perf_counter_d[240];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[239] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[239] <= perf_counter_d[239];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[238] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[238] <= perf_counter_d[238];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[237] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[237] <= perf_counter_d[237];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[236] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[236] <= perf_counter_d[236];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[235] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[235] <= perf_counter_d[235];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[234] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[234] <= perf_counter_d[234];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[233] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[233] <= perf_counter_d[233];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[232] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[232] <= perf_counter_d[232];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[231] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[231] <= perf_counter_d[231];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[230] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[230] <= perf_counter_d[230];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[229] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[229] <= perf_counter_d[229];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[228] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[228] <= perf_counter_d[228];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[227] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[227] <= perf_counter_d[227];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[226] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[226] <= perf_counter_d[226];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[225] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[225] <= perf_counter_d[225];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[224] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[224] <= perf_counter_d[224];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[223] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[223] <= perf_counter_d[223];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[222] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[222] <= perf_counter_d[222];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[221] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[221] <= perf_counter_d[221];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[220] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[220] <= perf_counter_d[220];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[219] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[219] <= perf_counter_d[219];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[218] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[218] <= perf_counter_d[218];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[217] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[217] <= perf_counter_d[217];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[216] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[216] <= perf_counter_d[216];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[215] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[215] <= perf_counter_d[215];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[214] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[214] <= perf_counter_d[214];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[213] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[213] <= perf_counter_d[213];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[212] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[212] <= perf_counter_d[212];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[211] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[211] <= perf_counter_d[211];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[210] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[210] <= perf_counter_d[210];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[209] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[209] <= perf_counter_d[209];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[208] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[208] <= perf_counter_d[208];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[207] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[207] <= perf_counter_d[207];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[206] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[206] <= perf_counter_d[206];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[205] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[205] <= perf_counter_d[205];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[204] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[204] <= perf_counter_d[204];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[203] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[203] <= perf_counter_d[203];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[202] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[202] <= perf_counter_d[202];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[201] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[201] <= perf_counter_d[201];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[200] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[200] <= perf_counter_d[200];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[199] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[199] <= perf_counter_d[199];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[198] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[198] <= perf_counter_d[198];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[197] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[197] <= perf_counter_d[197];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[196] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[196] <= perf_counter_d[196];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[195] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[195] <= perf_counter_d[195];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[194] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[194] <= perf_counter_d[194];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[193] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[193] <= perf_counter_d[193];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[192] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[192] <= perf_counter_d[192];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[191] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[191] <= perf_counter_d[191];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[190] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[190] <= perf_counter_d[190];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[189] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[189] <= perf_counter_d[189];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[188] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[188] <= perf_counter_d[188];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[187] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[187] <= perf_counter_d[187];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[186] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[186] <= perf_counter_d[186];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[185] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[185] <= perf_counter_d[185];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[184] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[184] <= perf_counter_d[184];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[183] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[183] <= perf_counter_d[183];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[182] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[182] <= perf_counter_d[182];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[181] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[181] <= perf_counter_d[181];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[180] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[180] <= perf_counter_d[180];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[179] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[179] <= perf_counter_d[179];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[178] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[178] <= perf_counter_d[178];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[177] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[177] <= perf_counter_d[177];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[176] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[176] <= perf_counter_d[176];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[175] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[175] <= perf_counter_d[175];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[174] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[174] <= perf_counter_d[174];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[173] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[173] <= perf_counter_d[173];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[172] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[172] <= perf_counter_d[172];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[171] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[171] <= perf_counter_d[171];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[170] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[170] <= perf_counter_d[170];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[169] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[169] <= perf_counter_d[169];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[168] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[168] <= perf_counter_d[168];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[167] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[167] <= perf_counter_d[167];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[166] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[166] <= perf_counter_d[166];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[165] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[165] <= perf_counter_d[165];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[164] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[164] <= perf_counter_d[164];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[163] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[163] <= perf_counter_d[163];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[162] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[162] <= perf_counter_d[162];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[161] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[161] <= perf_counter_d[161];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[160] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[160] <= perf_counter_d[160];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[159] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[159] <= perf_counter_d[159];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[158] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[158] <= perf_counter_d[158];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[157] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[157] <= perf_counter_d[157];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[156] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[156] <= perf_counter_d[156];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[155] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[155] <= perf_counter_d[155];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[154] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[154] <= perf_counter_d[154];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[153] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[153] <= perf_counter_d[153];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[152] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[152] <= perf_counter_d[152];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[151] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[151] <= perf_counter_d[151];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[150] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[150] <= perf_counter_d[150];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[149] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[149] <= perf_counter_d[149];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[148] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[148] <= perf_counter_d[148];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[147] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[147] <= perf_counter_d[147];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[146] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[146] <= perf_counter_d[146];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[145] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[145] <= perf_counter_d[145];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[144] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[144] <= perf_counter_d[144];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[143] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[143] <= perf_counter_d[143];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[142] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[142] <= perf_counter_d[142];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[141] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[141] <= perf_counter_d[141];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[140] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[140] <= perf_counter_d[140];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[139] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[139] <= perf_counter_d[139];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[138] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[138] <= perf_counter_d[138];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[137] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[137] <= perf_counter_d[137];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[136] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[136] <= perf_counter_d[136];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[135] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[135] <= perf_counter_d[135];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[134] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[134] <= perf_counter_d[134];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[133] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[133] <= perf_counter_d[133];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[132] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[132] <= perf_counter_d[132];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[131] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[131] <= perf_counter_d[131];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[130] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[130] <= perf_counter_d[130];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[129] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[129] <= perf_counter_d[129];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[128] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[128] <= perf_counter_d[128];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[127] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[127] <= perf_counter_d[127];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[126] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[126] <= perf_counter_d[126];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[125] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[125] <= perf_counter_d[125];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[124] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[124] <= perf_counter_d[124];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[123] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[123] <= perf_counter_d[123];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[122] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[122] <= perf_counter_d[122];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[121] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[121] <= perf_counter_d[121];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[120] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[120] <= perf_counter_d[120];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[119] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[119] <= perf_counter_d[119];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[118] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[118] <= perf_counter_d[118];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[117] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[117] <= perf_counter_d[117];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[116] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[116] <= perf_counter_d[116];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[115] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[115] <= perf_counter_d[115];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[114] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[114] <= perf_counter_d[114];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[113] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[113] <= perf_counter_d[113];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[112] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[112] <= perf_counter_d[112];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[111] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[111] <= perf_counter_d[111];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[110] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[110] <= perf_counter_d[110];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[109] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[109] <= perf_counter_d[109];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[108] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[108] <= perf_counter_d[108];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[107] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[107] <= perf_counter_d[107];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[106] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[106] <= perf_counter_d[106];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[105] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[105] <= perf_counter_d[105];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[104] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[104] <= perf_counter_d[104];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[103] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[103] <= perf_counter_d[103];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[102] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[102] <= perf_counter_d[102];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[101] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[101] <= perf_counter_d[101];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[100] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[100] <= perf_counter_d[100];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[99] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[99] <= perf_counter_d[99];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[98] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[98] <= perf_counter_d[98];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[97] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[97] <= perf_counter_d[97];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[96] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[96] <= perf_counter_d[96];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[95] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[95] <= perf_counter_d[95];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[94] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[94] <= perf_counter_d[94];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[93] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[93] <= perf_counter_d[93];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[92] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[92] <= perf_counter_d[92];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[91] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[91] <= perf_counter_d[91];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[90] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[90] <= perf_counter_d[90];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[89] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[89] <= perf_counter_d[89];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[88] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[88] <= perf_counter_d[88];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[87] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[87] <= perf_counter_d[87];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[86] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[86] <= perf_counter_d[86];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[85] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[85] <= perf_counter_d[85];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[84] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[84] <= perf_counter_d[84];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[83] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[83] <= perf_counter_d[83];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[82] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[82] <= perf_counter_d[82];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[81] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[81] <= perf_counter_d[81];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[80] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[80] <= perf_counter_d[80];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[79] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[79] <= perf_counter_d[79];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[78] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[78] <= perf_counter_d[78];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[77] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[77] <= perf_counter_d[77];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[76] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[76] <= perf_counter_d[76];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[75] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[75] <= perf_counter_d[75];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[74] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[74] <= perf_counter_d[74];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[73] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[73] <= perf_counter_d[73];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[72] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[72] <= perf_counter_d[72];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[71] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[71] <= perf_counter_d[71];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[70] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[70] <= perf_counter_d[70];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[69] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[69] <= perf_counter_d[69];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[68] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[68] <= perf_counter_d[68];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[67] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[67] <= perf_counter_d[67];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[66] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[66] <= perf_counter_d[66];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[65] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[65] <= perf_counter_d[65];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[64] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[64] <= perf_counter_d[64];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[63] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[63] <= perf_counter_d[63];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[62] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[62] <= perf_counter_d[62];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[61] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[61] <= perf_counter_d[61];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[60] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[60] <= perf_counter_d[60];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[59] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[59] <= perf_counter_d[59];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[58] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[58] <= perf_counter_d[58];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[57] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[57] <= perf_counter_d[57];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[56] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[56] <= perf_counter_d[56];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[55] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[55] <= perf_counter_d[55];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[54] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[54] <= perf_counter_d[54];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[53] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[53] <= perf_counter_d[53];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[52] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[52] <= perf_counter_d[52];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[51] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[51] <= perf_counter_d[51];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[50] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[50] <= perf_counter_d[50];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[49] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[49] <= perf_counter_d[49];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[48] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[48] <= perf_counter_d[48];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[47] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[47] <= perf_counter_d[47];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[46] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[46] <= perf_counter_d[46];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[45] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[45] <= perf_counter_d[45];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[44] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[44] <= perf_counter_d[44];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[43] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[43] <= perf_counter_d[43];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[42] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[42] <= perf_counter_d[42];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[41] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[41] <= perf_counter_d[41];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[40] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[40] <= perf_counter_d[40];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[39] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[39] <= perf_counter_d[39];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[38] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[38] <= perf_counter_d[38];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[37] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[37] <= perf_counter_d[37];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[36] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[36] <= perf_counter_d[36];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[35] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[35] <= perf_counter_d[35];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[34] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[34] <= perf_counter_d[34];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[33] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[33] <= perf_counter_d[33];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[32] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[32] <= perf_counter_d[32];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[31] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[31] <= perf_counter_d[31];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[30] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[30] <= perf_counter_d[30];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[29] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[29] <= perf_counter_d[29];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[28] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[28] <= perf_counter_d[28];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[27] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[27] <= perf_counter_d[27];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[26] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[26] <= perf_counter_d[26];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[25] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[25] <= perf_counter_d[25];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[24] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[24] <= perf_counter_d[24];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[23] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[23] <= perf_counter_d[23];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[22] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[22] <= perf_counter_d[22];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[21] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[21] <= perf_counter_d[21];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[20] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[20] <= perf_counter_d[20];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[19] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[19] <= perf_counter_d[19];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[18] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[18] <= perf_counter_d[18];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[17] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[17] <= perf_counter_d[17];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[16] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[16] <= perf_counter_d[16];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[15] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[15] <= perf_counter_d[15];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[14] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[14] <= perf_counter_d[14];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[13] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[13] <= perf_counter_d[13];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[12] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[12] <= perf_counter_d[12];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[11] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[11] <= perf_counter_d[11];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[10] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[10] <= perf_counter_d[10];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[9] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[9] <= perf_counter_d[9];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[8] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[8] <= perf_counter_d[8];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[7] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[7] <= perf_counter_d[7];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[6] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[6] <= perf_counter_d[6];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[5] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[5] <= perf_counter_d[5];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[4] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[4] <= perf_counter_d[4];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[3] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[3] <= perf_counter_d[3];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[2] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[2] <= perf_counter_d[2];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[1] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[1] <= perf_counter_d[1];
    end 
  end


  always @(posedge clk_i or posedge N4055) begin
    if(N4055) begin
      perf_counter_q[0] <= 1'b0;
    end else if(1'b1) begin
      perf_counter_q[0] <= perf_counter_d[0];
    end 
  end

  assign N4056 = ~commit_instr_i[293];
  assign N4057 = N4056 | commit_instr_i[294];
  assign N4058 = commit_instr_i[292] | N4057;
  assign N4059 = commit_instr_i[291] | N4058;
  assign N4060 = ~N4059;
  assign N4061 = ~commit_instr_i[292];
  assign N4062 = commit_instr_i[293] | commit_instr_i[294];
  assign N4063 = N4061 | N4062;
  assign N4064 = commit_instr_i[291] | N4063;
  assign N4065 = ~N4064;
  assign N4066 = ~commit_instr_i[291];
  assign N4067 = commit_instr_i[292] | N4062;
  assign N4068 = N4066 | N4067;
  assign N4069 = ~N4068;
  assign N4070 = ~commit_instr_i[288];
  assign N4071 = ~commit_instr_i[285];
  assign N4072 = ~commit_instr_i[284];
  assign N4073 = commit_instr_i[289] | commit_instr_i[290];
  assign N4074 = N4070 | N4073;
  assign N4075 = commit_instr_i[287] | N4074;
  assign N4076 = commit_instr_i[286] | N4075;
  assign N4077 = N4071 | N4076;
  assign N4078 = N4072 | N4077;
  assign N4079 = ~N4078;
  assign N4080 = ~commit_instr_i[278];
  assign N4081 = commit_instr_i[282] | commit_instr_i[283];
  assign N4082 = commit_instr_i[281] | N4081;
  assign N4083 = commit_instr_i[280] | N4082;
  assign N4084 = commit_instr_i[279] | N4083;
  assign N4085 = N4080 | N4084;
  assign N4086 = ~N4085;
  assign N4087 = commit_instr_i[288] | N4073;
  assign N4088 = commit_instr_i[287] | N4087;
  assign N4089 = commit_instr_i[286] | N4088;
  assign N4090 = commit_instr_i[285] | N4089;
  assign N4091 = commit_instr_i[284] | N4090;
  assign N4092 = ~N4091;
  assign N4093 = ~commit_instr_i[266];
  assign N4094 = commit_instr_i[270] | commit_instr_i[271];
  assign N4095 = commit_instr_i[269] | N4094;
  assign N4096 = commit_instr_i[268] | N4095;
  assign N4097 = commit_instr_i[267] | N4096;
  assign N4098 = N4093 | N4097;
  assign N4099 = ~N4098;
  assign { N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93 } = perf_counter_q[63:0] + 1'b1;
  assign { N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222 } = perf_counter_q[127:64] + 1'b1;
  assign { N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351 } = perf_counter_q[191:128] + 1'b1;
  assign { N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480 } = perf_counter_q[255:192] + 1'b1;
  assign { N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575 } = perf_counter_q[447:384] + 1'b1;
  assign { N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704 } = perf_counter_q[511:448] + 1'b1;
  assign { N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834 } = perf_counter_q[767:704] + 1'b1;
  assign { N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963 } = perf_counter_q[831:768] + 1'b1;
  assign { N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092 } = perf_counter_q[895:832] + 1'b1;
  assign { N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610 } = perf_counter_q[319:256] + 1'b1;
  assign { N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738 } = perf_counter_q[383:320] + 1'b1;
  assign { N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866 } = perf_counter_q[575:512] + 1'b1;
  assign { N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996 } = perf_counter_q[639:576] + 1'b1;
  assign { N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126 } = perf_counter_q[703:640] + 1'b1;
  assign N4100 = addr_i[2] & addr_i[3];
  assign N4101 = N0 & addr_i[3];
  assign N0 = ~addr_i[2];
  assign N4102 = addr_i[2] & N1;
  assign N1 = ~addr_i[3];
  assign N4103 = N2 & N3;
  assign N2 = ~addr_i[2];
  assign N3 = ~addr_i[3];
  assign N4104 = addr_i[0] & addr_i[1];
  assign N4105 = N4 & addr_i[1];
  assign N4 = ~addr_i[0];
  assign N4106 = addr_i[0] & N5;
  assign N5 = ~addr_i[1];
  assign N4107 = N6 & N7;
  assign N6 = ~addr_i[0];
  assign N7 = ~addr_i[1];
  assign N4108 = N4100 & N4104;
  assign N4109 = N4100 & N4105;
  assign N4110 = N4100 & N4106;
  assign N4111 = N4100 & N4107;
  assign N4112 = N4101 & N4104;
  assign N4113 = N4101 & N4105;
  assign N4114 = N4101 & N4106;
  assign N4115 = N4101 & N4107;
  assign N4116 = N4102 & N4104;
  assign N4117 = N4102 & N4105;
  assign N4118 = N4102 & N4106;
  assign N4119 = N4102 & N4107;
  assign N4120 = N4103 & N4104;
  assign N4121 = N4103 & N4107;
  assign N4122 = ~addr_i[4];
  assign N3131 = N4120 & N4122;
  assign N3132 = N4119 & N4122;
  assign N3133 = N4118 & N4122;
  assign N3134 = N4117 & N4122;
  assign N3135 = N4116 & N4122;
  assign N3136 = N4115 & N4122;
  assign N3137 = N4114 & N4122;
  assign N3138 = N4113 & N4122;
  assign N3139 = N4112 & N4122;
  assign N3140 = N4111 & N4122;
  assign N3141 = N4110 & N4122;
  assign N3142 = N4109 & N4122;
  assign N3143 = N4108 & N4122;
  assign N3144 = N4121 & addr_i[4];
  assign N3116 = N8 & N9 & N10;
  assign N8 = ~addr_i[3];
  assign N9 = ~addr_i[2];
  assign N10 = ~addr_i[0];
  assign N3117 = addr_i[3] & N11 & (N12 & N13);
  assign N11 = ~addr_i[2];
  assign N12 = ~addr_i[0];
  assign N13 = ~addr_i[1];
  assign N3120 = N14 & N15 & addr_i[0];
  assign N14 = ~addr_i[3];
  assign N15 = ~addr_i[2];
  assign N3122 = N16 & addr_i[2] & (N17 & N18);
  assign N16 = ~addr_i[3];
  assign N17 = ~addr_i[0];
  assign N18 = ~addr_i[1];
  assign N3124 = N19 & addr_i[0] & N20;
  assign N19 = ~addr_i[3];
  assign N20 = ~addr_i[1];
  assign N3126 = N21 & N22 & addr_i[1];
  assign N21 = ~addr_i[3];
  assign N22 = ~addr_i[0];
  assign N3128 = N23 & addr_i[2] & (addr_i[0] & addr_i[1]);
  assign N23 = ~addr_i[3];
  assign N3118 = N24 & addr_i[0] & N25;
  assign N24 = ~addr_i[2];
  assign N25 = ~addr_i[1];
  assign N3119 = N26 & N27 & addr_i[1];
  assign N26 = ~addr_i[2];
  assign N27 = ~addr_i[0];
  assign N3121 = addr_i[3] & N28 & (addr_i[0] & addr_i[1]);
  assign N28 = ~addr_i[2];
  assign N3123 = addr_i[3] & addr_i[2] & (N29 & N30);
  assign N29 = ~addr_i[0];
  assign N30 = ~addr_i[1];
  assign N3125 = addr_i[3] & addr_i[2] & (addr_i[0] & N31);
  assign N31 = ~addr_i[1];
  assign N3127 = addr_i[3] & addr_i[2] & (N32 & addr_i[1]);
  assign N32 = ~addr_i[0];
  assign N3129 = addr_i[3] & addr_i[2] & (addr_i[0] & addr_i[1]);
  assign { N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157 } = (N33)? { N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N34)? perf_counter_q[63:0] : 1'b0;
  assign N33 = l1_icache_miss_i;
  assign N34 = N92;
  assign { N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286 } = (N35)? { N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N36)? perf_counter_q[127:64] : 1'b0;
  assign N35 = l1_dcache_miss_i;
  assign N36 = N221;
  assign { N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415 } = (N37)? { N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N38)? perf_counter_q[191:128] : 1'b0;
  assign N37 = itlb_miss_i;
  assign N38 = N350;
  assign { N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544 } = (N39)? { N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N40)? perf_counter_q[255:192] : 1'b0;
  assign N39 = dtlb_miss_i;
  assign N40 = N479;
  assign { N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674 } = (N41)? { N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N42)? perf_counter_q[319:256] : 1'b0;
  assign N41 = N4069;
  assign N42 = N4068;
  assign { N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802 } = (N43)? { N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N44)? perf_counter_q[383:320] : 1'b0;
  assign N43 = N4065;
  assign N44 = N4064;
  assign { N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930 } = (N45)? { N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N46)? perf_counter_q[575:512] : 1'b0;
  assign N45 = N4060;
  assign N46 = N4059;
  assign { N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060 } = (N47)? { N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N995)? perf_counter_q[639:576] : 1'b0;
  assign N47 = N994;
  assign { N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190 } = (N48)? { N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1125)? perf_counter_q[703:640] : 1'b0;
  assign N48 = N1124;
  assign { N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254 } = (N49)? { N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N608)? { perf_counter_q[703:512], perf_counter_q[383:256] } : 1'b0;
  assign N49 = commit_ack_i[0];
  assign { N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639 } = (N50)? { N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1574)? perf_counter_q[447:384] : 1'b0;
  assign N50 = ex_i[0];
  assign { N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768 } = (N51)? { N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N52)? perf_counter_q[511:448] : 1'b0;
  assign N51 = eret_i;
  assign N52 = N1703;
  assign { N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898 } = (N53)? { N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1833)? perf_counter_q[767:704] : 1'b0;
  assign N53 = N1832;
  assign { N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027 } = (N54)? { N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N55)? perf_counter_q[831:768] : 1'b0;
  assign N54 = sb_full_i;
  assign N55 = N1962;
  assign { N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156 } = (N56)? { N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N57)? perf_counter_q[895:832] : 1'b0;
  assign N56 = if_empty_i;
  assign N57 = N2091;
  assign { N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220 } = (N58)? { N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N59)? perf_counter_q : 1'b0;
  assign N58 = N90;
  assign N59 = debug_mode_i;
  assign { N3209, N3208, N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, N3197, N3196, N3195, N3194, N3193, N3192, N3191, N3190, N3189, N3188, N3187, N3186, N3185, N3184, N3183, N3182, N3181, N3180, N3179, N3178, N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163, N3162, N3161, N3160, N3159, N3158, N3157, N3156, N3155, N3154, N3153, N3152, N3151, N3150, N3149, N3148, N3147, N3146 } = (N60)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3145)? { N2220, N2221, N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2229, N2230, N2231, N2232, N2233, N2234, N2235, N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, N2265, N2266, N2267, N2268, N2269, N2270, N2271, N2272, N2273, N2274, N2275, N2276, N2277, N2278, N2279, N2280, N2281, N2282, N2283 } : 1'b0;
  assign N60 = N3131;
  assign { N3274, N3273, N3272, N3271, N3270, N3269, N3268, N3267, N3266, N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252, N3251, N3250, N3249, N3248, N3247, N3246, N3245, N3244, N3243, N3242, N3241, N3240, N3239, N3238, N3237, N3236, N3235, N3234, N3233, N3232, N3231, N3230, N3229, N3228, N3227, N3226, N3225, N3224, N3223, N3222, N3221, N3220, N3219, N3218, N3217, N3216, N3215, N3214, N3213, N3212, N3211 } = (N61)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3210)? { N2284, N2285, N2286, N2287, N2288, N2289, N2290, N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315, N2316, N2317, N2318, N2319, N2320, N2321, N2322, N2323, N2324, N2325, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347 } : 1'b0;
  assign N61 = N3132;
  assign { N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331, N3330, N3329, N3328, N3327, N3326, N3325, N3324, N3323, N3322, N3321, N3320, N3319, N3318, N3317, N3316, N3315, N3314, N3313, N3312, N3311, N3310, N3309, N3308, N3307, N3306, N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, N3285, N3284, N3283, N3282, N3281, N3280, N3279, N3278, N3277, N3276 } = (N62)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3275)? { N2348, N2349, N2350, N2351, N2352, N2353, N2354, N2355, N2356, N2357, N2358, N2359, N2360, N2361, N2362, N2363, N2364, N2365, N2366, N2367, N2368, N2369, N2370, N2371, N2372, N2373, N2374, N2375, N2376, N2377, N2378, N2379, N2380, N2381, N2382, N2383, N2384, N2385, N2386, N2387, N2388, N2389, N2390, N2391, N2392, N2393, N2394, N2395, N2396, N2397, N2398, N2399, N2400, N2401, N2402, N2403, N2404, N2405, N2406, N2407, N2408, N2409, N2410, N2411 } : 1'b0;
  assign N62 = N3133;
  assign { N3404, N3403, N3402, N3401, N3400, N3399, N3398, N3397, N3396, N3395, N3394, N3393, N3392, N3391, N3390, N3389, N3388, N3387, N3386, N3385, N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, N3364, N3363, N3362, N3361, N3360, N3359, N3358, N3357, N3356, N3355, N3354, N3353, N3352, N3351, N3350, N3349, N3348, N3347, N3346, N3345, N3344, N3343, N3342, N3341 } = (N63)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3340)? { N2412, N2413, N2414, N2415, N2416, N2417, N2418, N2419, N2420, N2421, N2422, N2423, N2424, N2425, N2426, N2427, N2428, N2429, N2430, N2431, N2432, N2433, N2434, N2435, N2436, N2437, N2438, N2439, N2440, N2441, N2442, N2443, N2444, N2445, N2446, N2447, N2448, N2449, N2450, N2451, N2452, N2453, N2454, N2455, N2456, N2457, N2458, N2459, N2460, N2461, N2462, N2463, N2464, N2465, N2466, N2467, N2468, N2469, N2470, N2471, N2472, N2473, N2474, N2475 } : 1'b0;
  assign N63 = N3134;
  assign { N3469, N3468, N3467, N3466, N3465, N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, N3454, N3453, N3452, N3451, N3450, N3449, N3448, N3447, N3446, N3445, N3444, N3443, N3442, N3441, N3440, N3439, N3438, N3437, N3436, N3435, N3434, N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420, N3419, N3418, N3417, N3416, N3415, N3414, N3413, N3412, N3411, N3410, N3409, N3408, N3407, N3406 } = (N64)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3405)? { N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484, N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494, N2495, N2496, N2497, N2498, N2499, N2500, N2501, N2502, N2503, N2504, N2505, N2506, N2507, N2508, N2509, N2510, N2511, N2512, N2513, N2514, N2515, N2516, N2517, N2518, N2519, N2520, N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530, N2531, N2532, N2533, N2534, N2535, N2536, N2537, N2538, N2539 } : 1'b0;
  assign N64 = N3135;
  assign { N3534, N3533, N3532, N3531, N3530, N3529, N3528, N3527, N3526, N3525, N3524, N3523, N3522, N3521, N3520, N3519, N3518, N3517, N3516, N3515, N3514, N3513, N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499, N3498, N3497, N3496, N3495, N3494, N3493, N3492, N3491, N3490, N3489, N3488, N3487, N3486, N3485, N3484, N3483, N3482, N3481, N3480, N3479, N3478, N3477, N3476, N3475, N3474, N3473, N3472, N3471 } = (N65)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3470)? { N2540, N2541, N2542, N2543, N2544, N2545, N2546, N2547, N2548, N2549, N2550, N2551, N2552, N2553, N2554, N2555, N2556, N2557, N2558, N2559, N2560, N2561, N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569, N2570, N2571, N2572, N2573, N2574, N2575, N2576, N2577, N2578, N2579, N2580, N2581, N2582, N2583, N2584, N2585, N2586, N2587, N2588, N2589, N2590, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603 } : 1'b0;
  assign N65 = N3136;
  assign { N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588, N3587, N3586, N3585, N3584, N3583, N3582, N3581, N3580, N3579, N3578, N3577, N3576, N3575, N3574, N3573, N3572, N3571, N3570, N3569, N3568, N3567, N3566, N3565, N3564, N3563, N3562, N3561, N3560, N3559, N3558, N3557, N3556, N3555, N3554, N3553, N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536 } = (N66)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3535)? { N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2623, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667 } : 1'b0;
  assign N66 = N3137;
  assign { N3664, N3663, N3662, N3661, N3660, N3659, N3658, N3657, N3656, N3655, N3654, N3653, N3652, N3651, N3650, N3649, N3648, N3647, N3646, N3645, N3644, N3643, N3642, N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, N3622, N3621, N3620, N3619, N3618, N3617, N3616, N3615, N3614, N3613, N3612, N3611, N3610, N3609, N3608, N3607, N3606, N3605, N3604, N3603, N3602, N3601 } = (N67)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3600)? { N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683, N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695, N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705, N2706, N2707, N2708, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2723, N2724, N2725, N2726, N2727, N2728, N2729, N2730, N2731 } : 1'b0;
  assign N67 = N3138;
  assign { N3729, N3728, N3727, N3726, N3725, N3724, N3723, N3722, N3721, N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, N3701, N3700, N3699, N3698, N3697, N3696, N3695, N3694, N3693, N3692, N3691, N3690, N3689, N3688, N3687, N3686, N3685, N3684, N3683, N3682, N3681, N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667, N3666 } = (N68)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3665)? { N2732, N2733, N2734, N2735, N2736, N2737, N2738, N2739, N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2749, N2750, N2751, N2752, N2753, N2754, N2755, N2756, N2757, N2758, N2759, N2760, N2761, N2762, N2763, N2764, N2765, N2766, N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791, N2792, N2793, N2794, N2795 } : 1'b0;
  assign N68 = N3139;
  assign { N3794, N3793, N3792, N3791, N3790, N3789, N3788, N3787, N3786, N3785, N3784, N3783, N3782, N3781, N3780, N3779, N3778, N3777, N3776, N3775, N3774, N3773, N3772, N3771, N3770, N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756, N3755, N3754, N3753, N3752, N3751, N3750, N3749, N3748, N3747, N3746, N3745, N3744, N3743, N3742, N3741, N3740, N3739, N3738, N3737, N3736, N3735, N3734, N3733, N3732, N3731 } = (N69)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3730)? { N2796, N2797, N2798, N2799, N2800, N2801, N2802, N2803, N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811, N2812, N2813, N2814, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859 } : 1'b0;
  assign N69 = N3140;
  assign { N3859, N3858, N3857, N3856, N3855, N3854, N3853, N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838, N3837, N3836, N3835, N3834, N3833, N3832, N3831, N3830, N3829, N3828, N3827, N3826, N3825, N3824, N3823, N3822, N3821, N3820, N3819, N3818, N3817, N3816, N3815, N3814, N3813, N3812, N3811, N3810, N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, N3799, N3798, N3797, N3796 } = (N70)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3795)? { N2860, N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883, N2884, N2885, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2893, N2894, N2895, N2896, N2897, N2898, N2899, N2900, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923 } : 1'b0;
  assign N70 = N3141;
  assign { N3924, N3923, N3922, N3921, N3920, N3919, N3918, N3917, N3916, N3915, N3914, N3913, N3912, N3911, N3910, N3909, N3908, N3907, N3906, N3905, N3904, N3903, N3902, N3901, N3900, N3899, N3898, N3897, N3896, N3895, N3894, N3893, N3892, N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, N3871, N3870, N3869, N3868, N3867, N3866, N3865, N3864, N3863, N3862, N3861 } = (N71)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3860)? { N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2943, N2944, N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966, N2967, N2968, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987 } : 1'b0;
  assign N71 = N3142;
  assign { N3989, N3988, N3987, N3986, N3985, N3984, N3983, N3982, N3981, N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, N3960, N3959, N3958, N3957, N3956, N3955, N3954, N3953, N3952, N3951, N3950, N3949, N3948, N3947, N3946, N3945, N3944, N3943, N3942, N3941, N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927, N3926 } = (N72)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3925)? { N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3008, N3009, N3010, N3011, N3012, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038, N3039, N3040, N3041, N3042, N3043, N3044, N3045, N3046, N3047, N3048, N3049, N3050, N3051 } : 1'b0;
  assign N72 = N3143;
  assign { N4054, N4053, N4052, N4051, N4050, N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, N4039, N4038, N4037, N4036, N4035, N4034, N4033, N4032, N4031, N4030, N4029, N4028, N4027, N4026, N4025, N4024, N4023, N4022, N4021, N4020, N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006, N4005, N4004, N4003, N4002, N4001, N4000, N3999, N3998, N3997, N3996, N3995, N3994, N3993, N3992, N3991 } = (N73)? { data_i[0:0], data_i[1:1], data_i[2:2], data_i[3:3], data_i[4:4], data_i[5:5], data_i[6:6], data_i[7:7], data_i[8:8], data_i[9:9], data_i[10:10], data_i[11:11], data_i[12:12], data_i[13:13], data_i[14:14], data_i[15:15], data_i[16:16], data_i[17:17], data_i[18:18], data_i[19:19], data_i[20:20], data_i[21:21], data_i[22:22], data_i[23:23], data_i[24:24], data_i[25:25], data_i[26:26], data_i[27:27], data_i[28:28], data_i[29:29], data_i[30:30], data_i[31:31], data_i[32:32], data_i[33:33], data_i[34:34], data_i[35:35], data_i[36:36], data_i[37:37], data_i[38:38], data_i[39:39], data_i[40:40], data_i[41:41], data_i[42:42], data_i[43:43], data_i[44:44], data_i[45:45], data_i[46:46], data_i[47:47], data_i[48:48], data_i[49:49], data_i[50:50], data_i[51:51], data_i[52:52], data_i[53:53], data_i[54:54], data_i[55:55], data_i[56:56], data_i[57:57], data_i[58:58], data_i[59:59], data_i[60:60], data_i[61:61], data_i[62:62], data_i[63:63] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3990)? { N3052, N3053, N3054, N3055, N3056, N3057, N3058, N3059, N3060, N3061, N3062, N3063, N3064, N3065, N3066, N3067, N3068, N3069, N3070, N3071, N3072, N3073, N3074, N3075, N3076, N3077, N3078, N3079, N3080, N3081, N3082, N3083, N3084, N3085, N3086, N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096, N3097, N3098, N3099, N3100, N3101, N3102, N3103, N3104, N3105, N3106, N3107, N3108, N3109, N3110, N3111, N3112, N3113, N3114, N3115 } : 1'b0;
  assign N73 = N3144;
  assign perf_counter_d = (N74)? { N3991, N3992, N3993, N3994, N3995, N3996, N3997, N3998, N3999, N4000, N4001, N4002, N4003, N4004, N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4022, N4023, N4024, N4025, N4026, N4027, N4028, N4029, N4030, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051, N4052, N4053, N4054, N3926, N3927, N3928, N3929, N3930, N3931, N3932, N3933, N3934, N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942, N3943, N3944, N3945, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N3953, N3954, N3955, N3956, N3957, N3958, N3959, N3960, N3961, N3962, N3963, N3964, N3965, N3966, N3967, N3968, N3969, N3970, N3971, N3972, N3973, N3974, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3985, N3986, N3987, N3988, N3989, N3861, N3862, N3863, N3864, N3865, N3866, N3867, N3868, N3869, N3870, N3871, N3872, N3873, N3874, N3875, N3876, N3877, N3878, N3879, N3880, N3881, N3882, N3883, N3884, N3885, N3886, N3887, N3888, N3889, N3890, N3891, N3892, N3893, N3894, N3895, N3896, N3897, N3898, N3899, N3900, N3901, N3902, N3903, N3904, N3905, N3906, N3907, N3908, N3909, N3910, N3911, N3912, N3913, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3922, N3923, N3924, N3796, N3797, N3798, N3799, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3811, N3812, N3813, N3814, N3815, N3816, N3817, N3818, N3819, N3820, N3821, N3822, N3823, N3824, N3825, N3826, N3827, N3828, N3829, N3830, N3831, N3832, N3833, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3843, N3844, N3845, N3846, N3847, N3848, N3849, N3850, N3851, N3852, N3853, N3854, N3855, N3856, N3857, N3858, N3859, N3731, N3732, N3733, N3734, N3735, N3736, N3737, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3772, N3773, N3774, N3775, N3776, N3777, N3778, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3790, N3791, N3792, N3793, N3794, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3690, N3691, N3692, N3693, N3694, N3695, N3696, N3697, N3698, N3699, N3700, N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709, N3710, N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3601, N3602, N3603, N3604, N3605, N3606, N3607, N3608, N3609, N3610, N3611, N3612, N3613, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3536, N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546, N3547, N3548, N3549, N3550, N3551, N3552, N3553, N3554, N3555, N3556, N3557, N3558, N3559, N3560, N3561, N3562, N3563, N3564, N3565, N3566, N3567, N3568, N3569, N3570, N3571, N3572, N3573, N3574, N3575, N3576, N3577, N3578, N3579, N3580, N3581, N3582, N3583, N3584, N3585, N3586, N3587, N3588, N3589, N3590, N3591, N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3471, N3472, N3473, N3474, N3475, N3476, N3477, N3478, N3479, N3480, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3494, N3495, N3496, N3497, N3498, N3499, N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3516, N3517, N3518, N3519, N3520, N3521, N3522, N3523, N3524, N3525, N3526, N3527, N3528, N3529, N3530, N3531, N3532, N3533, N3534, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3417, N3418, N3419, N3420, N3421, N3422, N3423, N3424, N3425, N3426, N3427, N3428, N3429, N3430, N3431, N3432, N3433, N3434, N3435, N3436, N3437, N3438, N3439, N3440, N3441, N3442, N3443, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3467, N3468, N3469, N3341, N3342, N3343, N3344, N3345, N3346, N3347, N3348, N3349, N3350, N3351, N3352, N3353, N3354, N3355, N3356, N3357, N3358, N3359, N3360, N3361, N3362, N3363, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372, N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382, N3383, N3384, N3385, N3386, N3387, N3388, N3389, N3390, N3391, N3392, N3393, N3394, N3395, N3396, N3397, N3398, N3399, N3400, N3401, N3402, N3403, N3404, N3276, N3277, N3278, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3211, N3212, N3213, N3214, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270, N3271, N3272, N3273, N3274, N3146, N3147, N3148, N3149, N3150, N3151, N3152, N3153, N3154, N3155, N3156, N3157, N3158, N3159, N3160, N3161, N3162, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171, N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3179, N3180, N3181, N3182, N3183, N3184, N3185, N3186, N3187, N3188, N3189, N3190, N3191, N3192, N3193, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208, N3209 } : 
                          (N75)? { N3115, N3114, N3113, N3112, N3111, N3110, N3109, N3108, N3107, N3106, N3105, N3104, N3103, N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220 } : 1'b0;
  assign N74 = we_i;
  assign N75 = N3130;
  assign data_o[63] = (N76)? perf_counter_q[895] : 
                      (N77)? perf_counter_q[63] : 
                      (N78)? perf_counter_q[127] : 
                      (N79)? perf_counter_q[191] : 
                      (N80)? perf_counter_q[255] : 
                      (N81)? perf_counter_q[319] : 
                      (N82)? perf_counter_q[383] : 
                      (N83)? perf_counter_q[447] : 
                      (N84)? perf_counter_q[511] : 
                      (N85)? perf_counter_q[575] : 
                      (N86)? perf_counter_q[639] : 
                      (N87)? perf_counter_q[703] : 
                      (N88)? perf_counter_q[767] : 
                      (N89)? perf_counter_q[831] : 1'b0;
  assign N76 = N3116;
  assign N77 = N3120;
  assign N78 = N3122;
  assign N79 = N3124;
  assign N80 = N3126;
  assign N81 = N3128;
  assign N82 = N3117;
  assign N83 = N3118;
  assign N84 = N3119;
  assign N85 = N3121;
  assign N86 = N3123;
  assign N87 = N3125;
  assign N88 = N3127;
  assign N89 = N3129;
  assign data_o[62] = (N76)? perf_counter_q[894] : 
                      (N77)? perf_counter_q[62] : 
                      (N78)? perf_counter_q[126] : 
                      (N79)? perf_counter_q[190] : 
                      (N80)? perf_counter_q[254] : 
                      (N81)? perf_counter_q[318] : 
                      (N82)? perf_counter_q[382] : 
                      (N83)? perf_counter_q[446] : 
                      (N84)? perf_counter_q[510] : 
                      (N85)? perf_counter_q[574] : 
                      (N86)? perf_counter_q[638] : 
                      (N87)? perf_counter_q[702] : 
                      (N88)? perf_counter_q[766] : 
                      (N89)? perf_counter_q[830] : 1'b0;
  assign data_o[61] = (N76)? perf_counter_q[893] : 
                      (N77)? perf_counter_q[61] : 
                      (N78)? perf_counter_q[125] : 
                      (N79)? perf_counter_q[189] : 
                      (N80)? perf_counter_q[253] : 
                      (N81)? perf_counter_q[317] : 
                      (N82)? perf_counter_q[381] : 
                      (N83)? perf_counter_q[445] : 
                      (N84)? perf_counter_q[509] : 
                      (N85)? perf_counter_q[573] : 
                      (N86)? perf_counter_q[637] : 
                      (N87)? perf_counter_q[701] : 
                      (N88)? perf_counter_q[765] : 
                      (N89)? perf_counter_q[829] : 1'b0;
  assign data_o[60] = (N76)? perf_counter_q[892] : 
                      (N77)? perf_counter_q[60] : 
                      (N78)? perf_counter_q[124] : 
                      (N79)? perf_counter_q[188] : 
                      (N80)? perf_counter_q[252] : 
                      (N81)? perf_counter_q[316] : 
                      (N82)? perf_counter_q[380] : 
                      (N83)? perf_counter_q[444] : 
                      (N84)? perf_counter_q[508] : 
                      (N85)? perf_counter_q[572] : 
                      (N86)? perf_counter_q[636] : 
                      (N87)? perf_counter_q[700] : 
                      (N88)? perf_counter_q[764] : 
                      (N89)? perf_counter_q[828] : 1'b0;
  assign data_o[59] = (N76)? perf_counter_q[891] : 
                      (N77)? perf_counter_q[59] : 
                      (N78)? perf_counter_q[123] : 
                      (N79)? perf_counter_q[187] : 
                      (N80)? perf_counter_q[251] : 
                      (N81)? perf_counter_q[315] : 
                      (N82)? perf_counter_q[379] : 
                      (N83)? perf_counter_q[443] : 
                      (N84)? perf_counter_q[507] : 
                      (N85)? perf_counter_q[571] : 
                      (N86)? perf_counter_q[635] : 
                      (N87)? perf_counter_q[699] : 
                      (N88)? perf_counter_q[763] : 
                      (N89)? perf_counter_q[827] : 1'b0;
  assign data_o[58] = (N76)? perf_counter_q[890] : 
                      (N77)? perf_counter_q[58] : 
                      (N78)? perf_counter_q[122] : 
                      (N79)? perf_counter_q[186] : 
                      (N80)? perf_counter_q[250] : 
                      (N81)? perf_counter_q[314] : 
                      (N82)? perf_counter_q[378] : 
                      (N83)? perf_counter_q[442] : 
                      (N84)? perf_counter_q[506] : 
                      (N85)? perf_counter_q[570] : 
                      (N86)? perf_counter_q[634] : 
                      (N87)? perf_counter_q[698] : 
                      (N88)? perf_counter_q[762] : 
                      (N89)? perf_counter_q[826] : 1'b0;
  assign data_o[57] = (N76)? perf_counter_q[889] : 
                      (N77)? perf_counter_q[57] : 
                      (N78)? perf_counter_q[121] : 
                      (N79)? perf_counter_q[185] : 
                      (N80)? perf_counter_q[249] : 
                      (N81)? perf_counter_q[313] : 
                      (N82)? perf_counter_q[377] : 
                      (N83)? perf_counter_q[441] : 
                      (N84)? perf_counter_q[505] : 
                      (N85)? perf_counter_q[569] : 
                      (N86)? perf_counter_q[633] : 
                      (N87)? perf_counter_q[697] : 
                      (N88)? perf_counter_q[761] : 
                      (N89)? perf_counter_q[825] : 1'b0;
  assign data_o[56] = (N76)? perf_counter_q[888] : 
                      (N77)? perf_counter_q[56] : 
                      (N78)? perf_counter_q[120] : 
                      (N79)? perf_counter_q[184] : 
                      (N80)? perf_counter_q[248] : 
                      (N81)? perf_counter_q[312] : 
                      (N82)? perf_counter_q[376] : 
                      (N83)? perf_counter_q[440] : 
                      (N84)? perf_counter_q[504] : 
                      (N85)? perf_counter_q[568] : 
                      (N86)? perf_counter_q[632] : 
                      (N87)? perf_counter_q[696] : 
                      (N88)? perf_counter_q[760] : 
                      (N89)? perf_counter_q[824] : 1'b0;
  assign data_o[55] = (N76)? perf_counter_q[887] : 
                      (N77)? perf_counter_q[55] : 
                      (N78)? perf_counter_q[119] : 
                      (N79)? perf_counter_q[183] : 
                      (N80)? perf_counter_q[247] : 
                      (N81)? perf_counter_q[311] : 
                      (N82)? perf_counter_q[375] : 
                      (N83)? perf_counter_q[439] : 
                      (N84)? perf_counter_q[503] : 
                      (N85)? perf_counter_q[567] : 
                      (N86)? perf_counter_q[631] : 
                      (N87)? perf_counter_q[695] : 
                      (N88)? perf_counter_q[759] : 
                      (N89)? perf_counter_q[823] : 1'b0;
  assign data_o[54] = (N76)? perf_counter_q[886] : 
                      (N77)? perf_counter_q[54] : 
                      (N78)? perf_counter_q[118] : 
                      (N79)? perf_counter_q[182] : 
                      (N80)? perf_counter_q[246] : 
                      (N81)? perf_counter_q[310] : 
                      (N82)? perf_counter_q[374] : 
                      (N83)? perf_counter_q[438] : 
                      (N84)? perf_counter_q[502] : 
                      (N85)? perf_counter_q[566] : 
                      (N86)? perf_counter_q[630] : 
                      (N87)? perf_counter_q[694] : 
                      (N88)? perf_counter_q[758] : 
                      (N89)? perf_counter_q[822] : 1'b0;
  assign data_o[53] = (N76)? perf_counter_q[885] : 
                      (N77)? perf_counter_q[53] : 
                      (N78)? perf_counter_q[117] : 
                      (N79)? perf_counter_q[181] : 
                      (N80)? perf_counter_q[245] : 
                      (N81)? perf_counter_q[309] : 
                      (N82)? perf_counter_q[373] : 
                      (N83)? perf_counter_q[437] : 
                      (N84)? perf_counter_q[501] : 
                      (N85)? perf_counter_q[565] : 
                      (N86)? perf_counter_q[629] : 
                      (N87)? perf_counter_q[693] : 
                      (N88)? perf_counter_q[757] : 
                      (N89)? perf_counter_q[821] : 1'b0;
  assign data_o[52] = (N76)? perf_counter_q[884] : 
                      (N77)? perf_counter_q[52] : 
                      (N78)? perf_counter_q[116] : 
                      (N79)? perf_counter_q[180] : 
                      (N80)? perf_counter_q[244] : 
                      (N81)? perf_counter_q[308] : 
                      (N82)? perf_counter_q[372] : 
                      (N83)? perf_counter_q[436] : 
                      (N84)? perf_counter_q[500] : 
                      (N85)? perf_counter_q[564] : 
                      (N86)? perf_counter_q[628] : 
                      (N87)? perf_counter_q[692] : 
                      (N88)? perf_counter_q[756] : 
                      (N89)? perf_counter_q[820] : 1'b0;
  assign data_o[51] = (N76)? perf_counter_q[883] : 
                      (N77)? perf_counter_q[51] : 
                      (N78)? perf_counter_q[115] : 
                      (N79)? perf_counter_q[179] : 
                      (N80)? perf_counter_q[243] : 
                      (N81)? perf_counter_q[307] : 
                      (N82)? perf_counter_q[371] : 
                      (N83)? perf_counter_q[435] : 
                      (N84)? perf_counter_q[499] : 
                      (N85)? perf_counter_q[563] : 
                      (N86)? perf_counter_q[627] : 
                      (N87)? perf_counter_q[691] : 
                      (N88)? perf_counter_q[755] : 
                      (N89)? perf_counter_q[819] : 1'b0;
  assign data_o[50] = (N76)? perf_counter_q[882] : 
                      (N77)? perf_counter_q[50] : 
                      (N78)? perf_counter_q[114] : 
                      (N79)? perf_counter_q[178] : 
                      (N80)? perf_counter_q[242] : 
                      (N81)? perf_counter_q[306] : 
                      (N82)? perf_counter_q[370] : 
                      (N83)? perf_counter_q[434] : 
                      (N84)? perf_counter_q[498] : 
                      (N85)? perf_counter_q[562] : 
                      (N86)? perf_counter_q[626] : 
                      (N87)? perf_counter_q[690] : 
                      (N88)? perf_counter_q[754] : 
                      (N89)? perf_counter_q[818] : 1'b0;
  assign data_o[49] = (N76)? perf_counter_q[881] : 
                      (N77)? perf_counter_q[49] : 
                      (N78)? perf_counter_q[113] : 
                      (N79)? perf_counter_q[177] : 
                      (N80)? perf_counter_q[241] : 
                      (N81)? perf_counter_q[305] : 
                      (N82)? perf_counter_q[369] : 
                      (N83)? perf_counter_q[433] : 
                      (N84)? perf_counter_q[497] : 
                      (N85)? perf_counter_q[561] : 
                      (N86)? perf_counter_q[625] : 
                      (N87)? perf_counter_q[689] : 
                      (N88)? perf_counter_q[753] : 
                      (N89)? perf_counter_q[817] : 1'b0;
  assign data_o[48] = (N76)? perf_counter_q[880] : 
                      (N77)? perf_counter_q[48] : 
                      (N78)? perf_counter_q[112] : 
                      (N79)? perf_counter_q[176] : 
                      (N80)? perf_counter_q[240] : 
                      (N81)? perf_counter_q[304] : 
                      (N82)? perf_counter_q[368] : 
                      (N83)? perf_counter_q[432] : 
                      (N84)? perf_counter_q[496] : 
                      (N85)? perf_counter_q[560] : 
                      (N86)? perf_counter_q[624] : 
                      (N87)? perf_counter_q[688] : 
                      (N88)? perf_counter_q[752] : 
                      (N89)? perf_counter_q[816] : 1'b0;
  assign data_o[47] = (N76)? perf_counter_q[879] : 
                      (N77)? perf_counter_q[47] : 
                      (N78)? perf_counter_q[111] : 
                      (N79)? perf_counter_q[175] : 
                      (N80)? perf_counter_q[239] : 
                      (N81)? perf_counter_q[303] : 
                      (N82)? perf_counter_q[367] : 
                      (N83)? perf_counter_q[431] : 
                      (N84)? perf_counter_q[495] : 
                      (N85)? perf_counter_q[559] : 
                      (N86)? perf_counter_q[623] : 
                      (N87)? perf_counter_q[687] : 
                      (N88)? perf_counter_q[751] : 
                      (N89)? perf_counter_q[815] : 1'b0;
  assign data_o[46] = (N76)? perf_counter_q[878] : 
                      (N77)? perf_counter_q[46] : 
                      (N78)? perf_counter_q[110] : 
                      (N79)? perf_counter_q[174] : 
                      (N80)? perf_counter_q[238] : 
                      (N81)? perf_counter_q[302] : 
                      (N82)? perf_counter_q[366] : 
                      (N83)? perf_counter_q[430] : 
                      (N84)? perf_counter_q[494] : 
                      (N85)? perf_counter_q[558] : 
                      (N86)? perf_counter_q[622] : 
                      (N87)? perf_counter_q[686] : 
                      (N88)? perf_counter_q[750] : 
                      (N89)? perf_counter_q[814] : 1'b0;
  assign data_o[45] = (N76)? perf_counter_q[877] : 
                      (N77)? perf_counter_q[45] : 
                      (N78)? perf_counter_q[109] : 
                      (N79)? perf_counter_q[173] : 
                      (N80)? perf_counter_q[237] : 
                      (N81)? perf_counter_q[301] : 
                      (N82)? perf_counter_q[365] : 
                      (N83)? perf_counter_q[429] : 
                      (N84)? perf_counter_q[493] : 
                      (N85)? perf_counter_q[557] : 
                      (N86)? perf_counter_q[621] : 
                      (N87)? perf_counter_q[685] : 
                      (N88)? perf_counter_q[749] : 
                      (N89)? perf_counter_q[813] : 1'b0;
  assign data_o[44] = (N76)? perf_counter_q[876] : 
                      (N77)? perf_counter_q[44] : 
                      (N78)? perf_counter_q[108] : 
                      (N79)? perf_counter_q[172] : 
                      (N80)? perf_counter_q[236] : 
                      (N81)? perf_counter_q[300] : 
                      (N82)? perf_counter_q[364] : 
                      (N83)? perf_counter_q[428] : 
                      (N84)? perf_counter_q[492] : 
                      (N85)? perf_counter_q[556] : 
                      (N86)? perf_counter_q[620] : 
                      (N87)? perf_counter_q[684] : 
                      (N88)? perf_counter_q[748] : 
                      (N89)? perf_counter_q[812] : 1'b0;
  assign data_o[43] = (N76)? perf_counter_q[875] : 
                      (N77)? perf_counter_q[43] : 
                      (N78)? perf_counter_q[107] : 
                      (N79)? perf_counter_q[171] : 
                      (N80)? perf_counter_q[235] : 
                      (N81)? perf_counter_q[299] : 
                      (N82)? perf_counter_q[363] : 
                      (N83)? perf_counter_q[427] : 
                      (N84)? perf_counter_q[491] : 
                      (N85)? perf_counter_q[555] : 
                      (N86)? perf_counter_q[619] : 
                      (N87)? perf_counter_q[683] : 
                      (N88)? perf_counter_q[747] : 
                      (N89)? perf_counter_q[811] : 1'b0;
  assign data_o[42] = (N76)? perf_counter_q[874] : 
                      (N77)? perf_counter_q[42] : 
                      (N78)? perf_counter_q[106] : 
                      (N79)? perf_counter_q[170] : 
                      (N80)? perf_counter_q[234] : 
                      (N81)? perf_counter_q[298] : 
                      (N82)? perf_counter_q[362] : 
                      (N83)? perf_counter_q[426] : 
                      (N84)? perf_counter_q[490] : 
                      (N85)? perf_counter_q[554] : 
                      (N86)? perf_counter_q[618] : 
                      (N87)? perf_counter_q[682] : 
                      (N88)? perf_counter_q[746] : 
                      (N89)? perf_counter_q[810] : 1'b0;
  assign data_o[41] = (N76)? perf_counter_q[873] : 
                      (N77)? perf_counter_q[41] : 
                      (N78)? perf_counter_q[105] : 
                      (N79)? perf_counter_q[169] : 
                      (N80)? perf_counter_q[233] : 
                      (N81)? perf_counter_q[297] : 
                      (N82)? perf_counter_q[361] : 
                      (N83)? perf_counter_q[425] : 
                      (N84)? perf_counter_q[489] : 
                      (N85)? perf_counter_q[553] : 
                      (N86)? perf_counter_q[617] : 
                      (N87)? perf_counter_q[681] : 
                      (N88)? perf_counter_q[745] : 
                      (N89)? perf_counter_q[809] : 1'b0;
  assign data_o[40] = (N76)? perf_counter_q[872] : 
                      (N77)? perf_counter_q[40] : 
                      (N78)? perf_counter_q[104] : 
                      (N79)? perf_counter_q[168] : 
                      (N80)? perf_counter_q[232] : 
                      (N81)? perf_counter_q[296] : 
                      (N82)? perf_counter_q[360] : 
                      (N83)? perf_counter_q[424] : 
                      (N84)? perf_counter_q[488] : 
                      (N85)? perf_counter_q[552] : 
                      (N86)? perf_counter_q[616] : 
                      (N87)? perf_counter_q[680] : 
                      (N88)? perf_counter_q[744] : 
                      (N89)? perf_counter_q[808] : 1'b0;
  assign data_o[39] = (N76)? perf_counter_q[871] : 
                      (N77)? perf_counter_q[39] : 
                      (N78)? perf_counter_q[103] : 
                      (N79)? perf_counter_q[167] : 
                      (N80)? perf_counter_q[231] : 
                      (N81)? perf_counter_q[295] : 
                      (N82)? perf_counter_q[359] : 
                      (N83)? perf_counter_q[423] : 
                      (N84)? perf_counter_q[487] : 
                      (N85)? perf_counter_q[551] : 
                      (N86)? perf_counter_q[615] : 
                      (N87)? perf_counter_q[679] : 
                      (N88)? perf_counter_q[743] : 
                      (N89)? perf_counter_q[807] : 1'b0;
  assign data_o[38] = (N76)? perf_counter_q[870] : 
                      (N77)? perf_counter_q[38] : 
                      (N78)? perf_counter_q[102] : 
                      (N79)? perf_counter_q[166] : 
                      (N80)? perf_counter_q[230] : 
                      (N81)? perf_counter_q[294] : 
                      (N82)? perf_counter_q[358] : 
                      (N83)? perf_counter_q[422] : 
                      (N84)? perf_counter_q[486] : 
                      (N85)? perf_counter_q[550] : 
                      (N86)? perf_counter_q[614] : 
                      (N87)? perf_counter_q[678] : 
                      (N88)? perf_counter_q[742] : 
                      (N89)? perf_counter_q[806] : 1'b0;
  assign data_o[37] = (N76)? perf_counter_q[869] : 
                      (N77)? perf_counter_q[37] : 
                      (N78)? perf_counter_q[101] : 
                      (N79)? perf_counter_q[165] : 
                      (N80)? perf_counter_q[229] : 
                      (N81)? perf_counter_q[293] : 
                      (N82)? perf_counter_q[357] : 
                      (N83)? perf_counter_q[421] : 
                      (N84)? perf_counter_q[485] : 
                      (N85)? perf_counter_q[549] : 
                      (N86)? perf_counter_q[613] : 
                      (N87)? perf_counter_q[677] : 
                      (N88)? perf_counter_q[741] : 
                      (N89)? perf_counter_q[805] : 1'b0;
  assign data_o[36] = (N76)? perf_counter_q[868] : 
                      (N77)? perf_counter_q[36] : 
                      (N78)? perf_counter_q[100] : 
                      (N79)? perf_counter_q[164] : 
                      (N80)? perf_counter_q[228] : 
                      (N81)? perf_counter_q[292] : 
                      (N82)? perf_counter_q[356] : 
                      (N83)? perf_counter_q[420] : 
                      (N84)? perf_counter_q[484] : 
                      (N85)? perf_counter_q[548] : 
                      (N86)? perf_counter_q[612] : 
                      (N87)? perf_counter_q[676] : 
                      (N88)? perf_counter_q[740] : 
                      (N89)? perf_counter_q[804] : 1'b0;
  assign data_o[35] = (N76)? perf_counter_q[867] : 
                      (N77)? perf_counter_q[35] : 
                      (N78)? perf_counter_q[99] : 
                      (N79)? perf_counter_q[163] : 
                      (N80)? perf_counter_q[227] : 
                      (N81)? perf_counter_q[291] : 
                      (N82)? perf_counter_q[355] : 
                      (N83)? perf_counter_q[419] : 
                      (N84)? perf_counter_q[483] : 
                      (N85)? perf_counter_q[547] : 
                      (N86)? perf_counter_q[611] : 
                      (N87)? perf_counter_q[675] : 
                      (N88)? perf_counter_q[739] : 
                      (N89)? perf_counter_q[803] : 1'b0;
  assign data_o[34] = (N76)? perf_counter_q[866] : 
                      (N77)? perf_counter_q[34] : 
                      (N78)? perf_counter_q[98] : 
                      (N79)? perf_counter_q[162] : 
                      (N80)? perf_counter_q[226] : 
                      (N81)? perf_counter_q[290] : 
                      (N82)? perf_counter_q[354] : 
                      (N83)? perf_counter_q[418] : 
                      (N84)? perf_counter_q[482] : 
                      (N85)? perf_counter_q[546] : 
                      (N86)? perf_counter_q[610] : 
                      (N87)? perf_counter_q[674] : 
                      (N88)? perf_counter_q[738] : 
                      (N89)? perf_counter_q[802] : 1'b0;
  assign data_o[33] = (N76)? perf_counter_q[865] : 
                      (N77)? perf_counter_q[33] : 
                      (N78)? perf_counter_q[97] : 
                      (N79)? perf_counter_q[161] : 
                      (N80)? perf_counter_q[225] : 
                      (N81)? perf_counter_q[289] : 
                      (N82)? perf_counter_q[353] : 
                      (N83)? perf_counter_q[417] : 
                      (N84)? perf_counter_q[481] : 
                      (N85)? perf_counter_q[545] : 
                      (N86)? perf_counter_q[609] : 
                      (N87)? perf_counter_q[673] : 
                      (N88)? perf_counter_q[737] : 
                      (N89)? perf_counter_q[801] : 1'b0;
  assign data_o[32] = (N76)? perf_counter_q[864] : 
                      (N77)? perf_counter_q[32] : 
                      (N78)? perf_counter_q[96] : 
                      (N79)? perf_counter_q[160] : 
                      (N80)? perf_counter_q[224] : 
                      (N81)? perf_counter_q[288] : 
                      (N82)? perf_counter_q[352] : 
                      (N83)? perf_counter_q[416] : 
                      (N84)? perf_counter_q[480] : 
                      (N85)? perf_counter_q[544] : 
                      (N86)? perf_counter_q[608] : 
                      (N87)? perf_counter_q[672] : 
                      (N88)? perf_counter_q[736] : 
                      (N89)? perf_counter_q[800] : 1'b0;
  assign data_o[31] = (N76)? perf_counter_q[863] : 
                      (N77)? perf_counter_q[31] : 
                      (N78)? perf_counter_q[95] : 
                      (N79)? perf_counter_q[159] : 
                      (N80)? perf_counter_q[223] : 
                      (N81)? perf_counter_q[287] : 
                      (N82)? perf_counter_q[351] : 
                      (N83)? perf_counter_q[415] : 
                      (N84)? perf_counter_q[479] : 
                      (N85)? perf_counter_q[543] : 
                      (N86)? perf_counter_q[607] : 
                      (N87)? perf_counter_q[671] : 
                      (N88)? perf_counter_q[735] : 
                      (N89)? perf_counter_q[799] : 1'b0;
  assign data_o[30] = (N76)? perf_counter_q[862] : 
                      (N77)? perf_counter_q[30] : 
                      (N78)? perf_counter_q[94] : 
                      (N79)? perf_counter_q[158] : 
                      (N80)? perf_counter_q[222] : 
                      (N81)? perf_counter_q[286] : 
                      (N82)? perf_counter_q[350] : 
                      (N83)? perf_counter_q[414] : 
                      (N84)? perf_counter_q[478] : 
                      (N85)? perf_counter_q[542] : 
                      (N86)? perf_counter_q[606] : 
                      (N87)? perf_counter_q[670] : 
                      (N88)? perf_counter_q[734] : 
                      (N89)? perf_counter_q[798] : 1'b0;
  assign data_o[29] = (N76)? perf_counter_q[861] : 
                      (N77)? perf_counter_q[29] : 
                      (N78)? perf_counter_q[93] : 
                      (N79)? perf_counter_q[157] : 
                      (N80)? perf_counter_q[221] : 
                      (N81)? perf_counter_q[285] : 
                      (N82)? perf_counter_q[349] : 
                      (N83)? perf_counter_q[413] : 
                      (N84)? perf_counter_q[477] : 
                      (N85)? perf_counter_q[541] : 
                      (N86)? perf_counter_q[605] : 
                      (N87)? perf_counter_q[669] : 
                      (N88)? perf_counter_q[733] : 
                      (N89)? perf_counter_q[797] : 1'b0;
  assign data_o[28] = (N76)? perf_counter_q[860] : 
                      (N77)? perf_counter_q[28] : 
                      (N78)? perf_counter_q[92] : 
                      (N79)? perf_counter_q[156] : 
                      (N80)? perf_counter_q[220] : 
                      (N81)? perf_counter_q[284] : 
                      (N82)? perf_counter_q[348] : 
                      (N83)? perf_counter_q[412] : 
                      (N84)? perf_counter_q[476] : 
                      (N85)? perf_counter_q[540] : 
                      (N86)? perf_counter_q[604] : 
                      (N87)? perf_counter_q[668] : 
                      (N88)? perf_counter_q[732] : 
                      (N89)? perf_counter_q[796] : 1'b0;
  assign data_o[27] = (N76)? perf_counter_q[859] : 
                      (N77)? perf_counter_q[27] : 
                      (N78)? perf_counter_q[91] : 
                      (N79)? perf_counter_q[155] : 
                      (N80)? perf_counter_q[219] : 
                      (N81)? perf_counter_q[283] : 
                      (N82)? perf_counter_q[347] : 
                      (N83)? perf_counter_q[411] : 
                      (N84)? perf_counter_q[475] : 
                      (N85)? perf_counter_q[539] : 
                      (N86)? perf_counter_q[603] : 
                      (N87)? perf_counter_q[667] : 
                      (N88)? perf_counter_q[731] : 
                      (N89)? perf_counter_q[795] : 1'b0;
  assign data_o[26] = (N76)? perf_counter_q[858] : 
                      (N77)? perf_counter_q[26] : 
                      (N78)? perf_counter_q[90] : 
                      (N79)? perf_counter_q[154] : 
                      (N80)? perf_counter_q[218] : 
                      (N81)? perf_counter_q[282] : 
                      (N82)? perf_counter_q[346] : 
                      (N83)? perf_counter_q[410] : 
                      (N84)? perf_counter_q[474] : 
                      (N85)? perf_counter_q[538] : 
                      (N86)? perf_counter_q[602] : 
                      (N87)? perf_counter_q[666] : 
                      (N88)? perf_counter_q[730] : 
                      (N89)? perf_counter_q[794] : 1'b0;
  assign data_o[25] = (N76)? perf_counter_q[857] : 
                      (N77)? perf_counter_q[25] : 
                      (N78)? perf_counter_q[89] : 
                      (N79)? perf_counter_q[153] : 
                      (N80)? perf_counter_q[217] : 
                      (N81)? perf_counter_q[281] : 
                      (N82)? perf_counter_q[345] : 
                      (N83)? perf_counter_q[409] : 
                      (N84)? perf_counter_q[473] : 
                      (N85)? perf_counter_q[537] : 
                      (N86)? perf_counter_q[601] : 
                      (N87)? perf_counter_q[665] : 
                      (N88)? perf_counter_q[729] : 
                      (N89)? perf_counter_q[793] : 1'b0;
  assign data_o[24] = (N76)? perf_counter_q[856] : 
                      (N77)? perf_counter_q[24] : 
                      (N78)? perf_counter_q[88] : 
                      (N79)? perf_counter_q[152] : 
                      (N80)? perf_counter_q[216] : 
                      (N81)? perf_counter_q[280] : 
                      (N82)? perf_counter_q[344] : 
                      (N83)? perf_counter_q[408] : 
                      (N84)? perf_counter_q[472] : 
                      (N85)? perf_counter_q[536] : 
                      (N86)? perf_counter_q[600] : 
                      (N87)? perf_counter_q[664] : 
                      (N88)? perf_counter_q[728] : 
                      (N89)? perf_counter_q[792] : 1'b0;
  assign data_o[23] = (N76)? perf_counter_q[855] : 
                      (N77)? perf_counter_q[23] : 
                      (N78)? perf_counter_q[87] : 
                      (N79)? perf_counter_q[151] : 
                      (N80)? perf_counter_q[215] : 
                      (N81)? perf_counter_q[279] : 
                      (N82)? perf_counter_q[343] : 
                      (N83)? perf_counter_q[407] : 
                      (N84)? perf_counter_q[471] : 
                      (N85)? perf_counter_q[535] : 
                      (N86)? perf_counter_q[599] : 
                      (N87)? perf_counter_q[663] : 
                      (N88)? perf_counter_q[727] : 
                      (N89)? perf_counter_q[791] : 1'b0;
  assign data_o[22] = (N76)? perf_counter_q[854] : 
                      (N77)? perf_counter_q[22] : 
                      (N78)? perf_counter_q[86] : 
                      (N79)? perf_counter_q[150] : 
                      (N80)? perf_counter_q[214] : 
                      (N81)? perf_counter_q[278] : 
                      (N82)? perf_counter_q[342] : 
                      (N83)? perf_counter_q[406] : 
                      (N84)? perf_counter_q[470] : 
                      (N85)? perf_counter_q[534] : 
                      (N86)? perf_counter_q[598] : 
                      (N87)? perf_counter_q[662] : 
                      (N88)? perf_counter_q[726] : 
                      (N89)? perf_counter_q[790] : 1'b0;
  assign data_o[21] = (N76)? perf_counter_q[853] : 
                      (N77)? perf_counter_q[21] : 
                      (N78)? perf_counter_q[85] : 
                      (N79)? perf_counter_q[149] : 
                      (N80)? perf_counter_q[213] : 
                      (N81)? perf_counter_q[277] : 
                      (N82)? perf_counter_q[341] : 
                      (N83)? perf_counter_q[405] : 
                      (N84)? perf_counter_q[469] : 
                      (N85)? perf_counter_q[533] : 
                      (N86)? perf_counter_q[597] : 
                      (N87)? perf_counter_q[661] : 
                      (N88)? perf_counter_q[725] : 
                      (N89)? perf_counter_q[789] : 1'b0;
  assign data_o[20] = (N76)? perf_counter_q[852] : 
                      (N77)? perf_counter_q[20] : 
                      (N78)? perf_counter_q[84] : 
                      (N79)? perf_counter_q[148] : 
                      (N80)? perf_counter_q[212] : 
                      (N81)? perf_counter_q[276] : 
                      (N82)? perf_counter_q[340] : 
                      (N83)? perf_counter_q[404] : 
                      (N84)? perf_counter_q[468] : 
                      (N85)? perf_counter_q[532] : 
                      (N86)? perf_counter_q[596] : 
                      (N87)? perf_counter_q[660] : 
                      (N88)? perf_counter_q[724] : 
                      (N89)? perf_counter_q[788] : 1'b0;
  assign data_o[19] = (N76)? perf_counter_q[851] : 
                      (N77)? perf_counter_q[19] : 
                      (N78)? perf_counter_q[83] : 
                      (N79)? perf_counter_q[147] : 
                      (N80)? perf_counter_q[211] : 
                      (N81)? perf_counter_q[275] : 
                      (N82)? perf_counter_q[339] : 
                      (N83)? perf_counter_q[403] : 
                      (N84)? perf_counter_q[467] : 
                      (N85)? perf_counter_q[531] : 
                      (N86)? perf_counter_q[595] : 
                      (N87)? perf_counter_q[659] : 
                      (N88)? perf_counter_q[723] : 
                      (N89)? perf_counter_q[787] : 1'b0;
  assign data_o[18] = (N76)? perf_counter_q[850] : 
                      (N77)? perf_counter_q[18] : 
                      (N78)? perf_counter_q[82] : 
                      (N79)? perf_counter_q[146] : 
                      (N80)? perf_counter_q[210] : 
                      (N81)? perf_counter_q[274] : 
                      (N82)? perf_counter_q[338] : 
                      (N83)? perf_counter_q[402] : 
                      (N84)? perf_counter_q[466] : 
                      (N85)? perf_counter_q[530] : 
                      (N86)? perf_counter_q[594] : 
                      (N87)? perf_counter_q[658] : 
                      (N88)? perf_counter_q[722] : 
                      (N89)? perf_counter_q[786] : 1'b0;
  assign data_o[17] = (N76)? perf_counter_q[849] : 
                      (N77)? perf_counter_q[17] : 
                      (N78)? perf_counter_q[81] : 
                      (N79)? perf_counter_q[145] : 
                      (N80)? perf_counter_q[209] : 
                      (N81)? perf_counter_q[273] : 
                      (N82)? perf_counter_q[337] : 
                      (N83)? perf_counter_q[401] : 
                      (N84)? perf_counter_q[465] : 
                      (N85)? perf_counter_q[529] : 
                      (N86)? perf_counter_q[593] : 
                      (N87)? perf_counter_q[657] : 
                      (N88)? perf_counter_q[721] : 
                      (N89)? perf_counter_q[785] : 1'b0;
  assign data_o[16] = (N76)? perf_counter_q[848] : 
                      (N77)? perf_counter_q[16] : 
                      (N78)? perf_counter_q[80] : 
                      (N79)? perf_counter_q[144] : 
                      (N80)? perf_counter_q[208] : 
                      (N81)? perf_counter_q[272] : 
                      (N82)? perf_counter_q[336] : 
                      (N83)? perf_counter_q[400] : 
                      (N84)? perf_counter_q[464] : 
                      (N85)? perf_counter_q[528] : 
                      (N86)? perf_counter_q[592] : 
                      (N87)? perf_counter_q[656] : 
                      (N88)? perf_counter_q[720] : 
                      (N89)? perf_counter_q[784] : 1'b0;
  assign data_o[15] = (N76)? perf_counter_q[847] : 
                      (N77)? perf_counter_q[15] : 
                      (N78)? perf_counter_q[79] : 
                      (N79)? perf_counter_q[143] : 
                      (N80)? perf_counter_q[207] : 
                      (N81)? perf_counter_q[271] : 
                      (N82)? perf_counter_q[335] : 
                      (N83)? perf_counter_q[399] : 
                      (N84)? perf_counter_q[463] : 
                      (N85)? perf_counter_q[527] : 
                      (N86)? perf_counter_q[591] : 
                      (N87)? perf_counter_q[655] : 
                      (N88)? perf_counter_q[719] : 
                      (N89)? perf_counter_q[783] : 1'b0;
  assign data_o[14] = (N76)? perf_counter_q[846] : 
                      (N77)? perf_counter_q[14] : 
                      (N78)? perf_counter_q[78] : 
                      (N79)? perf_counter_q[142] : 
                      (N80)? perf_counter_q[206] : 
                      (N81)? perf_counter_q[270] : 
                      (N82)? perf_counter_q[334] : 
                      (N83)? perf_counter_q[398] : 
                      (N84)? perf_counter_q[462] : 
                      (N85)? perf_counter_q[526] : 
                      (N86)? perf_counter_q[590] : 
                      (N87)? perf_counter_q[654] : 
                      (N88)? perf_counter_q[718] : 
                      (N89)? perf_counter_q[782] : 1'b0;
  assign data_o[13] = (N76)? perf_counter_q[845] : 
                      (N77)? perf_counter_q[13] : 
                      (N78)? perf_counter_q[77] : 
                      (N79)? perf_counter_q[141] : 
                      (N80)? perf_counter_q[205] : 
                      (N81)? perf_counter_q[269] : 
                      (N82)? perf_counter_q[333] : 
                      (N83)? perf_counter_q[397] : 
                      (N84)? perf_counter_q[461] : 
                      (N85)? perf_counter_q[525] : 
                      (N86)? perf_counter_q[589] : 
                      (N87)? perf_counter_q[653] : 
                      (N88)? perf_counter_q[717] : 
                      (N89)? perf_counter_q[781] : 1'b0;
  assign data_o[12] = (N76)? perf_counter_q[844] : 
                      (N77)? perf_counter_q[12] : 
                      (N78)? perf_counter_q[76] : 
                      (N79)? perf_counter_q[140] : 
                      (N80)? perf_counter_q[204] : 
                      (N81)? perf_counter_q[268] : 
                      (N82)? perf_counter_q[332] : 
                      (N83)? perf_counter_q[396] : 
                      (N84)? perf_counter_q[460] : 
                      (N85)? perf_counter_q[524] : 
                      (N86)? perf_counter_q[588] : 
                      (N87)? perf_counter_q[652] : 
                      (N88)? perf_counter_q[716] : 
                      (N89)? perf_counter_q[780] : 1'b0;
  assign data_o[11] = (N76)? perf_counter_q[843] : 
                      (N77)? perf_counter_q[11] : 
                      (N78)? perf_counter_q[75] : 
                      (N79)? perf_counter_q[139] : 
                      (N80)? perf_counter_q[203] : 
                      (N81)? perf_counter_q[267] : 
                      (N82)? perf_counter_q[331] : 
                      (N83)? perf_counter_q[395] : 
                      (N84)? perf_counter_q[459] : 
                      (N85)? perf_counter_q[523] : 
                      (N86)? perf_counter_q[587] : 
                      (N87)? perf_counter_q[651] : 
                      (N88)? perf_counter_q[715] : 
                      (N89)? perf_counter_q[779] : 1'b0;
  assign data_o[10] = (N76)? perf_counter_q[842] : 
                      (N77)? perf_counter_q[10] : 
                      (N78)? perf_counter_q[74] : 
                      (N79)? perf_counter_q[138] : 
                      (N80)? perf_counter_q[202] : 
                      (N81)? perf_counter_q[266] : 
                      (N82)? perf_counter_q[330] : 
                      (N83)? perf_counter_q[394] : 
                      (N84)? perf_counter_q[458] : 
                      (N85)? perf_counter_q[522] : 
                      (N86)? perf_counter_q[586] : 
                      (N87)? perf_counter_q[650] : 
                      (N88)? perf_counter_q[714] : 
                      (N89)? perf_counter_q[778] : 1'b0;
  assign data_o[9] = (N76)? perf_counter_q[841] : 
                     (N77)? perf_counter_q[9] : 
                     (N78)? perf_counter_q[73] : 
                     (N79)? perf_counter_q[137] : 
                     (N80)? perf_counter_q[201] : 
                     (N81)? perf_counter_q[265] : 
                     (N82)? perf_counter_q[329] : 
                     (N83)? perf_counter_q[393] : 
                     (N84)? perf_counter_q[457] : 
                     (N85)? perf_counter_q[521] : 
                     (N86)? perf_counter_q[585] : 
                     (N87)? perf_counter_q[649] : 
                     (N88)? perf_counter_q[713] : 
                     (N89)? perf_counter_q[777] : 1'b0;
  assign data_o[8] = (N76)? perf_counter_q[840] : 
                     (N77)? perf_counter_q[8] : 
                     (N78)? perf_counter_q[72] : 
                     (N79)? perf_counter_q[136] : 
                     (N80)? perf_counter_q[200] : 
                     (N81)? perf_counter_q[264] : 
                     (N82)? perf_counter_q[328] : 
                     (N83)? perf_counter_q[392] : 
                     (N84)? perf_counter_q[456] : 
                     (N85)? perf_counter_q[520] : 
                     (N86)? perf_counter_q[584] : 
                     (N87)? perf_counter_q[648] : 
                     (N88)? perf_counter_q[712] : 
                     (N89)? perf_counter_q[776] : 1'b0;
  assign data_o[7] = (N76)? perf_counter_q[839] : 
                     (N77)? perf_counter_q[7] : 
                     (N78)? perf_counter_q[71] : 
                     (N79)? perf_counter_q[135] : 
                     (N80)? perf_counter_q[199] : 
                     (N81)? perf_counter_q[263] : 
                     (N82)? perf_counter_q[327] : 
                     (N83)? perf_counter_q[391] : 
                     (N84)? perf_counter_q[455] : 
                     (N85)? perf_counter_q[519] : 
                     (N86)? perf_counter_q[583] : 
                     (N87)? perf_counter_q[647] : 
                     (N88)? perf_counter_q[711] : 
                     (N89)? perf_counter_q[775] : 1'b0;
  assign data_o[6] = (N76)? perf_counter_q[838] : 
                     (N77)? perf_counter_q[6] : 
                     (N78)? perf_counter_q[70] : 
                     (N79)? perf_counter_q[134] : 
                     (N80)? perf_counter_q[198] : 
                     (N81)? perf_counter_q[262] : 
                     (N82)? perf_counter_q[326] : 
                     (N83)? perf_counter_q[390] : 
                     (N84)? perf_counter_q[454] : 
                     (N85)? perf_counter_q[518] : 
                     (N86)? perf_counter_q[582] : 
                     (N87)? perf_counter_q[646] : 
                     (N88)? perf_counter_q[710] : 
                     (N89)? perf_counter_q[774] : 1'b0;
  assign data_o[5] = (N76)? perf_counter_q[837] : 
                     (N77)? perf_counter_q[5] : 
                     (N78)? perf_counter_q[69] : 
                     (N79)? perf_counter_q[133] : 
                     (N80)? perf_counter_q[197] : 
                     (N81)? perf_counter_q[261] : 
                     (N82)? perf_counter_q[325] : 
                     (N83)? perf_counter_q[389] : 
                     (N84)? perf_counter_q[453] : 
                     (N85)? perf_counter_q[517] : 
                     (N86)? perf_counter_q[581] : 
                     (N87)? perf_counter_q[645] : 
                     (N88)? perf_counter_q[709] : 
                     (N89)? perf_counter_q[773] : 1'b0;
  assign data_o[4] = (N76)? perf_counter_q[836] : 
                     (N77)? perf_counter_q[4] : 
                     (N78)? perf_counter_q[68] : 
                     (N79)? perf_counter_q[132] : 
                     (N80)? perf_counter_q[196] : 
                     (N81)? perf_counter_q[260] : 
                     (N82)? perf_counter_q[324] : 
                     (N83)? perf_counter_q[388] : 
                     (N84)? perf_counter_q[452] : 
                     (N85)? perf_counter_q[516] : 
                     (N86)? perf_counter_q[580] : 
                     (N87)? perf_counter_q[644] : 
                     (N88)? perf_counter_q[708] : 
                     (N89)? perf_counter_q[772] : 1'b0;
  assign data_o[3] = (N76)? perf_counter_q[835] : 
                     (N77)? perf_counter_q[3] : 
                     (N78)? perf_counter_q[67] : 
                     (N79)? perf_counter_q[131] : 
                     (N80)? perf_counter_q[195] : 
                     (N81)? perf_counter_q[259] : 
                     (N82)? perf_counter_q[323] : 
                     (N83)? perf_counter_q[387] : 
                     (N84)? perf_counter_q[451] : 
                     (N85)? perf_counter_q[515] : 
                     (N86)? perf_counter_q[579] : 
                     (N87)? perf_counter_q[643] : 
                     (N88)? perf_counter_q[707] : 
                     (N89)? perf_counter_q[771] : 1'b0;
  assign data_o[2] = (N76)? perf_counter_q[834] : 
                     (N77)? perf_counter_q[2] : 
                     (N78)? perf_counter_q[66] : 
                     (N79)? perf_counter_q[130] : 
                     (N80)? perf_counter_q[194] : 
                     (N81)? perf_counter_q[258] : 
                     (N82)? perf_counter_q[322] : 
                     (N83)? perf_counter_q[386] : 
                     (N84)? perf_counter_q[450] : 
                     (N85)? perf_counter_q[514] : 
                     (N86)? perf_counter_q[578] : 
                     (N87)? perf_counter_q[642] : 
                     (N88)? perf_counter_q[706] : 
                     (N89)? perf_counter_q[770] : 1'b0;
  assign data_o[1] = (N76)? perf_counter_q[833] : 
                     (N77)? perf_counter_q[1] : 
                     (N78)? perf_counter_q[65] : 
                     (N79)? perf_counter_q[129] : 
                     (N80)? perf_counter_q[193] : 
                     (N81)? perf_counter_q[257] : 
                     (N82)? perf_counter_q[321] : 
                     (N83)? perf_counter_q[385] : 
                     (N84)? perf_counter_q[449] : 
                     (N85)? perf_counter_q[513] : 
                     (N86)? perf_counter_q[577] : 
                     (N87)? perf_counter_q[641] : 
                     (N88)? perf_counter_q[705] : 
                     (N89)? perf_counter_q[769] : 1'b0;
  assign data_o[0] = (N76)? perf_counter_q[832] : 
                     (N77)? perf_counter_q[0] : 
                     (N78)? perf_counter_q[64] : 
                     (N79)? perf_counter_q[128] : 
                     (N80)? perf_counter_q[192] : 
                     (N81)? perf_counter_q[256] : 
                     (N82)? perf_counter_q[320] : 
                     (N83)? perf_counter_q[384] : 
                     (N84)? perf_counter_q[448] : 
                     (N85)? perf_counter_q[512] : 
                     (N86)? perf_counter_q[576] : 
                     (N87)? perf_counter_q[640] : 
                     (N88)? perf_counter_q[704] : 
                     (N89)? perf_counter_q[768] : 1'b0;
  assign N90 = ~debug_mode_i;
  assign N91 = N90;
  assign N92 = ~l1_icache_miss_i;
  assign N221 = ~l1_dcache_miss_i;
  assign N350 = ~itlb_miss_i;
  assign N479 = ~dtlb_miss_i;
  assign N608 = ~commit_ack_i[0];
  assign N609 = N91 & commit_ack_i[0];
  assign N994 = N4123 & N4099;
  assign N4123 = N4060 & N4092;
  assign N995 = ~N994;
  assign N1124 = N4079 & N4086;
  assign N1125 = ~N1124;
  assign N1574 = ~ex_i[0];
  assign N1703 = ~eret_i;
  assign N1832 = resolved_branch_i[3] & resolved_branch_i[5];
  assign N1833 = ~N1832;
  assign N1962 = ~sb_full_i;
  assign N2091 = ~if_empty_i;
  assign N3130 = ~we_i;
  assign N3145 = ~N3131;
  assign N3210 = ~N3132;
  assign N3275 = ~N3133;
  assign N3340 = ~N3134;
  assign N3405 = ~N3135;
  assign N3470 = ~N3136;
  assign N3535 = ~N3137;
  assign N3600 = ~N3138;
  assign N3665 = ~N3139;
  assign N3730 = ~N3140;
  assign N3795 = ~N3141;
  assign N3860 = ~N3142;
  assign N3925 = ~N3143;
  assign N3990 = ~N3144;
  assign N4055 = ~rst_ni;

endmodule