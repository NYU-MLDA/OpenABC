module bsg_mem_1r1w_synth_width_p537_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [536:0] w_data_i;
  input [0:0] r_addr_i;
  output [536:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [536:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18;
  reg [1073:0] mem;
  assign r_data_o[536] = (N3)? mem[536] :
                         (N0)? mem[1073] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[535] = (N3)? mem[535] :
                         (N0)? mem[1072] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] :
                         (N0)? mem[1071] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] :
                         (N0)? mem[1070] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] :
                         (N0)? mem[1069] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] :
                         (N0)? mem[1068] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] :
                         (N0)? mem[1067] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] :
                         (N0)? mem[1066] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] :
                         (N0)? mem[1065] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] :
                         (N0)? mem[1064] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] :
                         (N0)? mem[1063] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] :
                         (N0)? mem[1062] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] :
                         (N0)? mem[1061] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] :
                         (N0)? mem[1060] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] :
                         (N0)? mem[1059] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] :
                         (N0)? mem[1058] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] :
                         (N0)? mem[1057] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] :
                         (N0)? mem[1056] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] :
                         (N0)? mem[1055] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] :
                         (N0)? mem[1054] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] :
                         (N0)? mem[1053] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] :
                         (N0)? mem[1052] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] :
                         (N0)? mem[1051] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] :
                         (N0)? mem[1050] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] :
                         (N0)? mem[1049] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] :
                         (N0)? mem[1048] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] :
                         (N0)? mem[1047] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] :
                         (N0)? mem[1046] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] :
                         (N0)? mem[1045] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] :
                         (N0)? mem[1044] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] :
                         (N0)? mem[1043] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] :
                         (N0)? mem[1042] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] :
                         (N0)? mem[1041] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] :
                         (N0)? mem[1040] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] :
                         (N0)? mem[1039] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] :
                         (N0)? mem[1038] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] :
                         (N0)? mem[1037] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] :
                         (N0)? mem[1036] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] :
                         (N0)? mem[1035] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] :
                         (N0)? mem[1034] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] :
                         (N0)? mem[1033] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] :
                         (N0)? mem[1032] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] :
                         (N0)? mem[1031] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] :
                         (N0)? mem[1030] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] :
                         (N0)? mem[1029] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] :
                         (N0)? mem[1028] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] :
                         (N0)? mem[1027] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] :
                         (N0)? mem[1026] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] :
                         (N0)? mem[1025] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] :
                         (N0)? mem[1024] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] :
                         (N0)? mem[1023] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] :
                         (N0)? mem[1022] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] :
                         (N0)? mem[1021] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] :
                         (N0)? mem[1020] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] :
                         (N0)? mem[1019] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] :
                         (N0)? mem[1018] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] :
                         (N0)? mem[1017] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] :
                         (N0)? mem[1016] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] :
                         (N0)? mem[1015] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] :
                         (N0)? mem[1014] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] :
                         (N0)? mem[1013] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] :
                         (N0)? mem[1012] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] :
                         (N0)? mem[1011] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] :
                         (N0)? mem[1010] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] :
                         (N0)? mem[1009] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] :
                         (N0)? mem[1008] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] :
                         (N0)? mem[1007] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] :
                         (N0)? mem[1006] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] :
                         (N0)? mem[1005] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] :
                         (N0)? mem[1004] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] :
                         (N0)? mem[1003] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] :
                         (N0)? mem[1002] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] :
                         (N0)? mem[1001] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] :
                         (N0)? mem[1000] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] :
                         (N0)? mem[999] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] :
                         (N0)? mem[998] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] :
                         (N0)? mem[997] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] :
                         (N0)? mem[996] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] :
                         (N0)? mem[995] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] :
                         (N0)? mem[994] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] :
                         (N0)? mem[993] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] :
                         (N0)? mem[992] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] :
                         (N0)? mem[991] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] :
                         (N0)? mem[990] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] :
                         (N0)? mem[989] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] :
                         (N0)? mem[988] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] :
                         (N0)? mem[987] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] :
                         (N0)? mem[986] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] :
                         (N0)? mem[985] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] :
                         (N0)? mem[984] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] :
                         (N0)? mem[983] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] :
                         (N0)? mem[982] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] :
                         (N0)? mem[981] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] :
                         (N0)? mem[980] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] :
                         (N0)? mem[979] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] :
                         (N0)? mem[978] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] :
                         (N0)? mem[977] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] :
                         (N0)? mem[976] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] :
                         (N0)? mem[975] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] :
                         (N0)? mem[974] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] :
                         (N0)? mem[973] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] :
                         (N0)? mem[972] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] :
                         (N0)? mem[971] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] :
                         (N0)? mem[970] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] :
                         (N0)? mem[969] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] :
                         (N0)? mem[968] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] :
                         (N0)? mem[967] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] :
                         (N0)? mem[966] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] :
                         (N0)? mem[965] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] :
                         (N0)? mem[964] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] :
                         (N0)? mem[963] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] :
                         (N0)? mem[962] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] :
                         (N0)? mem[961] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] :
                         (N0)? mem[960] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] :
                         (N0)? mem[959] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] :
                         (N0)? mem[958] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] :
                         (N0)? mem[957] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] :
                         (N0)? mem[956] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] :
                         (N0)? mem[955] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] :
                         (N0)? mem[954] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] :
                         (N0)? mem[953] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] :
                         (N0)? mem[952] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] :
                         (N0)? mem[951] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] :
                         (N0)? mem[950] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] :
                         (N0)? mem[949] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] :
                         (N0)? mem[948] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] :
                         (N0)? mem[947] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] :
                         (N0)? mem[946] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] :
                         (N0)? mem[945] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] :
                         (N0)? mem[944] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] :
                         (N0)? mem[943] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] :
                         (N0)? mem[942] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] :
                         (N0)? mem[941] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] :
                         (N0)? mem[940] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] :
                         (N0)? mem[939] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] :
                         (N0)? mem[938] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] :
                         (N0)? mem[937] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] :
                         (N0)? mem[936] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] :
                         (N0)? mem[935] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] :
                         (N0)? mem[934] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] :
                         (N0)? mem[933] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] :
                         (N0)? mem[932] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] :
                         (N0)? mem[931] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] :
                         (N0)? mem[930] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] :
                         (N0)? mem[929] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] :
                         (N0)? mem[928] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] :
                         (N0)? mem[927] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] :
                         (N0)? mem[926] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] :
                         (N0)? mem[925] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] :
                         (N0)? mem[924] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] :
                         (N0)? mem[923] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] :
                         (N0)? mem[922] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] :
                         (N0)? mem[921] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] :
                         (N0)? mem[920] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] :
                         (N0)? mem[919] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] :
                         (N0)? mem[918] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] :
                         (N0)? mem[917] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] :
                         (N0)? mem[916] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] :
                         (N0)? mem[915] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] :
                         (N0)? mem[914] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] :
                         (N0)? mem[913] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] :
                         (N0)? mem[912] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] :
                         (N0)? mem[911] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] :
                         (N0)? mem[910] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] :
                         (N0)? mem[909] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] :
                         (N0)? mem[908] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] :
                         (N0)? mem[907] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] :
                         (N0)? mem[906] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] :
                         (N0)? mem[905] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] :
                         (N0)? mem[904] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] :
                         (N0)? mem[903] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] :
                         (N0)? mem[902] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] :
                         (N0)? mem[901] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] :
                         (N0)? mem[900] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] :
                         (N0)? mem[899] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] :
                         (N0)? mem[898] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] :
                         (N0)? mem[897] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] :
                         (N0)? mem[896] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] :
                         (N0)? mem[895] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] :
                         (N0)? mem[894] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] :
                         (N0)? mem[893] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] :
                         (N0)? mem[892] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] :
                         (N0)? mem[891] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] :
                         (N0)? mem[890] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] :
                         (N0)? mem[889] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] :
                         (N0)? mem[888] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] :
                         (N0)? mem[887] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] :
                         (N0)? mem[886] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] :
                         (N0)? mem[885] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] :
                         (N0)? mem[884] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] :
                         (N0)? mem[883] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] :
                         (N0)? mem[882] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] :
                         (N0)? mem[881] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] :
                         (N0)? mem[880] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] :
                         (N0)? mem[879] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] :
                         (N0)? mem[878] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] :
                         (N0)? mem[877] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] :
                         (N0)? mem[876] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] :
                         (N0)? mem[875] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] :
                         (N0)? mem[874] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] :
                         (N0)? mem[873] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] :
                         (N0)? mem[872] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] :
                         (N0)? mem[871] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] :
                         (N0)? mem[870] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] :
                         (N0)? mem[869] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] :
                         (N0)? mem[868] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] :
                         (N0)? mem[867] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] :
                         (N0)? mem[866] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] :
                         (N0)? mem[865] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] :
                         (N0)? mem[864] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] :
                         (N0)? mem[863] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] :
                         (N0)? mem[862] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] :
                         (N0)? mem[861] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] :
                         (N0)? mem[860] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] :
                         (N0)? mem[859] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] :
                         (N0)? mem[858] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] :
                         (N0)? mem[857] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] :
                         (N0)? mem[856] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] :
                         (N0)? mem[855] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] :
                         (N0)? mem[854] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] :
                         (N0)? mem[853] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] :
                         (N0)? mem[852] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] :
                         (N0)? mem[851] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] :
                         (N0)? mem[850] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] :
                         (N0)? mem[849] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] :
                         (N0)? mem[848] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] :
                         (N0)? mem[847] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] :
                         (N0)? mem[846] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] :
                         (N0)? mem[845] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] :
                         (N0)? mem[844] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] :
                         (N0)? mem[843] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] :
                         (N0)? mem[842] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] :
                         (N0)? mem[841] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] :
                         (N0)? mem[840] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] :
                         (N0)? mem[839] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] :
                         (N0)? mem[838] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] :
                         (N0)? mem[837] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] :
                         (N0)? mem[836] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] :
                         (N0)? mem[835] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] :
                         (N0)? mem[834] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] :
                         (N0)? mem[833] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] :
                         (N0)? mem[832] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] :
                         (N0)? mem[831] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] :
                         (N0)? mem[830] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] :
                         (N0)? mem[829] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] :
                         (N0)? mem[828] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] :
                         (N0)? mem[827] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] :
                         (N0)? mem[826] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] :
                         (N0)? mem[825] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] :
                         (N0)? mem[824] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] :
                         (N0)? mem[823] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] :
                         (N0)? mem[822] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] :
                         (N0)? mem[821] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] :
                         (N0)? mem[820] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] :
                         (N0)? mem[819] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] :
                         (N0)? mem[818] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] :
                         (N0)? mem[817] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] :
                         (N0)? mem[816] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] :
                         (N0)? mem[815] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] :
                         (N0)? mem[814] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] :
                         (N0)? mem[813] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] :
                         (N0)? mem[812] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] :
                         (N0)? mem[811] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] :
                         (N0)? mem[810] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] :
                         (N0)? mem[809] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] :
                         (N0)? mem[808] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] :
                         (N0)? mem[807] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] :
                         (N0)? mem[806] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] :
                         (N0)? mem[805] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] :
                         (N0)? mem[804] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] :
                         (N0)? mem[803] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] :
                         (N0)? mem[802] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] :
                         (N0)? mem[801] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] :
                         (N0)? mem[800] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] :
                         (N0)? mem[799] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] :
                         (N0)? mem[798] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] :
                         (N0)? mem[797] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] :
                         (N0)? mem[796] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] :
                         (N0)? mem[795] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] :
                         (N0)? mem[794] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] :
                         (N0)? mem[793] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] :
                         (N0)? mem[792] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] :
                         (N0)? mem[791] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] :
                         (N0)? mem[790] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] :
                         (N0)? mem[789] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] :
                         (N0)? mem[788] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] :
                         (N0)? mem[787] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] :
                         (N0)? mem[786] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] :
                         (N0)? mem[785] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] :
                         (N0)? mem[784] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] :
                         (N0)? mem[783] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] :
                         (N0)? mem[782] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] :
                         (N0)? mem[781] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] :
                         (N0)? mem[780] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] :
                         (N0)? mem[779] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] :
                         (N0)? mem[778] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] :
                         (N0)? mem[777] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] :
                         (N0)? mem[776] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] :
                         (N0)? mem[775] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] :
                         (N0)? mem[774] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] :
                         (N0)? mem[773] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] :
                         (N0)? mem[772] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] :
                         (N0)? mem[771] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] :
                         (N0)? mem[770] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] :
                         (N0)? mem[769] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] :
                         (N0)? mem[768] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] :
                         (N0)? mem[767] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] :
                         (N0)? mem[766] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] :
                         (N0)? mem[765] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] :
                         (N0)? mem[764] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] :
                         (N0)? mem[763] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] :
                         (N0)? mem[762] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] :
                         (N0)? mem[761] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] :
                         (N0)? mem[760] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] :
                         (N0)? mem[759] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] :
                         (N0)? mem[758] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] :
                         (N0)? mem[757] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] :
                         (N0)? mem[756] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] :
                         (N0)? mem[755] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] :
                         (N0)? mem[754] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] :
                         (N0)? mem[753] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] :
                         (N0)? mem[752] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] :
                         (N0)? mem[751] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] :
                         (N0)? mem[750] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] :
                         (N0)? mem[749] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] :
                         (N0)? mem[748] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] :
                         (N0)? mem[747] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] :
                         (N0)? mem[746] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] :
                         (N0)? mem[745] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] :
                         (N0)? mem[744] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] :
                         (N0)? mem[743] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] :
                         (N0)? mem[742] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] :
                         (N0)? mem[741] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] :
                         (N0)? mem[740] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] :
                         (N0)? mem[739] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] :
                         (N0)? mem[738] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] :
                         (N0)? mem[737] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] :
                         (N0)? mem[736] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] :
                         (N0)? mem[735] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] :
                         (N0)? mem[734] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] :
                         (N0)? mem[733] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] :
                         (N0)? mem[732] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] :
                         (N0)? mem[731] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] :
                         (N0)? mem[730] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] :
                         (N0)? mem[729] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] :
                         (N0)? mem[728] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] :
                         (N0)? mem[727] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] :
                         (N0)? mem[726] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] :
                         (N0)? mem[725] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] :
                         (N0)? mem[724] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] :
                         (N0)? mem[723] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] :
                         (N0)? mem[722] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] :
                         (N0)? mem[721] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] :
                         (N0)? mem[720] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] :
                         (N0)? mem[719] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] :
                         (N0)? mem[718] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] :
                         (N0)? mem[717] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] :
                         (N0)? mem[716] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] :
                         (N0)? mem[715] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] :
                         (N0)? mem[714] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] :
                         (N0)? mem[713] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] :
                         (N0)? mem[712] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] :
                         (N0)? mem[711] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] :
                         (N0)? mem[710] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] :
                         (N0)? mem[709] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] :
                         (N0)? mem[708] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] :
                         (N0)? mem[707] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] :
                         (N0)? mem[706] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] :
                         (N0)? mem[705] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] :
                         (N0)? mem[704] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] :
                         (N0)? mem[703] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] :
                         (N0)? mem[702] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] :
                         (N0)? mem[701] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] :
                         (N0)? mem[700] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] :
                         (N0)? mem[699] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] :
                         (N0)? mem[698] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] :
                         (N0)? mem[697] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] :
                         (N0)? mem[696] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] :
                         (N0)? mem[695] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] :
                         (N0)? mem[694] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] :
                         (N0)? mem[693] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] :
                         (N0)? mem[692] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] :
                         (N0)? mem[691] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] :
                         (N0)? mem[690] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] :
                         (N0)? mem[689] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] :
                         (N0)? mem[688] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] :
                         (N0)? mem[687] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] :
                         (N0)? mem[686] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] :
                         (N0)? mem[685] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] :
                         (N0)? mem[684] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] :
                         (N0)? mem[683] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] :
                         (N0)? mem[682] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] :
                         (N0)? mem[681] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] :
                         (N0)? mem[680] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] :
                         (N0)? mem[679] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] :
                         (N0)? mem[678] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] :
                         (N0)? mem[677] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] :
                         (N0)? mem[676] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] :
                         (N0)? mem[675] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] :
                         (N0)? mem[674] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] :
                         (N0)? mem[673] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] :
                         (N0)? mem[672] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] :
                         (N0)? mem[671] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] :
                         (N0)? mem[670] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] :
                         (N0)? mem[669] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] :
                         (N0)? mem[668] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] :
                         (N0)? mem[667] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] :
                         (N0)? mem[666] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] :
                         (N0)? mem[665] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] :
                         (N0)? mem[664] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] :
                         (N0)? mem[663] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] :
                         (N0)? mem[662] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] :
                         (N0)? mem[661] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] :
                         (N0)? mem[660] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] :
                         (N0)? mem[659] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] :
                         (N0)? mem[658] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] :
                         (N0)? mem[657] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] :
                         (N0)? mem[656] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] :
                         (N0)? mem[655] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] :
                         (N0)? mem[654] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] :
                         (N0)? mem[653] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] :
                         (N0)? mem[652] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] :
                         (N0)? mem[651] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] :
                         (N0)? mem[650] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] :
                         (N0)? mem[649] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] :
                         (N0)? mem[648] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] :
                         (N0)? mem[647] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] :
                         (N0)? mem[646] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] :
                         (N0)? mem[645] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] :
                         (N0)? mem[644] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] :
                         (N0)? mem[643] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] :
                         (N0)? mem[642] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] :
                         (N0)? mem[641] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] :
                         (N0)? mem[640] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] :
                         (N0)? mem[639] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] :
                         (N0)? mem[638] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] :
                         (N0)? mem[637] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] :
                        (N0)? mem[636] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] :
                        (N0)? mem[635] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] :
                        (N0)? mem[634] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] :
                        (N0)? mem[633] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] :
                        (N0)? mem[632] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] :
                        (N0)? mem[631] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] :
                        (N0)? mem[630] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] :
                        (N0)? mem[629] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] :
                        (N0)? mem[628] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] :
                        (N0)? mem[627] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] :
                        (N0)? mem[626] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] :
                        (N0)? mem[625] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] :
                        (N0)? mem[624] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] :
                        (N0)? mem[623] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] :
                        (N0)? mem[622] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] :
                        (N0)? mem[621] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] :
                        (N0)? mem[620] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] :
                        (N0)? mem[619] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] :
                        (N0)? mem[618] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] :
                        (N0)? mem[617] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] :
                        (N0)? mem[616] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] :
                        (N0)? mem[615] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] :
                        (N0)? mem[614] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] :
                        (N0)? mem[613] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] :
                        (N0)? mem[612] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] :
                        (N0)? mem[611] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] :
                        (N0)? mem[610] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] :
                        (N0)? mem[609] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] :
                        (N0)? mem[608] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] :
                        (N0)? mem[607] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] :
                        (N0)? mem[606] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] :
                        (N0)? mem[605] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] :
                        (N0)? mem[604] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] :
                        (N0)? mem[603] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] :
                        (N0)? mem[602] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] :
                        (N0)? mem[601] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] :
                        (N0)? mem[600] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] :
                        (N0)? mem[599] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] :
                        (N0)? mem[598] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] :
                        (N0)? mem[597] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] :
                        (N0)? mem[596] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] :
                        (N0)? mem[595] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] :
                        (N0)? mem[594] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] :
                        (N0)? mem[593] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] :
                        (N0)? mem[592] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] :
                        (N0)? mem[591] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] :
                        (N0)? mem[590] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] :
                        (N0)? mem[589] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] :
                        (N0)? mem[588] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] :
                        (N0)? mem[587] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] :
                        (N0)? mem[586] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] :
                        (N0)? mem[585] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] :
                        (N0)? mem[584] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] :
                        (N0)? mem[583] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] :
                        (N0)? mem[582] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] :
                        (N0)? mem[581] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] :
                        (N0)? mem[580] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] :
                        (N0)? mem[579] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] :
                        (N0)? mem[578] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] :
                        (N0)? mem[577] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] :
                        (N0)? mem[576] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] :
                        (N0)? mem[575] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] :
                        (N0)? mem[574] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] :
                        (N0)? mem[573] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] :
                        (N0)? mem[572] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] :
                        (N0)? mem[571] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] :
                        (N0)? mem[570] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] :
                        (N0)? mem[569] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] :
                        (N0)? mem[568] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] :
                        (N0)? mem[567] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] :
                        (N0)? mem[566] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] :
                        (N0)? mem[565] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] :
                        (N0)? mem[564] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] :
                        (N0)? mem[563] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] :
                        (N0)? mem[562] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] :
                        (N0)? mem[561] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] :
                        (N0)? mem[560] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] :
                        (N0)? mem[559] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] :
                        (N0)? mem[558] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] :
                        (N0)? mem[557] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] :
                        (N0)? mem[556] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] :
                        (N0)? mem[555] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] :
                        (N0)? mem[554] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] :
                        (N0)? mem[553] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] :
                        (N0)? mem[552] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] :
                        (N0)? mem[551] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] :
                        (N0)? mem[550] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] :
                        (N0)? mem[549] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] :
                        (N0)? mem[548] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] :
                        (N0)? mem[547] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] :
                       (N0)? mem[546] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] :
                       (N0)? mem[545] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] :
                       (N0)? mem[544] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] :
                       (N0)? mem[543] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] :
                       (N0)? mem[542] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] :
                       (N0)? mem[541] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] :
                       (N0)? mem[540] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] :
                       (N0)? mem[539] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] :
                       (N0)? mem[538] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] :
                       (N0)? mem[537] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5 } :
                                                                       (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N13) begin
      { mem[1073:975], mem[537:537] } <= { w_data_i[536:438], w_data_i[0:0] };
    end
    if(N14) begin
      { mem[974:876], mem[538:538] } <= { w_data_i[437:339], w_data_i[1:1] };
    end
    if(N15) begin
      { mem[875:777], mem[539:539] } <= { w_data_i[338:240], w_data_i[2:2] };
    end
    if(N16) begin
      { mem[776:678], mem[540:540] } <= { w_data_i[239:141], w_data_i[3:3] };
    end
    if(N17) begin
      { mem[677:579], mem[541:541] } <= { w_data_i[140:42], w_data_i[4:4] };
    end
    if(N18) begin
      { mem[578:542] } <= { w_data_i[41:5] };
    end
    if(N7) begin
      { mem[536:438], mem[0:0] } <= { w_data_i[536:438], w_data_i[0:0] };
    end
    if(N8) begin
      { mem[437:339], mem[1:1] } <= { w_data_i[437:339], w_data_i[1:1] };
    end
    if(N9) begin
      { mem[338:240], mem[2:2] } <= { w_data_i[338:240], w_data_i[2:2] };
    end
    if(N10) begin
      { mem[239:141], mem[3:3] } <= { w_data_i[239:141], w_data_i[3:3] };
    end
    if(N11) begin
      { mem[140:42], mem[4:4] } <= { w_data_i[140:42], w_data_i[4:4] };
    end
    if(N12) begin
      { mem[41:5] } <= { w_data_i[41:5] };
    end
  end


endmodule