module ariane_regfile_64_2_00000002_1
(
  clk_i,
  rst_ni,
  test_en_i,
  raddr_i,
  rdata_o,
  waddr_i,
  wdata_i,
  we_i
);

  input [9:0] raddr_i;
  output [127:0] rdata_o;
  input [9:0] waddr_i;
  input [127:0] wdata_i;
  input [1:0] we_i;
  input clk_i;
  input rst_ni;
  input test_en_i;
  wire [127:0] rdata_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,we_dec_1__31_,we_dec_1__30_,we_dec_1__29_,we_dec_1__28_,
  we_dec_1__27_,we_dec_1__26_,we_dec_1__25_,we_dec_1__24_,we_dec_1__23_,we_dec_1__22_,
  we_dec_1__21_,we_dec_1__20_,we_dec_1__19_,we_dec_1__18_,we_dec_1__17_,we_dec_1__16_,
  we_dec_1__15_,we_dec_1__14_,we_dec_1__13_,we_dec_1__12_,we_dec_1__11_,
  we_dec_1__10_,we_dec_1__9_,we_dec_1__8_,we_dec_1__7_,we_dec_1__6_,we_dec_1__5_,
  we_dec_1__4_,we_dec_1__3_,we_dec_1__2_,we_dec_1__1_,we_dec_0__31_,we_dec_0__30_,
  we_dec_0__29_,we_dec_0__28_,we_dec_0__27_,we_dec_0__26_,we_dec_0__25_,we_dec_0__24_,
  we_dec_0__23_,we_dec_0__22_,we_dec_0__21_,we_dec_0__20_,we_dec_0__19_,we_dec_0__18_,
  we_dec_0__17_,we_dec_0__16_,we_dec_0__15_,we_dec_0__14_,we_dec_0__13_,we_dec_0__12_,
  we_dec_0__11_,we_dec_0__10_,we_dec_0__9_,we_dec_0__8_,we_dec_0__7_,we_dec_0__6_,
  we_dec_0__5_,we_dec_0__4_,we_dec_0__3_,we_dec_0__2_,we_dec_0__1_,N153,N154,N155,
  N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,
  N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,
  N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,
  N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,
  N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,
  N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,
  N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,
  N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,
  N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,
  N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,
  N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,
  N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,
  N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,
  N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,
  N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,
  N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,
  N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,
  N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,
  N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,
  N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,
  N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,
  N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,
  N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,
  N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,
  N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,
  N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,
  N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,
  N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,
  N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,
  N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,
  N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,
  N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,
  N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,
  N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,
  N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,
  N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,
  N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,
  N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
  N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,
  N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,
  N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,
  N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,
  N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,
  N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,
  N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,
  N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,
  N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,
  N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,
  N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,
  N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,
  N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,
  N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,
  N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,
  N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,
  N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,
  N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,
  N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,
  N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,
  N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,
  N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,
  N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,
  N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,
  N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,
  N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,
  N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,
  N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,
  N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,
  N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,
  N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,
  N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,
  N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,
  N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,
  N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,
  N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,
  N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,
  N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,
  N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,
  N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,
  N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,
  N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,
  N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,
  N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,
  N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,
  N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,
  N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,
  N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,
  N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,
  N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,
  N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
  N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,
  N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,
  N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,
  N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,
  N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,
  N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,
  N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,
  N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,
  N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,
  N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,
  N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,
  N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,
  N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,
  N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,
  N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,
  N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,
  N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,
  N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,
  N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,
  N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,
  N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,
  N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,
  N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,
  N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,
  N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,
  N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,
  N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,
  N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,
  N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,
  N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,
  N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,
  N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,
  N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,
  N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,
  N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,
  N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,
  N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,
  N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,
  N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,
  N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,
  N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,
  N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,
  N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,
  N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,
  N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,
  N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,
  N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,
  N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,
  N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,
  N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
  N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,
  N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,
  N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,
  N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,
  N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,
  N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,
  N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,
  N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,
  N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,
  N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,
  N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,
  N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,
  N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,
  N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,
  N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,
  N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,
  N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,
  N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,
  N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,
  N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,
  N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,
  N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,
  N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,
  N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,
  N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,
  N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,
  N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,
  N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,
  N2523,N2524,N2525;
  reg [2047:0] mem;

  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2047] <= 1'b0;
    end else if(N2137) begin
      mem[2047] <= N2201;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2046] <= 1'b0;
    end else if(N2137) begin
      mem[2046] <= N2200;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2045] <= 1'b0;
    end else if(N2137) begin
      mem[2045] <= N2199;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2044] <= 1'b0;
    end else if(N2137) begin
      mem[2044] <= N2198;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2043] <= 1'b0;
    end else if(N2137) begin
      mem[2043] <= N2197;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2042] <= 1'b0;
    end else if(N2137) begin
      mem[2042] <= N2196;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2041] <= 1'b0;
    end else if(N2137) begin
      mem[2041] <= N2195;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2040] <= 1'b0;
    end else if(N2137) begin
      mem[2040] <= N2194;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2039] <= 1'b0;
    end else if(N2137) begin
      mem[2039] <= N2193;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2038] <= 1'b0;
    end else if(N2137) begin
      mem[2038] <= N2192;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2037] <= 1'b0;
    end else if(N2137) begin
      mem[2037] <= N2191;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2036] <= 1'b0;
    end else if(N2137) begin
      mem[2036] <= N2190;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2035] <= 1'b0;
    end else if(N2137) begin
      mem[2035] <= N2189;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2034] <= 1'b0;
    end else if(N2137) begin
      mem[2034] <= N2188;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2033] <= 1'b0;
    end else if(N2137) begin
      mem[2033] <= N2187;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2032] <= 1'b0;
    end else if(N2137) begin
      mem[2032] <= N2186;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2031] <= 1'b0;
    end else if(N2137) begin
      mem[2031] <= N2185;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2030] <= 1'b0;
    end else if(N2137) begin
      mem[2030] <= N2184;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2029] <= 1'b0;
    end else if(N2137) begin
      mem[2029] <= N2183;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2028] <= 1'b0;
    end else if(N2137) begin
      mem[2028] <= N2182;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2027] <= 1'b0;
    end else if(N2137) begin
      mem[2027] <= N2181;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2026] <= 1'b0;
    end else if(N2137) begin
      mem[2026] <= N2180;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2025] <= 1'b0;
    end else if(N2137) begin
      mem[2025] <= N2179;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2024] <= 1'b0;
    end else if(N2137) begin
      mem[2024] <= N2178;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2023] <= 1'b0;
    end else if(N2137) begin
      mem[2023] <= N2177;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2022] <= 1'b0;
    end else if(N2137) begin
      mem[2022] <= N2176;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2021] <= 1'b0;
    end else if(N2137) begin
      mem[2021] <= N2175;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2020] <= 1'b0;
    end else if(N2137) begin
      mem[2020] <= N2174;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2019] <= 1'b0;
    end else if(N2137) begin
      mem[2019] <= N2173;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2018] <= 1'b0;
    end else if(N2137) begin
      mem[2018] <= N2172;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2017] <= 1'b0;
    end else if(N2137) begin
      mem[2017] <= N2171;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2016] <= 1'b0;
    end else if(N2137) begin
      mem[2016] <= N2170;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2015] <= 1'b0;
    end else if(N2137) begin
      mem[2015] <= N2169;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2014] <= 1'b0;
    end else if(N2137) begin
      mem[2014] <= N2168;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2013] <= 1'b0;
    end else if(N2137) begin
      mem[2013] <= N2167;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2012] <= 1'b0;
    end else if(N2137) begin
      mem[2012] <= N2166;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2011] <= 1'b0;
    end else if(N2137) begin
      mem[2011] <= N2165;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2010] <= 1'b0;
    end else if(N2137) begin
      mem[2010] <= N2164;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2009] <= 1'b0;
    end else if(N2137) begin
      mem[2009] <= N2163;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2008] <= 1'b0;
    end else if(N2137) begin
      mem[2008] <= N2162;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2007] <= 1'b0;
    end else if(N2137) begin
      mem[2007] <= N2161;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2006] <= 1'b0;
    end else if(N2137) begin
      mem[2006] <= N2160;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2005] <= 1'b0;
    end else if(N2137) begin
      mem[2005] <= N2159;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2004] <= 1'b0;
    end else if(N2137) begin
      mem[2004] <= N2158;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2003] <= 1'b0;
    end else if(N2137) begin
      mem[2003] <= N2157;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2002] <= 1'b0;
    end else if(N2137) begin
      mem[2002] <= N2156;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2001] <= 1'b0;
    end else if(N2137) begin
      mem[2001] <= N2155;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2000] <= 1'b0;
    end else if(N2137) begin
      mem[2000] <= N2154;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1999] <= 1'b0;
    end else if(N2137) begin
      mem[1999] <= N2153;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1998] <= 1'b0;
    end else if(N2137) begin
      mem[1998] <= N2152;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1997] <= 1'b0;
    end else if(N2137) begin
      mem[1997] <= N2151;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1996] <= 1'b0;
    end else if(N2137) begin
      mem[1996] <= N2150;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1995] <= 1'b0;
    end else if(N2137) begin
      mem[1995] <= N2149;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1994] <= 1'b0;
    end else if(N2137) begin
      mem[1994] <= N2148;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1993] <= 1'b0;
    end else if(N2137) begin
      mem[1993] <= N2147;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1992] <= 1'b0;
    end else if(N2137) begin
      mem[1992] <= N2146;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1991] <= 1'b0;
    end else if(N2137) begin
      mem[1991] <= N2145;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1990] <= 1'b0;
    end else if(N2137) begin
      mem[1990] <= N2144;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1989] <= 1'b0;
    end else if(N2137) begin
      mem[1989] <= N2143;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1988] <= 1'b0;
    end else if(N2137) begin
      mem[1988] <= N2142;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1987] <= 1'b0;
    end else if(N2137) begin
      mem[1987] <= N2141;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1986] <= 1'b0;
    end else if(N2137) begin
      mem[1986] <= N2140;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1985] <= 1'b0;
    end else if(N2137) begin
      mem[1985] <= N2139;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1984] <= 1'b0;
    end else if(N2137) begin
      mem[1984] <= N2138;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1983] <= 1'b0;
    end else if(N2071) begin
      mem[1983] <= N2135;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1982] <= 1'b0;
    end else if(N2071) begin
      mem[1982] <= N2134;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1981] <= 1'b0;
    end else if(N2071) begin
      mem[1981] <= N2133;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1980] <= 1'b0;
    end else if(N2071) begin
      mem[1980] <= N2132;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1979] <= 1'b0;
    end else if(N2071) begin
      mem[1979] <= N2131;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1978] <= 1'b0;
    end else if(N2071) begin
      mem[1978] <= N2130;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1977] <= 1'b0;
    end else if(N2071) begin
      mem[1977] <= N2129;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1976] <= 1'b0;
    end else if(N2071) begin
      mem[1976] <= N2128;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1975] <= 1'b0;
    end else if(N2071) begin
      mem[1975] <= N2127;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1974] <= 1'b0;
    end else if(N2071) begin
      mem[1974] <= N2126;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1973] <= 1'b0;
    end else if(N2071) begin
      mem[1973] <= N2125;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1972] <= 1'b0;
    end else if(N2071) begin
      mem[1972] <= N2124;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1971] <= 1'b0;
    end else if(N2071) begin
      mem[1971] <= N2123;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1970] <= 1'b0;
    end else if(N2071) begin
      mem[1970] <= N2122;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1969] <= 1'b0;
    end else if(N2071) begin
      mem[1969] <= N2121;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1968] <= 1'b0;
    end else if(N2071) begin
      mem[1968] <= N2120;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1967] <= 1'b0;
    end else if(N2071) begin
      mem[1967] <= N2119;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1966] <= 1'b0;
    end else if(N2071) begin
      mem[1966] <= N2118;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1965] <= 1'b0;
    end else if(N2071) begin
      mem[1965] <= N2117;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1964] <= 1'b0;
    end else if(N2071) begin
      mem[1964] <= N2116;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1963] <= 1'b0;
    end else if(N2071) begin
      mem[1963] <= N2115;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1962] <= 1'b0;
    end else if(N2071) begin
      mem[1962] <= N2114;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1961] <= 1'b0;
    end else if(N2071) begin
      mem[1961] <= N2113;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1960] <= 1'b0;
    end else if(N2071) begin
      mem[1960] <= N2112;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1959] <= 1'b0;
    end else if(N2071) begin
      mem[1959] <= N2111;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1958] <= 1'b0;
    end else if(N2071) begin
      mem[1958] <= N2110;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1957] <= 1'b0;
    end else if(N2071) begin
      mem[1957] <= N2109;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1956] <= 1'b0;
    end else if(N2071) begin
      mem[1956] <= N2108;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1955] <= 1'b0;
    end else if(N2071) begin
      mem[1955] <= N2107;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1954] <= 1'b0;
    end else if(N2071) begin
      mem[1954] <= N2106;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1953] <= 1'b0;
    end else if(N2071) begin
      mem[1953] <= N2105;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1952] <= 1'b0;
    end else if(N2071) begin
      mem[1952] <= N2104;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1951] <= 1'b0;
    end else if(N2071) begin
      mem[1951] <= N2103;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1950] <= 1'b0;
    end else if(N2071) begin
      mem[1950] <= N2102;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1949] <= 1'b0;
    end else if(N2071) begin
      mem[1949] <= N2101;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1948] <= 1'b0;
    end else if(N2071) begin
      mem[1948] <= N2100;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1947] <= 1'b0;
    end else if(N2071) begin
      mem[1947] <= N2099;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1946] <= 1'b0;
    end else if(N2071) begin
      mem[1946] <= N2098;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1945] <= 1'b0;
    end else if(N2071) begin
      mem[1945] <= N2097;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1944] <= 1'b0;
    end else if(N2071) begin
      mem[1944] <= N2096;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1943] <= 1'b0;
    end else if(N2071) begin
      mem[1943] <= N2095;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1942] <= 1'b0;
    end else if(N2071) begin
      mem[1942] <= N2094;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1941] <= 1'b0;
    end else if(N2071) begin
      mem[1941] <= N2093;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1940] <= 1'b0;
    end else if(N2071) begin
      mem[1940] <= N2092;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1939] <= 1'b0;
    end else if(N2071) begin
      mem[1939] <= N2091;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1938] <= 1'b0;
    end else if(N2071) begin
      mem[1938] <= N2090;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1937] <= 1'b0;
    end else if(N2071) begin
      mem[1937] <= N2089;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1936] <= 1'b0;
    end else if(N2071) begin
      mem[1936] <= N2088;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1935] <= 1'b0;
    end else if(N2071) begin
      mem[1935] <= N2087;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1934] <= 1'b0;
    end else if(N2071) begin
      mem[1934] <= N2086;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1933] <= 1'b0;
    end else if(N2071) begin
      mem[1933] <= N2085;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1932] <= 1'b0;
    end else if(N2071) begin
      mem[1932] <= N2084;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1931] <= 1'b0;
    end else if(N2071) begin
      mem[1931] <= N2083;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1930] <= 1'b0;
    end else if(N2071) begin
      mem[1930] <= N2082;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1929] <= 1'b0;
    end else if(N2071) begin
      mem[1929] <= N2081;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1928] <= 1'b0;
    end else if(N2071) begin
      mem[1928] <= N2080;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1927] <= 1'b0;
    end else if(N2071) begin
      mem[1927] <= N2079;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1926] <= 1'b0;
    end else if(N2071) begin
      mem[1926] <= N2078;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1925] <= 1'b0;
    end else if(N2071) begin
      mem[1925] <= N2077;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1924] <= 1'b0;
    end else if(N2071) begin
      mem[1924] <= N2076;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1923] <= 1'b0;
    end else if(N2071) begin
      mem[1923] <= N2075;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1922] <= 1'b0;
    end else if(N2071) begin
      mem[1922] <= N2074;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1921] <= 1'b0;
    end else if(N2071) begin
      mem[1921] <= N2073;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1920] <= 1'b0;
    end else if(N2071) begin
      mem[1920] <= N2072;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1919] <= 1'b0;
    end else if(N2005) begin
      mem[1919] <= N2069;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1918] <= 1'b0;
    end else if(N2005) begin
      mem[1918] <= N2068;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1917] <= 1'b0;
    end else if(N2005) begin
      mem[1917] <= N2067;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1916] <= 1'b0;
    end else if(N2005) begin
      mem[1916] <= N2066;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1915] <= 1'b0;
    end else if(N2005) begin
      mem[1915] <= N2065;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1914] <= 1'b0;
    end else if(N2005) begin
      mem[1914] <= N2064;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1913] <= 1'b0;
    end else if(N2005) begin
      mem[1913] <= N2063;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1912] <= 1'b0;
    end else if(N2005) begin
      mem[1912] <= N2062;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1911] <= 1'b0;
    end else if(N2005) begin
      mem[1911] <= N2061;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1910] <= 1'b0;
    end else if(N2005) begin
      mem[1910] <= N2060;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1909] <= 1'b0;
    end else if(N2005) begin
      mem[1909] <= N2059;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1908] <= 1'b0;
    end else if(N2005) begin
      mem[1908] <= N2058;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1907] <= 1'b0;
    end else if(N2005) begin
      mem[1907] <= N2057;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1906] <= 1'b0;
    end else if(N2005) begin
      mem[1906] <= N2056;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1905] <= 1'b0;
    end else if(N2005) begin
      mem[1905] <= N2055;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1904] <= 1'b0;
    end else if(N2005) begin
      mem[1904] <= N2054;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1903] <= 1'b0;
    end else if(N2005) begin
      mem[1903] <= N2053;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1902] <= 1'b0;
    end else if(N2005) begin
      mem[1902] <= N2052;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1901] <= 1'b0;
    end else if(N2005) begin
      mem[1901] <= N2051;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1900] <= 1'b0;
    end else if(N2005) begin
      mem[1900] <= N2050;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1899] <= 1'b0;
    end else if(N2005) begin
      mem[1899] <= N2049;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1898] <= 1'b0;
    end else if(N2005) begin
      mem[1898] <= N2048;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1897] <= 1'b0;
    end else if(N2005) begin
      mem[1897] <= N2047;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1896] <= 1'b0;
    end else if(N2005) begin
      mem[1896] <= N2046;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1895] <= 1'b0;
    end else if(N2005) begin
      mem[1895] <= N2045;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1894] <= 1'b0;
    end else if(N2005) begin
      mem[1894] <= N2044;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1893] <= 1'b0;
    end else if(N2005) begin
      mem[1893] <= N2043;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1892] <= 1'b0;
    end else if(N2005) begin
      mem[1892] <= N2042;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1891] <= 1'b0;
    end else if(N2005) begin
      mem[1891] <= N2041;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1890] <= 1'b0;
    end else if(N2005) begin
      mem[1890] <= N2040;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1889] <= 1'b0;
    end else if(N2005) begin
      mem[1889] <= N2039;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1888] <= 1'b0;
    end else if(N2005) begin
      mem[1888] <= N2038;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1887] <= 1'b0;
    end else if(N2005) begin
      mem[1887] <= N2037;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1886] <= 1'b0;
    end else if(N2005) begin
      mem[1886] <= N2036;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1885] <= 1'b0;
    end else if(N2005) begin
      mem[1885] <= N2035;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1884] <= 1'b0;
    end else if(N2005) begin
      mem[1884] <= N2034;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1883] <= 1'b0;
    end else if(N2005) begin
      mem[1883] <= N2033;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1882] <= 1'b0;
    end else if(N2005) begin
      mem[1882] <= N2032;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1881] <= 1'b0;
    end else if(N2005) begin
      mem[1881] <= N2031;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1880] <= 1'b0;
    end else if(N2005) begin
      mem[1880] <= N2030;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1879] <= 1'b0;
    end else if(N2005) begin
      mem[1879] <= N2029;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1878] <= 1'b0;
    end else if(N2005) begin
      mem[1878] <= N2028;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1877] <= 1'b0;
    end else if(N2005) begin
      mem[1877] <= N2027;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1876] <= 1'b0;
    end else if(N2005) begin
      mem[1876] <= N2026;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1875] <= 1'b0;
    end else if(N2005) begin
      mem[1875] <= N2025;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1874] <= 1'b0;
    end else if(N2005) begin
      mem[1874] <= N2024;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1873] <= 1'b0;
    end else if(N2005) begin
      mem[1873] <= N2023;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1872] <= 1'b0;
    end else if(N2005) begin
      mem[1872] <= N2022;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1871] <= 1'b0;
    end else if(N2005) begin
      mem[1871] <= N2021;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1870] <= 1'b0;
    end else if(N2005) begin
      mem[1870] <= N2020;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1869] <= 1'b0;
    end else if(N2005) begin
      mem[1869] <= N2019;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1868] <= 1'b0;
    end else if(N2005) begin
      mem[1868] <= N2018;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1867] <= 1'b0;
    end else if(N2005) begin
      mem[1867] <= N2017;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1866] <= 1'b0;
    end else if(N2005) begin
      mem[1866] <= N2016;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1865] <= 1'b0;
    end else if(N2005) begin
      mem[1865] <= N2015;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1864] <= 1'b0;
    end else if(N2005) begin
      mem[1864] <= N2014;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1863] <= 1'b0;
    end else if(N2005) begin
      mem[1863] <= N2013;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1862] <= 1'b0;
    end else if(N2005) begin
      mem[1862] <= N2012;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1861] <= 1'b0;
    end else if(N2005) begin
      mem[1861] <= N2011;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1860] <= 1'b0;
    end else if(N2005) begin
      mem[1860] <= N2010;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1859] <= 1'b0;
    end else if(N2005) begin
      mem[1859] <= N2009;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1858] <= 1'b0;
    end else if(N2005) begin
      mem[1858] <= N2008;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1857] <= 1'b0;
    end else if(N2005) begin
      mem[1857] <= N2007;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1856] <= 1'b0;
    end else if(N2005) begin
      mem[1856] <= N2006;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1855] <= 1'b0;
    end else if(N1939) begin
      mem[1855] <= N2003;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1854] <= 1'b0;
    end else if(N1939) begin
      mem[1854] <= N2002;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1853] <= 1'b0;
    end else if(N1939) begin
      mem[1853] <= N2001;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1852] <= 1'b0;
    end else if(N1939) begin
      mem[1852] <= N2000;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1851] <= 1'b0;
    end else if(N1939) begin
      mem[1851] <= N1999;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1850] <= 1'b0;
    end else if(N1939) begin
      mem[1850] <= N1998;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1849] <= 1'b0;
    end else if(N1939) begin
      mem[1849] <= N1997;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1848] <= 1'b0;
    end else if(N1939) begin
      mem[1848] <= N1996;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1847] <= 1'b0;
    end else if(N1939) begin
      mem[1847] <= N1995;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1846] <= 1'b0;
    end else if(N1939) begin
      mem[1846] <= N1994;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1845] <= 1'b0;
    end else if(N1939) begin
      mem[1845] <= N1993;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1844] <= 1'b0;
    end else if(N1939) begin
      mem[1844] <= N1992;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1843] <= 1'b0;
    end else if(N1939) begin
      mem[1843] <= N1991;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1842] <= 1'b0;
    end else if(N1939) begin
      mem[1842] <= N1990;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1841] <= 1'b0;
    end else if(N1939) begin
      mem[1841] <= N1989;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1840] <= 1'b0;
    end else if(N1939) begin
      mem[1840] <= N1988;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1839] <= 1'b0;
    end else if(N1939) begin
      mem[1839] <= N1987;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1838] <= 1'b0;
    end else if(N1939) begin
      mem[1838] <= N1986;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1837] <= 1'b0;
    end else if(N1939) begin
      mem[1837] <= N1985;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1836] <= 1'b0;
    end else if(N1939) begin
      mem[1836] <= N1984;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1835] <= 1'b0;
    end else if(N1939) begin
      mem[1835] <= N1983;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1834] <= 1'b0;
    end else if(N1939) begin
      mem[1834] <= N1982;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1833] <= 1'b0;
    end else if(N1939) begin
      mem[1833] <= N1981;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1832] <= 1'b0;
    end else if(N1939) begin
      mem[1832] <= N1980;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1831] <= 1'b0;
    end else if(N1939) begin
      mem[1831] <= N1979;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1830] <= 1'b0;
    end else if(N1939) begin
      mem[1830] <= N1978;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1829] <= 1'b0;
    end else if(N1939) begin
      mem[1829] <= N1977;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1828] <= 1'b0;
    end else if(N1939) begin
      mem[1828] <= N1976;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1827] <= 1'b0;
    end else if(N1939) begin
      mem[1827] <= N1975;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1826] <= 1'b0;
    end else if(N1939) begin
      mem[1826] <= N1974;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1825] <= 1'b0;
    end else if(N1939) begin
      mem[1825] <= N1973;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1824] <= 1'b0;
    end else if(N1939) begin
      mem[1824] <= N1972;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1823] <= 1'b0;
    end else if(N1939) begin
      mem[1823] <= N1971;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1822] <= 1'b0;
    end else if(N1939) begin
      mem[1822] <= N1970;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1821] <= 1'b0;
    end else if(N1939) begin
      mem[1821] <= N1969;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1820] <= 1'b0;
    end else if(N1939) begin
      mem[1820] <= N1968;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1819] <= 1'b0;
    end else if(N1939) begin
      mem[1819] <= N1967;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1818] <= 1'b0;
    end else if(N1939) begin
      mem[1818] <= N1966;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1817] <= 1'b0;
    end else if(N1939) begin
      mem[1817] <= N1965;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1816] <= 1'b0;
    end else if(N1939) begin
      mem[1816] <= N1964;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1815] <= 1'b0;
    end else if(N1939) begin
      mem[1815] <= N1963;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1814] <= 1'b0;
    end else if(N1939) begin
      mem[1814] <= N1962;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1813] <= 1'b0;
    end else if(N1939) begin
      mem[1813] <= N1961;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1812] <= 1'b0;
    end else if(N1939) begin
      mem[1812] <= N1960;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1811] <= 1'b0;
    end else if(N1939) begin
      mem[1811] <= N1959;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1810] <= 1'b0;
    end else if(N1939) begin
      mem[1810] <= N1958;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1809] <= 1'b0;
    end else if(N1939) begin
      mem[1809] <= N1957;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1808] <= 1'b0;
    end else if(N1939) begin
      mem[1808] <= N1956;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1807] <= 1'b0;
    end else if(N1939) begin
      mem[1807] <= N1955;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1806] <= 1'b0;
    end else if(N1939) begin
      mem[1806] <= N1954;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1805] <= 1'b0;
    end else if(N1939) begin
      mem[1805] <= N1953;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1804] <= 1'b0;
    end else if(N1939) begin
      mem[1804] <= N1952;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1803] <= 1'b0;
    end else if(N1939) begin
      mem[1803] <= N1951;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1802] <= 1'b0;
    end else if(N1939) begin
      mem[1802] <= N1950;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1801] <= 1'b0;
    end else if(N1939) begin
      mem[1801] <= N1949;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1800] <= 1'b0;
    end else if(N1939) begin
      mem[1800] <= N1948;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1799] <= 1'b0;
    end else if(N1939) begin
      mem[1799] <= N1947;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1798] <= 1'b0;
    end else if(N1939) begin
      mem[1798] <= N1946;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1797] <= 1'b0;
    end else if(N1939) begin
      mem[1797] <= N1945;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1796] <= 1'b0;
    end else if(N1939) begin
      mem[1796] <= N1944;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1795] <= 1'b0;
    end else if(N1939) begin
      mem[1795] <= N1943;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1794] <= 1'b0;
    end else if(N1939) begin
      mem[1794] <= N1942;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1793] <= 1'b0;
    end else if(N1939) begin
      mem[1793] <= N1941;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1792] <= 1'b0;
    end else if(N1939) begin
      mem[1792] <= N1940;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1791] <= 1'b0;
    end else if(N1873) begin
      mem[1791] <= N1937;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1790] <= 1'b0;
    end else if(N1873) begin
      mem[1790] <= N1936;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1789] <= 1'b0;
    end else if(N1873) begin
      mem[1789] <= N1935;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1788] <= 1'b0;
    end else if(N1873) begin
      mem[1788] <= N1934;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1787] <= 1'b0;
    end else if(N1873) begin
      mem[1787] <= N1933;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1786] <= 1'b0;
    end else if(N1873) begin
      mem[1786] <= N1932;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1785] <= 1'b0;
    end else if(N1873) begin
      mem[1785] <= N1931;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1784] <= 1'b0;
    end else if(N1873) begin
      mem[1784] <= N1930;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1783] <= 1'b0;
    end else if(N1873) begin
      mem[1783] <= N1929;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1782] <= 1'b0;
    end else if(N1873) begin
      mem[1782] <= N1928;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1781] <= 1'b0;
    end else if(N1873) begin
      mem[1781] <= N1927;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1780] <= 1'b0;
    end else if(N1873) begin
      mem[1780] <= N1926;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1779] <= 1'b0;
    end else if(N1873) begin
      mem[1779] <= N1925;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1778] <= 1'b0;
    end else if(N1873) begin
      mem[1778] <= N1924;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1777] <= 1'b0;
    end else if(N1873) begin
      mem[1777] <= N1923;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1776] <= 1'b0;
    end else if(N1873) begin
      mem[1776] <= N1922;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1775] <= 1'b0;
    end else if(N1873) begin
      mem[1775] <= N1921;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1774] <= 1'b0;
    end else if(N1873) begin
      mem[1774] <= N1920;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1773] <= 1'b0;
    end else if(N1873) begin
      mem[1773] <= N1919;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1772] <= 1'b0;
    end else if(N1873) begin
      mem[1772] <= N1918;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1771] <= 1'b0;
    end else if(N1873) begin
      mem[1771] <= N1917;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1770] <= 1'b0;
    end else if(N1873) begin
      mem[1770] <= N1916;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1769] <= 1'b0;
    end else if(N1873) begin
      mem[1769] <= N1915;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1768] <= 1'b0;
    end else if(N1873) begin
      mem[1768] <= N1914;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1767] <= 1'b0;
    end else if(N1873) begin
      mem[1767] <= N1913;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1766] <= 1'b0;
    end else if(N1873) begin
      mem[1766] <= N1912;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1765] <= 1'b0;
    end else if(N1873) begin
      mem[1765] <= N1911;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1764] <= 1'b0;
    end else if(N1873) begin
      mem[1764] <= N1910;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1763] <= 1'b0;
    end else if(N1873) begin
      mem[1763] <= N1909;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1762] <= 1'b0;
    end else if(N1873) begin
      mem[1762] <= N1908;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1761] <= 1'b0;
    end else if(N1873) begin
      mem[1761] <= N1907;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1760] <= 1'b0;
    end else if(N1873) begin
      mem[1760] <= N1906;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1759] <= 1'b0;
    end else if(N1873) begin
      mem[1759] <= N1905;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1758] <= 1'b0;
    end else if(N1873) begin
      mem[1758] <= N1904;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1757] <= 1'b0;
    end else if(N1873) begin
      mem[1757] <= N1903;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1756] <= 1'b0;
    end else if(N1873) begin
      mem[1756] <= N1902;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1755] <= 1'b0;
    end else if(N1873) begin
      mem[1755] <= N1901;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1754] <= 1'b0;
    end else if(N1873) begin
      mem[1754] <= N1900;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1753] <= 1'b0;
    end else if(N1873) begin
      mem[1753] <= N1899;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1752] <= 1'b0;
    end else if(N1873) begin
      mem[1752] <= N1898;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1751] <= 1'b0;
    end else if(N1873) begin
      mem[1751] <= N1897;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1750] <= 1'b0;
    end else if(N1873) begin
      mem[1750] <= N1896;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1749] <= 1'b0;
    end else if(N1873) begin
      mem[1749] <= N1895;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1748] <= 1'b0;
    end else if(N1873) begin
      mem[1748] <= N1894;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1747] <= 1'b0;
    end else if(N1873) begin
      mem[1747] <= N1893;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1746] <= 1'b0;
    end else if(N1873) begin
      mem[1746] <= N1892;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1745] <= 1'b0;
    end else if(N1873) begin
      mem[1745] <= N1891;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1744] <= 1'b0;
    end else if(N1873) begin
      mem[1744] <= N1890;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1743] <= 1'b0;
    end else if(N1873) begin
      mem[1743] <= N1889;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1742] <= 1'b0;
    end else if(N1873) begin
      mem[1742] <= N1888;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1741] <= 1'b0;
    end else if(N1873) begin
      mem[1741] <= N1887;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1740] <= 1'b0;
    end else if(N1873) begin
      mem[1740] <= N1886;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1739] <= 1'b0;
    end else if(N1873) begin
      mem[1739] <= N1885;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1738] <= 1'b0;
    end else if(N1873) begin
      mem[1738] <= N1884;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1737] <= 1'b0;
    end else if(N1873) begin
      mem[1737] <= N1883;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1736] <= 1'b0;
    end else if(N1873) begin
      mem[1736] <= N1882;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1735] <= 1'b0;
    end else if(N1873) begin
      mem[1735] <= N1881;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1734] <= 1'b0;
    end else if(N1873) begin
      mem[1734] <= N1880;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1733] <= 1'b0;
    end else if(N1873) begin
      mem[1733] <= N1879;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1732] <= 1'b0;
    end else if(N1873) begin
      mem[1732] <= N1878;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1731] <= 1'b0;
    end else if(N1873) begin
      mem[1731] <= N1877;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1730] <= 1'b0;
    end else if(N1873) begin
      mem[1730] <= N1876;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1729] <= 1'b0;
    end else if(N1873) begin
      mem[1729] <= N1875;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1728] <= 1'b0;
    end else if(N1873) begin
      mem[1728] <= N1874;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1727] <= 1'b0;
    end else if(N1807) begin
      mem[1727] <= N1871;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1726] <= 1'b0;
    end else if(N1807) begin
      mem[1726] <= N1870;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1725] <= 1'b0;
    end else if(N1807) begin
      mem[1725] <= N1869;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1724] <= 1'b0;
    end else if(N1807) begin
      mem[1724] <= N1868;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1723] <= 1'b0;
    end else if(N1807) begin
      mem[1723] <= N1867;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1722] <= 1'b0;
    end else if(N1807) begin
      mem[1722] <= N1866;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1721] <= 1'b0;
    end else if(N1807) begin
      mem[1721] <= N1865;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1720] <= 1'b0;
    end else if(N1807) begin
      mem[1720] <= N1864;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1719] <= 1'b0;
    end else if(N1807) begin
      mem[1719] <= N1863;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1718] <= 1'b0;
    end else if(N1807) begin
      mem[1718] <= N1862;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1717] <= 1'b0;
    end else if(N1807) begin
      mem[1717] <= N1861;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1716] <= 1'b0;
    end else if(N1807) begin
      mem[1716] <= N1860;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1715] <= 1'b0;
    end else if(N1807) begin
      mem[1715] <= N1859;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1714] <= 1'b0;
    end else if(N1807) begin
      mem[1714] <= N1858;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1713] <= 1'b0;
    end else if(N1807) begin
      mem[1713] <= N1857;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1712] <= 1'b0;
    end else if(N1807) begin
      mem[1712] <= N1856;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1711] <= 1'b0;
    end else if(N1807) begin
      mem[1711] <= N1855;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1710] <= 1'b0;
    end else if(N1807) begin
      mem[1710] <= N1854;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1709] <= 1'b0;
    end else if(N1807) begin
      mem[1709] <= N1853;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1708] <= 1'b0;
    end else if(N1807) begin
      mem[1708] <= N1852;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1707] <= 1'b0;
    end else if(N1807) begin
      mem[1707] <= N1851;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1706] <= 1'b0;
    end else if(N1807) begin
      mem[1706] <= N1850;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1705] <= 1'b0;
    end else if(N1807) begin
      mem[1705] <= N1849;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1704] <= 1'b0;
    end else if(N1807) begin
      mem[1704] <= N1848;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1703] <= 1'b0;
    end else if(N1807) begin
      mem[1703] <= N1847;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1702] <= 1'b0;
    end else if(N1807) begin
      mem[1702] <= N1846;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1701] <= 1'b0;
    end else if(N1807) begin
      mem[1701] <= N1845;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1700] <= 1'b0;
    end else if(N1807) begin
      mem[1700] <= N1844;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1699] <= 1'b0;
    end else if(N1807) begin
      mem[1699] <= N1843;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1698] <= 1'b0;
    end else if(N1807) begin
      mem[1698] <= N1842;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1697] <= 1'b0;
    end else if(N1807) begin
      mem[1697] <= N1841;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1696] <= 1'b0;
    end else if(N1807) begin
      mem[1696] <= N1840;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1695] <= 1'b0;
    end else if(N1807) begin
      mem[1695] <= N1839;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1694] <= 1'b0;
    end else if(N1807) begin
      mem[1694] <= N1838;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1693] <= 1'b0;
    end else if(N1807) begin
      mem[1693] <= N1837;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1692] <= 1'b0;
    end else if(N1807) begin
      mem[1692] <= N1836;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1691] <= 1'b0;
    end else if(N1807) begin
      mem[1691] <= N1835;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1690] <= 1'b0;
    end else if(N1807) begin
      mem[1690] <= N1834;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1689] <= 1'b0;
    end else if(N1807) begin
      mem[1689] <= N1833;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1688] <= 1'b0;
    end else if(N1807) begin
      mem[1688] <= N1832;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1687] <= 1'b0;
    end else if(N1807) begin
      mem[1687] <= N1831;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1686] <= 1'b0;
    end else if(N1807) begin
      mem[1686] <= N1830;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1685] <= 1'b0;
    end else if(N1807) begin
      mem[1685] <= N1829;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1684] <= 1'b0;
    end else if(N1807) begin
      mem[1684] <= N1828;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1683] <= 1'b0;
    end else if(N1807) begin
      mem[1683] <= N1827;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1682] <= 1'b0;
    end else if(N1807) begin
      mem[1682] <= N1826;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1681] <= 1'b0;
    end else if(N1807) begin
      mem[1681] <= N1825;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1680] <= 1'b0;
    end else if(N1807) begin
      mem[1680] <= N1824;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1679] <= 1'b0;
    end else if(N1807) begin
      mem[1679] <= N1823;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1678] <= 1'b0;
    end else if(N1807) begin
      mem[1678] <= N1822;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1677] <= 1'b0;
    end else if(N1807) begin
      mem[1677] <= N1821;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1676] <= 1'b0;
    end else if(N1807) begin
      mem[1676] <= N1820;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1675] <= 1'b0;
    end else if(N1807) begin
      mem[1675] <= N1819;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1674] <= 1'b0;
    end else if(N1807) begin
      mem[1674] <= N1818;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1673] <= 1'b0;
    end else if(N1807) begin
      mem[1673] <= N1817;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1672] <= 1'b0;
    end else if(N1807) begin
      mem[1672] <= N1816;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1671] <= 1'b0;
    end else if(N1807) begin
      mem[1671] <= N1815;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1670] <= 1'b0;
    end else if(N1807) begin
      mem[1670] <= N1814;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1669] <= 1'b0;
    end else if(N1807) begin
      mem[1669] <= N1813;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1668] <= 1'b0;
    end else if(N1807) begin
      mem[1668] <= N1812;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1667] <= 1'b0;
    end else if(N1807) begin
      mem[1667] <= N1811;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1666] <= 1'b0;
    end else if(N1807) begin
      mem[1666] <= N1810;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1665] <= 1'b0;
    end else if(N1807) begin
      mem[1665] <= N1809;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1664] <= 1'b0;
    end else if(N1807) begin
      mem[1664] <= N1808;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1663] <= 1'b0;
    end else if(N1741) begin
      mem[1663] <= N1805;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1662] <= 1'b0;
    end else if(N1741) begin
      mem[1662] <= N1804;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1661] <= 1'b0;
    end else if(N1741) begin
      mem[1661] <= N1803;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1660] <= 1'b0;
    end else if(N1741) begin
      mem[1660] <= N1802;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1659] <= 1'b0;
    end else if(N1741) begin
      mem[1659] <= N1801;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1658] <= 1'b0;
    end else if(N1741) begin
      mem[1658] <= N1800;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1657] <= 1'b0;
    end else if(N1741) begin
      mem[1657] <= N1799;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1656] <= 1'b0;
    end else if(N1741) begin
      mem[1656] <= N1798;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1655] <= 1'b0;
    end else if(N1741) begin
      mem[1655] <= N1797;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1654] <= 1'b0;
    end else if(N1741) begin
      mem[1654] <= N1796;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1653] <= 1'b0;
    end else if(N1741) begin
      mem[1653] <= N1795;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1652] <= 1'b0;
    end else if(N1741) begin
      mem[1652] <= N1794;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1651] <= 1'b0;
    end else if(N1741) begin
      mem[1651] <= N1793;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1650] <= 1'b0;
    end else if(N1741) begin
      mem[1650] <= N1792;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1649] <= 1'b0;
    end else if(N1741) begin
      mem[1649] <= N1791;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1648] <= 1'b0;
    end else if(N1741) begin
      mem[1648] <= N1790;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1647] <= 1'b0;
    end else if(N1741) begin
      mem[1647] <= N1789;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1646] <= 1'b0;
    end else if(N1741) begin
      mem[1646] <= N1788;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1645] <= 1'b0;
    end else if(N1741) begin
      mem[1645] <= N1787;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1644] <= 1'b0;
    end else if(N1741) begin
      mem[1644] <= N1786;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1643] <= 1'b0;
    end else if(N1741) begin
      mem[1643] <= N1785;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1642] <= 1'b0;
    end else if(N1741) begin
      mem[1642] <= N1784;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1641] <= 1'b0;
    end else if(N1741) begin
      mem[1641] <= N1783;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1640] <= 1'b0;
    end else if(N1741) begin
      mem[1640] <= N1782;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1639] <= 1'b0;
    end else if(N1741) begin
      mem[1639] <= N1781;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1638] <= 1'b0;
    end else if(N1741) begin
      mem[1638] <= N1780;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1637] <= 1'b0;
    end else if(N1741) begin
      mem[1637] <= N1779;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1636] <= 1'b0;
    end else if(N1741) begin
      mem[1636] <= N1778;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1635] <= 1'b0;
    end else if(N1741) begin
      mem[1635] <= N1777;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1634] <= 1'b0;
    end else if(N1741) begin
      mem[1634] <= N1776;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1633] <= 1'b0;
    end else if(N1741) begin
      mem[1633] <= N1775;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1632] <= 1'b0;
    end else if(N1741) begin
      mem[1632] <= N1774;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1631] <= 1'b0;
    end else if(N1741) begin
      mem[1631] <= N1773;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1630] <= 1'b0;
    end else if(N1741) begin
      mem[1630] <= N1772;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1629] <= 1'b0;
    end else if(N1741) begin
      mem[1629] <= N1771;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1628] <= 1'b0;
    end else if(N1741) begin
      mem[1628] <= N1770;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1627] <= 1'b0;
    end else if(N1741) begin
      mem[1627] <= N1769;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1626] <= 1'b0;
    end else if(N1741) begin
      mem[1626] <= N1768;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1625] <= 1'b0;
    end else if(N1741) begin
      mem[1625] <= N1767;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1624] <= 1'b0;
    end else if(N1741) begin
      mem[1624] <= N1766;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1623] <= 1'b0;
    end else if(N1741) begin
      mem[1623] <= N1765;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1622] <= 1'b0;
    end else if(N1741) begin
      mem[1622] <= N1764;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1621] <= 1'b0;
    end else if(N1741) begin
      mem[1621] <= N1763;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1620] <= 1'b0;
    end else if(N1741) begin
      mem[1620] <= N1762;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1619] <= 1'b0;
    end else if(N1741) begin
      mem[1619] <= N1761;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1618] <= 1'b0;
    end else if(N1741) begin
      mem[1618] <= N1760;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1617] <= 1'b0;
    end else if(N1741) begin
      mem[1617] <= N1759;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1616] <= 1'b0;
    end else if(N1741) begin
      mem[1616] <= N1758;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1615] <= 1'b0;
    end else if(N1741) begin
      mem[1615] <= N1757;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1614] <= 1'b0;
    end else if(N1741) begin
      mem[1614] <= N1756;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1613] <= 1'b0;
    end else if(N1741) begin
      mem[1613] <= N1755;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1612] <= 1'b0;
    end else if(N1741) begin
      mem[1612] <= N1754;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1611] <= 1'b0;
    end else if(N1741) begin
      mem[1611] <= N1753;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1610] <= 1'b0;
    end else if(N1741) begin
      mem[1610] <= N1752;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1609] <= 1'b0;
    end else if(N1741) begin
      mem[1609] <= N1751;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1608] <= 1'b0;
    end else if(N1741) begin
      mem[1608] <= N1750;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1607] <= 1'b0;
    end else if(N1741) begin
      mem[1607] <= N1749;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1606] <= 1'b0;
    end else if(N1741) begin
      mem[1606] <= N1748;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1605] <= 1'b0;
    end else if(N1741) begin
      mem[1605] <= N1747;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1604] <= 1'b0;
    end else if(N1741) begin
      mem[1604] <= N1746;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1603] <= 1'b0;
    end else if(N1741) begin
      mem[1603] <= N1745;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1602] <= 1'b0;
    end else if(N1741) begin
      mem[1602] <= N1744;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1601] <= 1'b0;
    end else if(N1741) begin
      mem[1601] <= N1743;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1600] <= 1'b0;
    end else if(N1741) begin
      mem[1600] <= N1742;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1599] <= 1'b0;
    end else if(N1675) begin
      mem[1599] <= N1739;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1598] <= 1'b0;
    end else if(N1675) begin
      mem[1598] <= N1738;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1597] <= 1'b0;
    end else if(N1675) begin
      mem[1597] <= N1737;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1596] <= 1'b0;
    end else if(N1675) begin
      mem[1596] <= N1736;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1595] <= 1'b0;
    end else if(N1675) begin
      mem[1595] <= N1735;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1594] <= 1'b0;
    end else if(N1675) begin
      mem[1594] <= N1734;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1593] <= 1'b0;
    end else if(N1675) begin
      mem[1593] <= N1733;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1592] <= 1'b0;
    end else if(N1675) begin
      mem[1592] <= N1732;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1591] <= 1'b0;
    end else if(N1675) begin
      mem[1591] <= N1731;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1590] <= 1'b0;
    end else if(N1675) begin
      mem[1590] <= N1730;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1589] <= 1'b0;
    end else if(N1675) begin
      mem[1589] <= N1729;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1588] <= 1'b0;
    end else if(N1675) begin
      mem[1588] <= N1728;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1587] <= 1'b0;
    end else if(N1675) begin
      mem[1587] <= N1727;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1586] <= 1'b0;
    end else if(N1675) begin
      mem[1586] <= N1726;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1585] <= 1'b0;
    end else if(N1675) begin
      mem[1585] <= N1725;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1584] <= 1'b0;
    end else if(N1675) begin
      mem[1584] <= N1724;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1583] <= 1'b0;
    end else if(N1675) begin
      mem[1583] <= N1723;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1582] <= 1'b0;
    end else if(N1675) begin
      mem[1582] <= N1722;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1581] <= 1'b0;
    end else if(N1675) begin
      mem[1581] <= N1721;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1580] <= 1'b0;
    end else if(N1675) begin
      mem[1580] <= N1720;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1579] <= 1'b0;
    end else if(N1675) begin
      mem[1579] <= N1719;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1578] <= 1'b0;
    end else if(N1675) begin
      mem[1578] <= N1718;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1577] <= 1'b0;
    end else if(N1675) begin
      mem[1577] <= N1717;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1576] <= 1'b0;
    end else if(N1675) begin
      mem[1576] <= N1716;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1575] <= 1'b0;
    end else if(N1675) begin
      mem[1575] <= N1715;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1574] <= 1'b0;
    end else if(N1675) begin
      mem[1574] <= N1714;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1573] <= 1'b0;
    end else if(N1675) begin
      mem[1573] <= N1713;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1572] <= 1'b0;
    end else if(N1675) begin
      mem[1572] <= N1712;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1571] <= 1'b0;
    end else if(N1675) begin
      mem[1571] <= N1711;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1570] <= 1'b0;
    end else if(N1675) begin
      mem[1570] <= N1710;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1569] <= 1'b0;
    end else if(N1675) begin
      mem[1569] <= N1709;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1568] <= 1'b0;
    end else if(N1675) begin
      mem[1568] <= N1708;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1567] <= 1'b0;
    end else if(N1675) begin
      mem[1567] <= N1707;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1566] <= 1'b0;
    end else if(N1675) begin
      mem[1566] <= N1706;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1565] <= 1'b0;
    end else if(N1675) begin
      mem[1565] <= N1705;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1564] <= 1'b0;
    end else if(N1675) begin
      mem[1564] <= N1704;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1563] <= 1'b0;
    end else if(N1675) begin
      mem[1563] <= N1703;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1562] <= 1'b0;
    end else if(N1675) begin
      mem[1562] <= N1702;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1561] <= 1'b0;
    end else if(N1675) begin
      mem[1561] <= N1701;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1560] <= 1'b0;
    end else if(N1675) begin
      mem[1560] <= N1700;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1559] <= 1'b0;
    end else if(N1675) begin
      mem[1559] <= N1699;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1558] <= 1'b0;
    end else if(N1675) begin
      mem[1558] <= N1698;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1557] <= 1'b0;
    end else if(N1675) begin
      mem[1557] <= N1697;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1556] <= 1'b0;
    end else if(N1675) begin
      mem[1556] <= N1696;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1555] <= 1'b0;
    end else if(N1675) begin
      mem[1555] <= N1695;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1554] <= 1'b0;
    end else if(N1675) begin
      mem[1554] <= N1694;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1553] <= 1'b0;
    end else if(N1675) begin
      mem[1553] <= N1693;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1552] <= 1'b0;
    end else if(N1675) begin
      mem[1552] <= N1692;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1551] <= 1'b0;
    end else if(N1675) begin
      mem[1551] <= N1691;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1550] <= 1'b0;
    end else if(N1675) begin
      mem[1550] <= N1690;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1549] <= 1'b0;
    end else if(N1675) begin
      mem[1549] <= N1689;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1548] <= 1'b0;
    end else if(N1675) begin
      mem[1548] <= N1688;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1547] <= 1'b0;
    end else if(N1675) begin
      mem[1547] <= N1687;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1546] <= 1'b0;
    end else if(N1675) begin
      mem[1546] <= N1686;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1545] <= 1'b0;
    end else if(N1675) begin
      mem[1545] <= N1685;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1544] <= 1'b0;
    end else if(N1675) begin
      mem[1544] <= N1684;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1543] <= 1'b0;
    end else if(N1675) begin
      mem[1543] <= N1683;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1542] <= 1'b0;
    end else if(N1675) begin
      mem[1542] <= N1682;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1541] <= 1'b0;
    end else if(N1675) begin
      mem[1541] <= N1681;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1540] <= 1'b0;
    end else if(N1675) begin
      mem[1540] <= N1680;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1539] <= 1'b0;
    end else if(N1675) begin
      mem[1539] <= N1679;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1538] <= 1'b0;
    end else if(N1675) begin
      mem[1538] <= N1678;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1537] <= 1'b0;
    end else if(N1675) begin
      mem[1537] <= N1677;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1536] <= 1'b0;
    end else if(N1675) begin
      mem[1536] <= N1676;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1535] <= 1'b0;
    end else if(N1609) begin
      mem[1535] <= N1673;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1534] <= 1'b0;
    end else if(N1609) begin
      mem[1534] <= N1672;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1533] <= 1'b0;
    end else if(N1609) begin
      mem[1533] <= N1671;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1532] <= 1'b0;
    end else if(N1609) begin
      mem[1532] <= N1670;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1531] <= 1'b0;
    end else if(N1609) begin
      mem[1531] <= N1669;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1530] <= 1'b0;
    end else if(N1609) begin
      mem[1530] <= N1668;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1529] <= 1'b0;
    end else if(N1609) begin
      mem[1529] <= N1667;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1528] <= 1'b0;
    end else if(N1609) begin
      mem[1528] <= N1666;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1527] <= 1'b0;
    end else if(N1609) begin
      mem[1527] <= N1665;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1526] <= 1'b0;
    end else if(N1609) begin
      mem[1526] <= N1664;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1525] <= 1'b0;
    end else if(N1609) begin
      mem[1525] <= N1663;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1524] <= 1'b0;
    end else if(N1609) begin
      mem[1524] <= N1662;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1523] <= 1'b0;
    end else if(N1609) begin
      mem[1523] <= N1661;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1522] <= 1'b0;
    end else if(N1609) begin
      mem[1522] <= N1660;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1521] <= 1'b0;
    end else if(N1609) begin
      mem[1521] <= N1659;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1520] <= 1'b0;
    end else if(N1609) begin
      mem[1520] <= N1658;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1519] <= 1'b0;
    end else if(N1609) begin
      mem[1519] <= N1657;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1518] <= 1'b0;
    end else if(N1609) begin
      mem[1518] <= N1656;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1517] <= 1'b0;
    end else if(N1609) begin
      mem[1517] <= N1655;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1516] <= 1'b0;
    end else if(N1609) begin
      mem[1516] <= N1654;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1515] <= 1'b0;
    end else if(N1609) begin
      mem[1515] <= N1653;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1514] <= 1'b0;
    end else if(N1609) begin
      mem[1514] <= N1652;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1513] <= 1'b0;
    end else if(N1609) begin
      mem[1513] <= N1651;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1512] <= 1'b0;
    end else if(N1609) begin
      mem[1512] <= N1650;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1511] <= 1'b0;
    end else if(N1609) begin
      mem[1511] <= N1649;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1510] <= 1'b0;
    end else if(N1609) begin
      mem[1510] <= N1648;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1509] <= 1'b0;
    end else if(N1609) begin
      mem[1509] <= N1647;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1508] <= 1'b0;
    end else if(N1609) begin
      mem[1508] <= N1646;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1507] <= 1'b0;
    end else if(N1609) begin
      mem[1507] <= N1645;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1506] <= 1'b0;
    end else if(N1609) begin
      mem[1506] <= N1644;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1505] <= 1'b0;
    end else if(N1609) begin
      mem[1505] <= N1643;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1504] <= 1'b0;
    end else if(N1609) begin
      mem[1504] <= N1642;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1503] <= 1'b0;
    end else if(N1609) begin
      mem[1503] <= N1641;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1502] <= 1'b0;
    end else if(N1609) begin
      mem[1502] <= N1640;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1501] <= 1'b0;
    end else if(N1609) begin
      mem[1501] <= N1639;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1500] <= 1'b0;
    end else if(N1609) begin
      mem[1500] <= N1638;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1499] <= 1'b0;
    end else if(N1609) begin
      mem[1499] <= N1637;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1498] <= 1'b0;
    end else if(N1609) begin
      mem[1498] <= N1636;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1497] <= 1'b0;
    end else if(N1609) begin
      mem[1497] <= N1635;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1496] <= 1'b0;
    end else if(N1609) begin
      mem[1496] <= N1634;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1495] <= 1'b0;
    end else if(N1609) begin
      mem[1495] <= N1633;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1494] <= 1'b0;
    end else if(N1609) begin
      mem[1494] <= N1632;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1493] <= 1'b0;
    end else if(N1609) begin
      mem[1493] <= N1631;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1492] <= 1'b0;
    end else if(N1609) begin
      mem[1492] <= N1630;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1491] <= 1'b0;
    end else if(N1609) begin
      mem[1491] <= N1629;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1490] <= 1'b0;
    end else if(N1609) begin
      mem[1490] <= N1628;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1489] <= 1'b0;
    end else if(N1609) begin
      mem[1489] <= N1627;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1488] <= 1'b0;
    end else if(N1609) begin
      mem[1488] <= N1626;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1487] <= 1'b0;
    end else if(N1609) begin
      mem[1487] <= N1625;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1486] <= 1'b0;
    end else if(N1609) begin
      mem[1486] <= N1624;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1485] <= 1'b0;
    end else if(N1609) begin
      mem[1485] <= N1623;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1484] <= 1'b0;
    end else if(N1609) begin
      mem[1484] <= N1622;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1483] <= 1'b0;
    end else if(N1609) begin
      mem[1483] <= N1621;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1482] <= 1'b0;
    end else if(N1609) begin
      mem[1482] <= N1620;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1481] <= 1'b0;
    end else if(N1609) begin
      mem[1481] <= N1619;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1480] <= 1'b0;
    end else if(N1609) begin
      mem[1480] <= N1618;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1479] <= 1'b0;
    end else if(N1609) begin
      mem[1479] <= N1617;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1478] <= 1'b0;
    end else if(N1609) begin
      mem[1478] <= N1616;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1477] <= 1'b0;
    end else if(N1609) begin
      mem[1477] <= N1615;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1476] <= 1'b0;
    end else if(N1609) begin
      mem[1476] <= N1614;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1475] <= 1'b0;
    end else if(N1609) begin
      mem[1475] <= N1613;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1474] <= 1'b0;
    end else if(N1609) begin
      mem[1474] <= N1612;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1473] <= 1'b0;
    end else if(N1609) begin
      mem[1473] <= N1611;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1472] <= 1'b0;
    end else if(N1609) begin
      mem[1472] <= N1610;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1471] <= 1'b0;
    end else if(N1543) begin
      mem[1471] <= N1607;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1470] <= 1'b0;
    end else if(N1543) begin
      mem[1470] <= N1606;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1469] <= 1'b0;
    end else if(N1543) begin
      mem[1469] <= N1605;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1468] <= 1'b0;
    end else if(N1543) begin
      mem[1468] <= N1604;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1467] <= 1'b0;
    end else if(N1543) begin
      mem[1467] <= N1603;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1466] <= 1'b0;
    end else if(N1543) begin
      mem[1466] <= N1602;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1465] <= 1'b0;
    end else if(N1543) begin
      mem[1465] <= N1601;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1464] <= 1'b0;
    end else if(N1543) begin
      mem[1464] <= N1600;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1463] <= 1'b0;
    end else if(N1543) begin
      mem[1463] <= N1599;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1462] <= 1'b0;
    end else if(N1543) begin
      mem[1462] <= N1598;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1461] <= 1'b0;
    end else if(N1543) begin
      mem[1461] <= N1597;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1460] <= 1'b0;
    end else if(N1543) begin
      mem[1460] <= N1596;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1459] <= 1'b0;
    end else if(N1543) begin
      mem[1459] <= N1595;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1458] <= 1'b0;
    end else if(N1543) begin
      mem[1458] <= N1594;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1457] <= 1'b0;
    end else if(N1543) begin
      mem[1457] <= N1593;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1456] <= 1'b0;
    end else if(N1543) begin
      mem[1456] <= N1592;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1455] <= 1'b0;
    end else if(N1543) begin
      mem[1455] <= N1591;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1454] <= 1'b0;
    end else if(N1543) begin
      mem[1454] <= N1590;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1453] <= 1'b0;
    end else if(N1543) begin
      mem[1453] <= N1589;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1452] <= 1'b0;
    end else if(N1543) begin
      mem[1452] <= N1588;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1451] <= 1'b0;
    end else if(N1543) begin
      mem[1451] <= N1587;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1450] <= 1'b0;
    end else if(N1543) begin
      mem[1450] <= N1586;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1449] <= 1'b0;
    end else if(N1543) begin
      mem[1449] <= N1585;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1448] <= 1'b0;
    end else if(N1543) begin
      mem[1448] <= N1584;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1447] <= 1'b0;
    end else if(N1543) begin
      mem[1447] <= N1583;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1446] <= 1'b0;
    end else if(N1543) begin
      mem[1446] <= N1582;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1445] <= 1'b0;
    end else if(N1543) begin
      mem[1445] <= N1581;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1444] <= 1'b0;
    end else if(N1543) begin
      mem[1444] <= N1580;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1443] <= 1'b0;
    end else if(N1543) begin
      mem[1443] <= N1579;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1442] <= 1'b0;
    end else if(N1543) begin
      mem[1442] <= N1578;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1441] <= 1'b0;
    end else if(N1543) begin
      mem[1441] <= N1577;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1440] <= 1'b0;
    end else if(N1543) begin
      mem[1440] <= N1576;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1439] <= 1'b0;
    end else if(N1543) begin
      mem[1439] <= N1575;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1438] <= 1'b0;
    end else if(N1543) begin
      mem[1438] <= N1574;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1437] <= 1'b0;
    end else if(N1543) begin
      mem[1437] <= N1573;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1436] <= 1'b0;
    end else if(N1543) begin
      mem[1436] <= N1572;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1435] <= 1'b0;
    end else if(N1543) begin
      mem[1435] <= N1571;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1434] <= 1'b0;
    end else if(N1543) begin
      mem[1434] <= N1570;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1433] <= 1'b0;
    end else if(N1543) begin
      mem[1433] <= N1569;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1432] <= 1'b0;
    end else if(N1543) begin
      mem[1432] <= N1568;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1431] <= 1'b0;
    end else if(N1543) begin
      mem[1431] <= N1567;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1430] <= 1'b0;
    end else if(N1543) begin
      mem[1430] <= N1566;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1429] <= 1'b0;
    end else if(N1543) begin
      mem[1429] <= N1565;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1428] <= 1'b0;
    end else if(N1543) begin
      mem[1428] <= N1564;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1427] <= 1'b0;
    end else if(N1543) begin
      mem[1427] <= N1563;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1426] <= 1'b0;
    end else if(N1543) begin
      mem[1426] <= N1562;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1425] <= 1'b0;
    end else if(N1543) begin
      mem[1425] <= N1561;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1424] <= 1'b0;
    end else if(N1543) begin
      mem[1424] <= N1560;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1423] <= 1'b0;
    end else if(N1543) begin
      mem[1423] <= N1559;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1422] <= 1'b0;
    end else if(N1543) begin
      mem[1422] <= N1558;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1421] <= 1'b0;
    end else if(N1543) begin
      mem[1421] <= N1557;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1420] <= 1'b0;
    end else if(N1543) begin
      mem[1420] <= N1556;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1419] <= 1'b0;
    end else if(N1543) begin
      mem[1419] <= N1555;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1418] <= 1'b0;
    end else if(N1543) begin
      mem[1418] <= N1554;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1417] <= 1'b0;
    end else if(N1543) begin
      mem[1417] <= N1553;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1416] <= 1'b0;
    end else if(N1543) begin
      mem[1416] <= N1552;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1415] <= 1'b0;
    end else if(N1543) begin
      mem[1415] <= N1551;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1414] <= 1'b0;
    end else if(N1543) begin
      mem[1414] <= N1550;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1413] <= 1'b0;
    end else if(N1543) begin
      mem[1413] <= N1549;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1412] <= 1'b0;
    end else if(N1543) begin
      mem[1412] <= N1548;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1411] <= 1'b0;
    end else if(N1543) begin
      mem[1411] <= N1547;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1410] <= 1'b0;
    end else if(N1543) begin
      mem[1410] <= N1546;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1409] <= 1'b0;
    end else if(N1543) begin
      mem[1409] <= N1545;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1408] <= 1'b0;
    end else if(N1543) begin
      mem[1408] <= N1544;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1407] <= 1'b0;
    end else if(N1477) begin
      mem[1407] <= N1541;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1406] <= 1'b0;
    end else if(N1477) begin
      mem[1406] <= N1540;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1405] <= 1'b0;
    end else if(N1477) begin
      mem[1405] <= N1539;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1404] <= 1'b0;
    end else if(N1477) begin
      mem[1404] <= N1538;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1403] <= 1'b0;
    end else if(N1477) begin
      mem[1403] <= N1537;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1402] <= 1'b0;
    end else if(N1477) begin
      mem[1402] <= N1536;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1401] <= 1'b0;
    end else if(N1477) begin
      mem[1401] <= N1535;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1400] <= 1'b0;
    end else if(N1477) begin
      mem[1400] <= N1534;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1399] <= 1'b0;
    end else if(N1477) begin
      mem[1399] <= N1533;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1398] <= 1'b0;
    end else if(N1477) begin
      mem[1398] <= N1532;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1397] <= 1'b0;
    end else if(N1477) begin
      mem[1397] <= N1531;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1396] <= 1'b0;
    end else if(N1477) begin
      mem[1396] <= N1530;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1395] <= 1'b0;
    end else if(N1477) begin
      mem[1395] <= N1529;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1394] <= 1'b0;
    end else if(N1477) begin
      mem[1394] <= N1528;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1393] <= 1'b0;
    end else if(N1477) begin
      mem[1393] <= N1527;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1392] <= 1'b0;
    end else if(N1477) begin
      mem[1392] <= N1526;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1391] <= 1'b0;
    end else if(N1477) begin
      mem[1391] <= N1525;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1390] <= 1'b0;
    end else if(N1477) begin
      mem[1390] <= N1524;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1389] <= 1'b0;
    end else if(N1477) begin
      mem[1389] <= N1523;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1388] <= 1'b0;
    end else if(N1477) begin
      mem[1388] <= N1522;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1387] <= 1'b0;
    end else if(N1477) begin
      mem[1387] <= N1521;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1386] <= 1'b0;
    end else if(N1477) begin
      mem[1386] <= N1520;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1385] <= 1'b0;
    end else if(N1477) begin
      mem[1385] <= N1519;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1384] <= 1'b0;
    end else if(N1477) begin
      mem[1384] <= N1518;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1383] <= 1'b0;
    end else if(N1477) begin
      mem[1383] <= N1517;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1382] <= 1'b0;
    end else if(N1477) begin
      mem[1382] <= N1516;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1381] <= 1'b0;
    end else if(N1477) begin
      mem[1381] <= N1515;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1380] <= 1'b0;
    end else if(N1477) begin
      mem[1380] <= N1514;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1379] <= 1'b0;
    end else if(N1477) begin
      mem[1379] <= N1513;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1378] <= 1'b0;
    end else if(N1477) begin
      mem[1378] <= N1512;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1377] <= 1'b0;
    end else if(N1477) begin
      mem[1377] <= N1511;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1376] <= 1'b0;
    end else if(N1477) begin
      mem[1376] <= N1510;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1375] <= 1'b0;
    end else if(N1477) begin
      mem[1375] <= N1509;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1374] <= 1'b0;
    end else if(N1477) begin
      mem[1374] <= N1508;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1373] <= 1'b0;
    end else if(N1477) begin
      mem[1373] <= N1507;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1372] <= 1'b0;
    end else if(N1477) begin
      mem[1372] <= N1506;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1371] <= 1'b0;
    end else if(N1477) begin
      mem[1371] <= N1505;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1370] <= 1'b0;
    end else if(N1477) begin
      mem[1370] <= N1504;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1369] <= 1'b0;
    end else if(N1477) begin
      mem[1369] <= N1503;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1368] <= 1'b0;
    end else if(N1477) begin
      mem[1368] <= N1502;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1367] <= 1'b0;
    end else if(N1477) begin
      mem[1367] <= N1501;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1366] <= 1'b0;
    end else if(N1477) begin
      mem[1366] <= N1500;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1365] <= 1'b0;
    end else if(N1477) begin
      mem[1365] <= N1499;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1364] <= 1'b0;
    end else if(N1477) begin
      mem[1364] <= N1498;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1363] <= 1'b0;
    end else if(N1477) begin
      mem[1363] <= N1497;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1362] <= 1'b0;
    end else if(N1477) begin
      mem[1362] <= N1496;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1361] <= 1'b0;
    end else if(N1477) begin
      mem[1361] <= N1495;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1360] <= 1'b0;
    end else if(N1477) begin
      mem[1360] <= N1494;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1359] <= 1'b0;
    end else if(N1477) begin
      mem[1359] <= N1493;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1358] <= 1'b0;
    end else if(N1477) begin
      mem[1358] <= N1492;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1357] <= 1'b0;
    end else if(N1477) begin
      mem[1357] <= N1491;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1356] <= 1'b0;
    end else if(N1477) begin
      mem[1356] <= N1490;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1355] <= 1'b0;
    end else if(N1477) begin
      mem[1355] <= N1489;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1354] <= 1'b0;
    end else if(N1477) begin
      mem[1354] <= N1488;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1353] <= 1'b0;
    end else if(N1477) begin
      mem[1353] <= N1487;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1352] <= 1'b0;
    end else if(N1477) begin
      mem[1352] <= N1486;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1351] <= 1'b0;
    end else if(N1477) begin
      mem[1351] <= N1485;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1350] <= 1'b0;
    end else if(N1477) begin
      mem[1350] <= N1484;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1349] <= 1'b0;
    end else if(N1477) begin
      mem[1349] <= N1483;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1348] <= 1'b0;
    end else if(N1477) begin
      mem[1348] <= N1482;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1347] <= 1'b0;
    end else if(N1477) begin
      mem[1347] <= N1481;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1346] <= 1'b0;
    end else if(N1477) begin
      mem[1346] <= N1480;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1345] <= 1'b0;
    end else if(N1477) begin
      mem[1345] <= N1479;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1344] <= 1'b0;
    end else if(N1477) begin
      mem[1344] <= N1478;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1343] <= 1'b0;
    end else if(N1411) begin
      mem[1343] <= N1475;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1342] <= 1'b0;
    end else if(N1411) begin
      mem[1342] <= N1474;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1341] <= 1'b0;
    end else if(N1411) begin
      mem[1341] <= N1473;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1340] <= 1'b0;
    end else if(N1411) begin
      mem[1340] <= N1472;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1339] <= 1'b0;
    end else if(N1411) begin
      mem[1339] <= N1471;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1338] <= 1'b0;
    end else if(N1411) begin
      mem[1338] <= N1470;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1337] <= 1'b0;
    end else if(N1411) begin
      mem[1337] <= N1469;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1336] <= 1'b0;
    end else if(N1411) begin
      mem[1336] <= N1468;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1335] <= 1'b0;
    end else if(N1411) begin
      mem[1335] <= N1467;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1334] <= 1'b0;
    end else if(N1411) begin
      mem[1334] <= N1466;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1333] <= 1'b0;
    end else if(N1411) begin
      mem[1333] <= N1465;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1332] <= 1'b0;
    end else if(N1411) begin
      mem[1332] <= N1464;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1331] <= 1'b0;
    end else if(N1411) begin
      mem[1331] <= N1463;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1330] <= 1'b0;
    end else if(N1411) begin
      mem[1330] <= N1462;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1329] <= 1'b0;
    end else if(N1411) begin
      mem[1329] <= N1461;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1328] <= 1'b0;
    end else if(N1411) begin
      mem[1328] <= N1460;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1327] <= 1'b0;
    end else if(N1411) begin
      mem[1327] <= N1459;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1326] <= 1'b0;
    end else if(N1411) begin
      mem[1326] <= N1458;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1325] <= 1'b0;
    end else if(N1411) begin
      mem[1325] <= N1457;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1324] <= 1'b0;
    end else if(N1411) begin
      mem[1324] <= N1456;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1323] <= 1'b0;
    end else if(N1411) begin
      mem[1323] <= N1455;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1322] <= 1'b0;
    end else if(N1411) begin
      mem[1322] <= N1454;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1321] <= 1'b0;
    end else if(N1411) begin
      mem[1321] <= N1453;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1320] <= 1'b0;
    end else if(N1411) begin
      mem[1320] <= N1452;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1319] <= 1'b0;
    end else if(N1411) begin
      mem[1319] <= N1451;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1318] <= 1'b0;
    end else if(N1411) begin
      mem[1318] <= N1450;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1317] <= 1'b0;
    end else if(N1411) begin
      mem[1317] <= N1449;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1316] <= 1'b0;
    end else if(N1411) begin
      mem[1316] <= N1448;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1315] <= 1'b0;
    end else if(N1411) begin
      mem[1315] <= N1447;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1314] <= 1'b0;
    end else if(N1411) begin
      mem[1314] <= N1446;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1313] <= 1'b0;
    end else if(N1411) begin
      mem[1313] <= N1445;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1312] <= 1'b0;
    end else if(N1411) begin
      mem[1312] <= N1444;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1311] <= 1'b0;
    end else if(N1411) begin
      mem[1311] <= N1443;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1310] <= 1'b0;
    end else if(N1411) begin
      mem[1310] <= N1442;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1309] <= 1'b0;
    end else if(N1411) begin
      mem[1309] <= N1441;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1308] <= 1'b0;
    end else if(N1411) begin
      mem[1308] <= N1440;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1307] <= 1'b0;
    end else if(N1411) begin
      mem[1307] <= N1439;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1306] <= 1'b0;
    end else if(N1411) begin
      mem[1306] <= N1438;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1305] <= 1'b0;
    end else if(N1411) begin
      mem[1305] <= N1437;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1304] <= 1'b0;
    end else if(N1411) begin
      mem[1304] <= N1436;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1303] <= 1'b0;
    end else if(N1411) begin
      mem[1303] <= N1435;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1302] <= 1'b0;
    end else if(N1411) begin
      mem[1302] <= N1434;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1301] <= 1'b0;
    end else if(N1411) begin
      mem[1301] <= N1433;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1300] <= 1'b0;
    end else if(N1411) begin
      mem[1300] <= N1432;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1299] <= 1'b0;
    end else if(N1411) begin
      mem[1299] <= N1431;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1298] <= 1'b0;
    end else if(N1411) begin
      mem[1298] <= N1430;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1297] <= 1'b0;
    end else if(N1411) begin
      mem[1297] <= N1429;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1296] <= 1'b0;
    end else if(N1411) begin
      mem[1296] <= N1428;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1295] <= 1'b0;
    end else if(N1411) begin
      mem[1295] <= N1427;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1294] <= 1'b0;
    end else if(N1411) begin
      mem[1294] <= N1426;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1293] <= 1'b0;
    end else if(N1411) begin
      mem[1293] <= N1425;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1292] <= 1'b0;
    end else if(N1411) begin
      mem[1292] <= N1424;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1291] <= 1'b0;
    end else if(N1411) begin
      mem[1291] <= N1423;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1290] <= 1'b0;
    end else if(N1411) begin
      mem[1290] <= N1422;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1289] <= 1'b0;
    end else if(N1411) begin
      mem[1289] <= N1421;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1288] <= 1'b0;
    end else if(N1411) begin
      mem[1288] <= N1420;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1287] <= 1'b0;
    end else if(N1411) begin
      mem[1287] <= N1419;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1286] <= 1'b0;
    end else if(N1411) begin
      mem[1286] <= N1418;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1285] <= 1'b0;
    end else if(N1411) begin
      mem[1285] <= N1417;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1284] <= 1'b0;
    end else if(N1411) begin
      mem[1284] <= N1416;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1283] <= 1'b0;
    end else if(N1411) begin
      mem[1283] <= N1415;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1282] <= 1'b0;
    end else if(N1411) begin
      mem[1282] <= N1414;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1281] <= 1'b0;
    end else if(N1411) begin
      mem[1281] <= N1413;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1280] <= 1'b0;
    end else if(N1411) begin
      mem[1280] <= N1412;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1279] <= 1'b0;
    end else if(N1345) begin
      mem[1279] <= N1409;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1278] <= 1'b0;
    end else if(N1345) begin
      mem[1278] <= N1408;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1277] <= 1'b0;
    end else if(N1345) begin
      mem[1277] <= N1407;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1276] <= 1'b0;
    end else if(N1345) begin
      mem[1276] <= N1406;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1275] <= 1'b0;
    end else if(N1345) begin
      mem[1275] <= N1405;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1274] <= 1'b0;
    end else if(N1345) begin
      mem[1274] <= N1404;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1273] <= 1'b0;
    end else if(N1345) begin
      mem[1273] <= N1403;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1272] <= 1'b0;
    end else if(N1345) begin
      mem[1272] <= N1402;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1271] <= 1'b0;
    end else if(N1345) begin
      mem[1271] <= N1401;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1270] <= 1'b0;
    end else if(N1345) begin
      mem[1270] <= N1400;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1269] <= 1'b0;
    end else if(N1345) begin
      mem[1269] <= N1399;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1268] <= 1'b0;
    end else if(N1345) begin
      mem[1268] <= N1398;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1267] <= 1'b0;
    end else if(N1345) begin
      mem[1267] <= N1397;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1266] <= 1'b0;
    end else if(N1345) begin
      mem[1266] <= N1396;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1265] <= 1'b0;
    end else if(N1345) begin
      mem[1265] <= N1395;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1264] <= 1'b0;
    end else if(N1345) begin
      mem[1264] <= N1394;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1263] <= 1'b0;
    end else if(N1345) begin
      mem[1263] <= N1393;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1262] <= 1'b0;
    end else if(N1345) begin
      mem[1262] <= N1392;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1261] <= 1'b0;
    end else if(N1345) begin
      mem[1261] <= N1391;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1260] <= 1'b0;
    end else if(N1345) begin
      mem[1260] <= N1390;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1259] <= 1'b0;
    end else if(N1345) begin
      mem[1259] <= N1389;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1258] <= 1'b0;
    end else if(N1345) begin
      mem[1258] <= N1388;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1257] <= 1'b0;
    end else if(N1345) begin
      mem[1257] <= N1387;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1256] <= 1'b0;
    end else if(N1345) begin
      mem[1256] <= N1386;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1255] <= 1'b0;
    end else if(N1345) begin
      mem[1255] <= N1385;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1254] <= 1'b0;
    end else if(N1345) begin
      mem[1254] <= N1384;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1253] <= 1'b0;
    end else if(N1345) begin
      mem[1253] <= N1383;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1252] <= 1'b0;
    end else if(N1345) begin
      mem[1252] <= N1382;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1251] <= 1'b0;
    end else if(N1345) begin
      mem[1251] <= N1381;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1250] <= 1'b0;
    end else if(N1345) begin
      mem[1250] <= N1380;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1249] <= 1'b0;
    end else if(N1345) begin
      mem[1249] <= N1379;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1248] <= 1'b0;
    end else if(N1345) begin
      mem[1248] <= N1378;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1247] <= 1'b0;
    end else if(N1345) begin
      mem[1247] <= N1377;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1246] <= 1'b0;
    end else if(N1345) begin
      mem[1246] <= N1376;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1245] <= 1'b0;
    end else if(N1345) begin
      mem[1245] <= N1375;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1244] <= 1'b0;
    end else if(N1345) begin
      mem[1244] <= N1374;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1243] <= 1'b0;
    end else if(N1345) begin
      mem[1243] <= N1373;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1242] <= 1'b0;
    end else if(N1345) begin
      mem[1242] <= N1372;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1241] <= 1'b0;
    end else if(N1345) begin
      mem[1241] <= N1371;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1240] <= 1'b0;
    end else if(N1345) begin
      mem[1240] <= N1370;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1239] <= 1'b0;
    end else if(N1345) begin
      mem[1239] <= N1369;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1238] <= 1'b0;
    end else if(N1345) begin
      mem[1238] <= N1368;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1237] <= 1'b0;
    end else if(N1345) begin
      mem[1237] <= N1367;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1236] <= 1'b0;
    end else if(N1345) begin
      mem[1236] <= N1366;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1235] <= 1'b0;
    end else if(N1345) begin
      mem[1235] <= N1365;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1234] <= 1'b0;
    end else if(N1345) begin
      mem[1234] <= N1364;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1233] <= 1'b0;
    end else if(N1345) begin
      mem[1233] <= N1363;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1232] <= 1'b0;
    end else if(N1345) begin
      mem[1232] <= N1362;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1231] <= 1'b0;
    end else if(N1345) begin
      mem[1231] <= N1361;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1230] <= 1'b0;
    end else if(N1345) begin
      mem[1230] <= N1360;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1229] <= 1'b0;
    end else if(N1345) begin
      mem[1229] <= N1359;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1228] <= 1'b0;
    end else if(N1345) begin
      mem[1228] <= N1358;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1227] <= 1'b0;
    end else if(N1345) begin
      mem[1227] <= N1357;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1226] <= 1'b0;
    end else if(N1345) begin
      mem[1226] <= N1356;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1225] <= 1'b0;
    end else if(N1345) begin
      mem[1225] <= N1355;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1224] <= 1'b0;
    end else if(N1345) begin
      mem[1224] <= N1354;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1223] <= 1'b0;
    end else if(N1345) begin
      mem[1223] <= N1353;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1222] <= 1'b0;
    end else if(N1345) begin
      mem[1222] <= N1352;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1221] <= 1'b0;
    end else if(N1345) begin
      mem[1221] <= N1351;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1220] <= 1'b0;
    end else if(N1345) begin
      mem[1220] <= N1350;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1219] <= 1'b0;
    end else if(N1345) begin
      mem[1219] <= N1349;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1218] <= 1'b0;
    end else if(N1345) begin
      mem[1218] <= N1348;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1217] <= 1'b0;
    end else if(N1345) begin
      mem[1217] <= N1347;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1216] <= 1'b0;
    end else if(N1345) begin
      mem[1216] <= N1346;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1215] <= 1'b0;
    end else if(N1279) begin
      mem[1215] <= N1343;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1214] <= 1'b0;
    end else if(N1279) begin
      mem[1214] <= N1342;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1213] <= 1'b0;
    end else if(N1279) begin
      mem[1213] <= N1341;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1212] <= 1'b0;
    end else if(N1279) begin
      mem[1212] <= N1340;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1211] <= 1'b0;
    end else if(N1279) begin
      mem[1211] <= N1339;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1210] <= 1'b0;
    end else if(N1279) begin
      mem[1210] <= N1338;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1209] <= 1'b0;
    end else if(N1279) begin
      mem[1209] <= N1337;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1208] <= 1'b0;
    end else if(N1279) begin
      mem[1208] <= N1336;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1207] <= 1'b0;
    end else if(N1279) begin
      mem[1207] <= N1335;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1206] <= 1'b0;
    end else if(N1279) begin
      mem[1206] <= N1334;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1205] <= 1'b0;
    end else if(N1279) begin
      mem[1205] <= N1333;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1204] <= 1'b0;
    end else if(N1279) begin
      mem[1204] <= N1332;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1203] <= 1'b0;
    end else if(N1279) begin
      mem[1203] <= N1331;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1202] <= 1'b0;
    end else if(N1279) begin
      mem[1202] <= N1330;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1201] <= 1'b0;
    end else if(N1279) begin
      mem[1201] <= N1329;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1200] <= 1'b0;
    end else if(N1279) begin
      mem[1200] <= N1328;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1199] <= 1'b0;
    end else if(N1279) begin
      mem[1199] <= N1327;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1198] <= 1'b0;
    end else if(N1279) begin
      mem[1198] <= N1326;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1197] <= 1'b0;
    end else if(N1279) begin
      mem[1197] <= N1325;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1196] <= 1'b0;
    end else if(N1279) begin
      mem[1196] <= N1324;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1195] <= 1'b0;
    end else if(N1279) begin
      mem[1195] <= N1323;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1194] <= 1'b0;
    end else if(N1279) begin
      mem[1194] <= N1322;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1193] <= 1'b0;
    end else if(N1279) begin
      mem[1193] <= N1321;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1192] <= 1'b0;
    end else if(N1279) begin
      mem[1192] <= N1320;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1191] <= 1'b0;
    end else if(N1279) begin
      mem[1191] <= N1319;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1190] <= 1'b0;
    end else if(N1279) begin
      mem[1190] <= N1318;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1189] <= 1'b0;
    end else if(N1279) begin
      mem[1189] <= N1317;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1188] <= 1'b0;
    end else if(N1279) begin
      mem[1188] <= N1316;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1187] <= 1'b0;
    end else if(N1279) begin
      mem[1187] <= N1315;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1186] <= 1'b0;
    end else if(N1279) begin
      mem[1186] <= N1314;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1185] <= 1'b0;
    end else if(N1279) begin
      mem[1185] <= N1313;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1184] <= 1'b0;
    end else if(N1279) begin
      mem[1184] <= N1312;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1183] <= 1'b0;
    end else if(N1279) begin
      mem[1183] <= N1311;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1182] <= 1'b0;
    end else if(N1279) begin
      mem[1182] <= N1310;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1181] <= 1'b0;
    end else if(N1279) begin
      mem[1181] <= N1309;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1180] <= 1'b0;
    end else if(N1279) begin
      mem[1180] <= N1308;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1179] <= 1'b0;
    end else if(N1279) begin
      mem[1179] <= N1307;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1178] <= 1'b0;
    end else if(N1279) begin
      mem[1178] <= N1306;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1177] <= 1'b0;
    end else if(N1279) begin
      mem[1177] <= N1305;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1176] <= 1'b0;
    end else if(N1279) begin
      mem[1176] <= N1304;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1175] <= 1'b0;
    end else if(N1279) begin
      mem[1175] <= N1303;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1174] <= 1'b0;
    end else if(N1279) begin
      mem[1174] <= N1302;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1173] <= 1'b0;
    end else if(N1279) begin
      mem[1173] <= N1301;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1172] <= 1'b0;
    end else if(N1279) begin
      mem[1172] <= N1300;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1171] <= 1'b0;
    end else if(N1279) begin
      mem[1171] <= N1299;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1170] <= 1'b0;
    end else if(N1279) begin
      mem[1170] <= N1298;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1169] <= 1'b0;
    end else if(N1279) begin
      mem[1169] <= N1297;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1168] <= 1'b0;
    end else if(N1279) begin
      mem[1168] <= N1296;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1167] <= 1'b0;
    end else if(N1279) begin
      mem[1167] <= N1295;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1166] <= 1'b0;
    end else if(N1279) begin
      mem[1166] <= N1294;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1165] <= 1'b0;
    end else if(N1279) begin
      mem[1165] <= N1293;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1164] <= 1'b0;
    end else if(N1279) begin
      mem[1164] <= N1292;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1163] <= 1'b0;
    end else if(N1279) begin
      mem[1163] <= N1291;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1162] <= 1'b0;
    end else if(N1279) begin
      mem[1162] <= N1290;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1161] <= 1'b0;
    end else if(N1279) begin
      mem[1161] <= N1289;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1160] <= 1'b0;
    end else if(N1279) begin
      mem[1160] <= N1288;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1159] <= 1'b0;
    end else if(N1279) begin
      mem[1159] <= N1287;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1158] <= 1'b0;
    end else if(N1279) begin
      mem[1158] <= N1286;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1157] <= 1'b0;
    end else if(N1279) begin
      mem[1157] <= N1285;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1156] <= 1'b0;
    end else if(N1279) begin
      mem[1156] <= N1284;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1155] <= 1'b0;
    end else if(N1279) begin
      mem[1155] <= N1283;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1154] <= 1'b0;
    end else if(N1279) begin
      mem[1154] <= N1282;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1153] <= 1'b0;
    end else if(N1279) begin
      mem[1153] <= N1281;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1152] <= 1'b0;
    end else if(N1279) begin
      mem[1152] <= N1280;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1151] <= 1'b0;
    end else if(N1213) begin
      mem[1151] <= N1277;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1150] <= 1'b0;
    end else if(N1213) begin
      mem[1150] <= N1276;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1149] <= 1'b0;
    end else if(N1213) begin
      mem[1149] <= N1275;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1148] <= 1'b0;
    end else if(N1213) begin
      mem[1148] <= N1274;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1147] <= 1'b0;
    end else if(N1213) begin
      mem[1147] <= N1273;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1146] <= 1'b0;
    end else if(N1213) begin
      mem[1146] <= N1272;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1145] <= 1'b0;
    end else if(N1213) begin
      mem[1145] <= N1271;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1144] <= 1'b0;
    end else if(N1213) begin
      mem[1144] <= N1270;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1143] <= 1'b0;
    end else if(N1213) begin
      mem[1143] <= N1269;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1142] <= 1'b0;
    end else if(N1213) begin
      mem[1142] <= N1268;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1141] <= 1'b0;
    end else if(N1213) begin
      mem[1141] <= N1267;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1140] <= 1'b0;
    end else if(N1213) begin
      mem[1140] <= N1266;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1139] <= 1'b0;
    end else if(N1213) begin
      mem[1139] <= N1265;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1138] <= 1'b0;
    end else if(N1213) begin
      mem[1138] <= N1264;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1137] <= 1'b0;
    end else if(N1213) begin
      mem[1137] <= N1263;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1136] <= 1'b0;
    end else if(N1213) begin
      mem[1136] <= N1262;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1135] <= 1'b0;
    end else if(N1213) begin
      mem[1135] <= N1261;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1134] <= 1'b0;
    end else if(N1213) begin
      mem[1134] <= N1260;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1133] <= 1'b0;
    end else if(N1213) begin
      mem[1133] <= N1259;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1132] <= 1'b0;
    end else if(N1213) begin
      mem[1132] <= N1258;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1131] <= 1'b0;
    end else if(N1213) begin
      mem[1131] <= N1257;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1130] <= 1'b0;
    end else if(N1213) begin
      mem[1130] <= N1256;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1129] <= 1'b0;
    end else if(N1213) begin
      mem[1129] <= N1255;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1128] <= 1'b0;
    end else if(N1213) begin
      mem[1128] <= N1254;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1127] <= 1'b0;
    end else if(N1213) begin
      mem[1127] <= N1253;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1126] <= 1'b0;
    end else if(N1213) begin
      mem[1126] <= N1252;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1125] <= 1'b0;
    end else if(N1213) begin
      mem[1125] <= N1251;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1124] <= 1'b0;
    end else if(N1213) begin
      mem[1124] <= N1250;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1123] <= 1'b0;
    end else if(N1213) begin
      mem[1123] <= N1249;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1122] <= 1'b0;
    end else if(N1213) begin
      mem[1122] <= N1248;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1121] <= 1'b0;
    end else if(N1213) begin
      mem[1121] <= N1247;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1120] <= 1'b0;
    end else if(N1213) begin
      mem[1120] <= N1246;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1119] <= 1'b0;
    end else if(N1213) begin
      mem[1119] <= N1245;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1118] <= 1'b0;
    end else if(N1213) begin
      mem[1118] <= N1244;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1117] <= 1'b0;
    end else if(N1213) begin
      mem[1117] <= N1243;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1116] <= 1'b0;
    end else if(N1213) begin
      mem[1116] <= N1242;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1115] <= 1'b0;
    end else if(N1213) begin
      mem[1115] <= N1241;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1114] <= 1'b0;
    end else if(N1213) begin
      mem[1114] <= N1240;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1113] <= 1'b0;
    end else if(N1213) begin
      mem[1113] <= N1239;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1112] <= 1'b0;
    end else if(N1213) begin
      mem[1112] <= N1238;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1111] <= 1'b0;
    end else if(N1213) begin
      mem[1111] <= N1237;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1110] <= 1'b0;
    end else if(N1213) begin
      mem[1110] <= N1236;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1109] <= 1'b0;
    end else if(N1213) begin
      mem[1109] <= N1235;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1108] <= 1'b0;
    end else if(N1213) begin
      mem[1108] <= N1234;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1107] <= 1'b0;
    end else if(N1213) begin
      mem[1107] <= N1233;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1106] <= 1'b0;
    end else if(N1213) begin
      mem[1106] <= N1232;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1105] <= 1'b0;
    end else if(N1213) begin
      mem[1105] <= N1231;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1104] <= 1'b0;
    end else if(N1213) begin
      mem[1104] <= N1230;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1103] <= 1'b0;
    end else if(N1213) begin
      mem[1103] <= N1229;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1102] <= 1'b0;
    end else if(N1213) begin
      mem[1102] <= N1228;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1101] <= 1'b0;
    end else if(N1213) begin
      mem[1101] <= N1227;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1100] <= 1'b0;
    end else if(N1213) begin
      mem[1100] <= N1226;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1099] <= 1'b0;
    end else if(N1213) begin
      mem[1099] <= N1225;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1098] <= 1'b0;
    end else if(N1213) begin
      mem[1098] <= N1224;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1097] <= 1'b0;
    end else if(N1213) begin
      mem[1097] <= N1223;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1096] <= 1'b0;
    end else if(N1213) begin
      mem[1096] <= N1222;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1095] <= 1'b0;
    end else if(N1213) begin
      mem[1095] <= N1221;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1094] <= 1'b0;
    end else if(N1213) begin
      mem[1094] <= N1220;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1093] <= 1'b0;
    end else if(N1213) begin
      mem[1093] <= N1219;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1092] <= 1'b0;
    end else if(N1213) begin
      mem[1092] <= N1218;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1091] <= 1'b0;
    end else if(N1213) begin
      mem[1091] <= N1217;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1090] <= 1'b0;
    end else if(N1213) begin
      mem[1090] <= N1216;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1089] <= 1'b0;
    end else if(N1213) begin
      mem[1089] <= N1215;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1088] <= 1'b0;
    end else if(N1213) begin
      mem[1088] <= N1214;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1087] <= 1'b0;
    end else if(N1147) begin
      mem[1087] <= N1211;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1086] <= 1'b0;
    end else if(N1147) begin
      mem[1086] <= N1210;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1085] <= 1'b0;
    end else if(N1147) begin
      mem[1085] <= N1209;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1084] <= 1'b0;
    end else if(N1147) begin
      mem[1084] <= N1208;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1083] <= 1'b0;
    end else if(N1147) begin
      mem[1083] <= N1207;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1082] <= 1'b0;
    end else if(N1147) begin
      mem[1082] <= N1206;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1081] <= 1'b0;
    end else if(N1147) begin
      mem[1081] <= N1205;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1080] <= 1'b0;
    end else if(N1147) begin
      mem[1080] <= N1204;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1079] <= 1'b0;
    end else if(N1147) begin
      mem[1079] <= N1203;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1078] <= 1'b0;
    end else if(N1147) begin
      mem[1078] <= N1202;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1077] <= 1'b0;
    end else if(N1147) begin
      mem[1077] <= N1201;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1076] <= 1'b0;
    end else if(N1147) begin
      mem[1076] <= N1200;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1075] <= 1'b0;
    end else if(N1147) begin
      mem[1075] <= N1199;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1074] <= 1'b0;
    end else if(N1147) begin
      mem[1074] <= N1198;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1073] <= 1'b0;
    end else if(N1147) begin
      mem[1073] <= N1197;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1072] <= 1'b0;
    end else if(N1147) begin
      mem[1072] <= N1196;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1071] <= 1'b0;
    end else if(N1147) begin
      mem[1071] <= N1195;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1070] <= 1'b0;
    end else if(N1147) begin
      mem[1070] <= N1194;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1069] <= 1'b0;
    end else if(N1147) begin
      mem[1069] <= N1193;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1068] <= 1'b0;
    end else if(N1147) begin
      mem[1068] <= N1192;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1067] <= 1'b0;
    end else if(N1147) begin
      mem[1067] <= N1191;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1066] <= 1'b0;
    end else if(N1147) begin
      mem[1066] <= N1190;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1065] <= 1'b0;
    end else if(N1147) begin
      mem[1065] <= N1189;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1064] <= 1'b0;
    end else if(N1147) begin
      mem[1064] <= N1188;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1063] <= 1'b0;
    end else if(N1147) begin
      mem[1063] <= N1187;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1062] <= 1'b0;
    end else if(N1147) begin
      mem[1062] <= N1186;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1061] <= 1'b0;
    end else if(N1147) begin
      mem[1061] <= N1185;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1060] <= 1'b0;
    end else if(N1147) begin
      mem[1060] <= N1184;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1059] <= 1'b0;
    end else if(N1147) begin
      mem[1059] <= N1183;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1058] <= 1'b0;
    end else if(N1147) begin
      mem[1058] <= N1182;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1057] <= 1'b0;
    end else if(N1147) begin
      mem[1057] <= N1181;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1056] <= 1'b0;
    end else if(N1147) begin
      mem[1056] <= N1180;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1055] <= 1'b0;
    end else if(N1147) begin
      mem[1055] <= N1179;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1054] <= 1'b0;
    end else if(N1147) begin
      mem[1054] <= N1178;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1053] <= 1'b0;
    end else if(N1147) begin
      mem[1053] <= N1177;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1052] <= 1'b0;
    end else if(N1147) begin
      mem[1052] <= N1176;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1051] <= 1'b0;
    end else if(N1147) begin
      mem[1051] <= N1175;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1050] <= 1'b0;
    end else if(N1147) begin
      mem[1050] <= N1174;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1049] <= 1'b0;
    end else if(N1147) begin
      mem[1049] <= N1173;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1048] <= 1'b0;
    end else if(N1147) begin
      mem[1048] <= N1172;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1047] <= 1'b0;
    end else if(N1147) begin
      mem[1047] <= N1171;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1046] <= 1'b0;
    end else if(N1147) begin
      mem[1046] <= N1170;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1045] <= 1'b0;
    end else if(N1147) begin
      mem[1045] <= N1169;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1044] <= 1'b0;
    end else if(N1147) begin
      mem[1044] <= N1168;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1043] <= 1'b0;
    end else if(N1147) begin
      mem[1043] <= N1167;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1042] <= 1'b0;
    end else if(N1147) begin
      mem[1042] <= N1166;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1041] <= 1'b0;
    end else if(N1147) begin
      mem[1041] <= N1165;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1040] <= 1'b0;
    end else if(N1147) begin
      mem[1040] <= N1164;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1039] <= 1'b0;
    end else if(N1147) begin
      mem[1039] <= N1163;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1038] <= 1'b0;
    end else if(N1147) begin
      mem[1038] <= N1162;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1037] <= 1'b0;
    end else if(N1147) begin
      mem[1037] <= N1161;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1036] <= 1'b0;
    end else if(N1147) begin
      mem[1036] <= N1160;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1035] <= 1'b0;
    end else if(N1147) begin
      mem[1035] <= N1159;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1034] <= 1'b0;
    end else if(N1147) begin
      mem[1034] <= N1158;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1033] <= 1'b0;
    end else if(N1147) begin
      mem[1033] <= N1157;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1032] <= 1'b0;
    end else if(N1147) begin
      mem[1032] <= N1156;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1031] <= 1'b0;
    end else if(N1147) begin
      mem[1031] <= N1155;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1030] <= 1'b0;
    end else if(N1147) begin
      mem[1030] <= N1154;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1029] <= 1'b0;
    end else if(N1147) begin
      mem[1029] <= N1153;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1028] <= 1'b0;
    end else if(N1147) begin
      mem[1028] <= N1152;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1027] <= 1'b0;
    end else if(N1147) begin
      mem[1027] <= N1151;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1026] <= 1'b0;
    end else if(N1147) begin
      mem[1026] <= N1150;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1025] <= 1'b0;
    end else if(N1147) begin
      mem[1025] <= N1149;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1024] <= 1'b0;
    end else if(N1147) begin
      mem[1024] <= N1148;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1023] <= 1'b0;
    end else if(N1081) begin
      mem[1023] <= N1145;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1022] <= 1'b0;
    end else if(N1081) begin
      mem[1022] <= N1144;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1021] <= 1'b0;
    end else if(N1081) begin
      mem[1021] <= N1143;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1020] <= 1'b0;
    end else if(N1081) begin
      mem[1020] <= N1142;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1019] <= 1'b0;
    end else if(N1081) begin
      mem[1019] <= N1141;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1018] <= 1'b0;
    end else if(N1081) begin
      mem[1018] <= N1140;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1017] <= 1'b0;
    end else if(N1081) begin
      mem[1017] <= N1139;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1016] <= 1'b0;
    end else if(N1081) begin
      mem[1016] <= N1138;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1015] <= 1'b0;
    end else if(N1081) begin
      mem[1015] <= N1137;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1014] <= 1'b0;
    end else if(N1081) begin
      mem[1014] <= N1136;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1013] <= 1'b0;
    end else if(N1081) begin
      mem[1013] <= N1135;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1012] <= 1'b0;
    end else if(N1081) begin
      mem[1012] <= N1134;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1011] <= 1'b0;
    end else if(N1081) begin
      mem[1011] <= N1133;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1010] <= 1'b0;
    end else if(N1081) begin
      mem[1010] <= N1132;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1009] <= 1'b0;
    end else if(N1081) begin
      mem[1009] <= N1131;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1008] <= 1'b0;
    end else if(N1081) begin
      mem[1008] <= N1130;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1007] <= 1'b0;
    end else if(N1081) begin
      mem[1007] <= N1129;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1006] <= 1'b0;
    end else if(N1081) begin
      mem[1006] <= N1128;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1005] <= 1'b0;
    end else if(N1081) begin
      mem[1005] <= N1127;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1004] <= 1'b0;
    end else if(N1081) begin
      mem[1004] <= N1126;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1003] <= 1'b0;
    end else if(N1081) begin
      mem[1003] <= N1125;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1002] <= 1'b0;
    end else if(N1081) begin
      mem[1002] <= N1124;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1001] <= 1'b0;
    end else if(N1081) begin
      mem[1001] <= N1123;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1000] <= 1'b0;
    end else if(N1081) begin
      mem[1000] <= N1122;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[999] <= 1'b0;
    end else if(N1081) begin
      mem[999] <= N1121;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[998] <= 1'b0;
    end else if(N1081) begin
      mem[998] <= N1120;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[997] <= 1'b0;
    end else if(N1081) begin
      mem[997] <= N1119;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[996] <= 1'b0;
    end else if(N1081) begin
      mem[996] <= N1118;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[995] <= 1'b0;
    end else if(N1081) begin
      mem[995] <= N1117;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[994] <= 1'b0;
    end else if(N1081) begin
      mem[994] <= N1116;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[993] <= 1'b0;
    end else if(N1081) begin
      mem[993] <= N1115;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[992] <= 1'b0;
    end else if(N1081) begin
      mem[992] <= N1114;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[991] <= 1'b0;
    end else if(N1081) begin
      mem[991] <= N1113;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[990] <= 1'b0;
    end else if(N1081) begin
      mem[990] <= N1112;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[989] <= 1'b0;
    end else if(N1081) begin
      mem[989] <= N1111;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[988] <= 1'b0;
    end else if(N1081) begin
      mem[988] <= N1110;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[987] <= 1'b0;
    end else if(N1081) begin
      mem[987] <= N1109;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[986] <= 1'b0;
    end else if(N1081) begin
      mem[986] <= N1108;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[985] <= 1'b0;
    end else if(N1081) begin
      mem[985] <= N1107;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[984] <= 1'b0;
    end else if(N1081) begin
      mem[984] <= N1106;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[983] <= 1'b0;
    end else if(N1081) begin
      mem[983] <= N1105;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[982] <= 1'b0;
    end else if(N1081) begin
      mem[982] <= N1104;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[981] <= 1'b0;
    end else if(N1081) begin
      mem[981] <= N1103;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[980] <= 1'b0;
    end else if(N1081) begin
      mem[980] <= N1102;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[979] <= 1'b0;
    end else if(N1081) begin
      mem[979] <= N1101;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[978] <= 1'b0;
    end else if(N1081) begin
      mem[978] <= N1100;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[977] <= 1'b0;
    end else if(N1081) begin
      mem[977] <= N1099;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[976] <= 1'b0;
    end else if(N1081) begin
      mem[976] <= N1098;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[975] <= 1'b0;
    end else if(N1081) begin
      mem[975] <= N1097;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[974] <= 1'b0;
    end else if(N1081) begin
      mem[974] <= N1096;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[973] <= 1'b0;
    end else if(N1081) begin
      mem[973] <= N1095;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[972] <= 1'b0;
    end else if(N1081) begin
      mem[972] <= N1094;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[971] <= 1'b0;
    end else if(N1081) begin
      mem[971] <= N1093;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[970] <= 1'b0;
    end else if(N1081) begin
      mem[970] <= N1092;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[969] <= 1'b0;
    end else if(N1081) begin
      mem[969] <= N1091;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[968] <= 1'b0;
    end else if(N1081) begin
      mem[968] <= N1090;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[967] <= 1'b0;
    end else if(N1081) begin
      mem[967] <= N1089;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[966] <= 1'b0;
    end else if(N1081) begin
      mem[966] <= N1088;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[965] <= 1'b0;
    end else if(N1081) begin
      mem[965] <= N1087;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[964] <= 1'b0;
    end else if(N1081) begin
      mem[964] <= N1086;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[963] <= 1'b0;
    end else if(N1081) begin
      mem[963] <= N1085;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[962] <= 1'b0;
    end else if(N1081) begin
      mem[962] <= N1084;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[961] <= 1'b0;
    end else if(N1081) begin
      mem[961] <= N1083;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[960] <= 1'b0;
    end else if(N1081) begin
      mem[960] <= N1082;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[959] <= 1'b0;
    end else if(N1015) begin
      mem[959] <= N1079;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[958] <= 1'b0;
    end else if(N1015) begin
      mem[958] <= N1078;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[957] <= 1'b0;
    end else if(N1015) begin
      mem[957] <= N1077;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[956] <= 1'b0;
    end else if(N1015) begin
      mem[956] <= N1076;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[955] <= 1'b0;
    end else if(N1015) begin
      mem[955] <= N1075;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[954] <= 1'b0;
    end else if(N1015) begin
      mem[954] <= N1074;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[953] <= 1'b0;
    end else if(N1015) begin
      mem[953] <= N1073;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[952] <= 1'b0;
    end else if(N1015) begin
      mem[952] <= N1072;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[951] <= 1'b0;
    end else if(N1015) begin
      mem[951] <= N1071;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[950] <= 1'b0;
    end else if(N1015) begin
      mem[950] <= N1070;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[949] <= 1'b0;
    end else if(N1015) begin
      mem[949] <= N1069;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[948] <= 1'b0;
    end else if(N1015) begin
      mem[948] <= N1068;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[947] <= 1'b0;
    end else if(N1015) begin
      mem[947] <= N1067;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[946] <= 1'b0;
    end else if(N1015) begin
      mem[946] <= N1066;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[945] <= 1'b0;
    end else if(N1015) begin
      mem[945] <= N1065;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[944] <= 1'b0;
    end else if(N1015) begin
      mem[944] <= N1064;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[943] <= 1'b0;
    end else if(N1015) begin
      mem[943] <= N1063;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[942] <= 1'b0;
    end else if(N1015) begin
      mem[942] <= N1062;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[941] <= 1'b0;
    end else if(N1015) begin
      mem[941] <= N1061;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[940] <= 1'b0;
    end else if(N1015) begin
      mem[940] <= N1060;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[939] <= 1'b0;
    end else if(N1015) begin
      mem[939] <= N1059;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[938] <= 1'b0;
    end else if(N1015) begin
      mem[938] <= N1058;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[937] <= 1'b0;
    end else if(N1015) begin
      mem[937] <= N1057;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[936] <= 1'b0;
    end else if(N1015) begin
      mem[936] <= N1056;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[935] <= 1'b0;
    end else if(N1015) begin
      mem[935] <= N1055;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[934] <= 1'b0;
    end else if(N1015) begin
      mem[934] <= N1054;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[933] <= 1'b0;
    end else if(N1015) begin
      mem[933] <= N1053;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[932] <= 1'b0;
    end else if(N1015) begin
      mem[932] <= N1052;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[931] <= 1'b0;
    end else if(N1015) begin
      mem[931] <= N1051;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[930] <= 1'b0;
    end else if(N1015) begin
      mem[930] <= N1050;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[929] <= 1'b0;
    end else if(N1015) begin
      mem[929] <= N1049;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[928] <= 1'b0;
    end else if(N1015) begin
      mem[928] <= N1048;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[927] <= 1'b0;
    end else if(N1015) begin
      mem[927] <= N1047;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[926] <= 1'b0;
    end else if(N1015) begin
      mem[926] <= N1046;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[925] <= 1'b0;
    end else if(N1015) begin
      mem[925] <= N1045;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[924] <= 1'b0;
    end else if(N1015) begin
      mem[924] <= N1044;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[923] <= 1'b0;
    end else if(N1015) begin
      mem[923] <= N1043;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[922] <= 1'b0;
    end else if(N1015) begin
      mem[922] <= N1042;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[921] <= 1'b0;
    end else if(N1015) begin
      mem[921] <= N1041;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[920] <= 1'b0;
    end else if(N1015) begin
      mem[920] <= N1040;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[919] <= 1'b0;
    end else if(N1015) begin
      mem[919] <= N1039;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[918] <= 1'b0;
    end else if(N1015) begin
      mem[918] <= N1038;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[917] <= 1'b0;
    end else if(N1015) begin
      mem[917] <= N1037;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[916] <= 1'b0;
    end else if(N1015) begin
      mem[916] <= N1036;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[915] <= 1'b0;
    end else if(N1015) begin
      mem[915] <= N1035;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[914] <= 1'b0;
    end else if(N1015) begin
      mem[914] <= N1034;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[913] <= 1'b0;
    end else if(N1015) begin
      mem[913] <= N1033;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[912] <= 1'b0;
    end else if(N1015) begin
      mem[912] <= N1032;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[911] <= 1'b0;
    end else if(N1015) begin
      mem[911] <= N1031;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[910] <= 1'b0;
    end else if(N1015) begin
      mem[910] <= N1030;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[909] <= 1'b0;
    end else if(N1015) begin
      mem[909] <= N1029;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[908] <= 1'b0;
    end else if(N1015) begin
      mem[908] <= N1028;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[907] <= 1'b0;
    end else if(N1015) begin
      mem[907] <= N1027;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[906] <= 1'b0;
    end else if(N1015) begin
      mem[906] <= N1026;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[905] <= 1'b0;
    end else if(N1015) begin
      mem[905] <= N1025;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[904] <= 1'b0;
    end else if(N1015) begin
      mem[904] <= N1024;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[903] <= 1'b0;
    end else if(N1015) begin
      mem[903] <= N1023;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[902] <= 1'b0;
    end else if(N1015) begin
      mem[902] <= N1022;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[901] <= 1'b0;
    end else if(N1015) begin
      mem[901] <= N1021;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[900] <= 1'b0;
    end else if(N1015) begin
      mem[900] <= N1020;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[899] <= 1'b0;
    end else if(N1015) begin
      mem[899] <= N1019;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[898] <= 1'b0;
    end else if(N1015) begin
      mem[898] <= N1018;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[897] <= 1'b0;
    end else if(N1015) begin
      mem[897] <= N1017;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[896] <= 1'b0;
    end else if(N1015) begin
      mem[896] <= N1016;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[895] <= 1'b0;
    end else if(N949) begin
      mem[895] <= N1013;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[894] <= 1'b0;
    end else if(N949) begin
      mem[894] <= N1012;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[893] <= 1'b0;
    end else if(N949) begin
      mem[893] <= N1011;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[892] <= 1'b0;
    end else if(N949) begin
      mem[892] <= N1010;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[891] <= 1'b0;
    end else if(N949) begin
      mem[891] <= N1009;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[890] <= 1'b0;
    end else if(N949) begin
      mem[890] <= N1008;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[889] <= 1'b0;
    end else if(N949) begin
      mem[889] <= N1007;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[888] <= 1'b0;
    end else if(N949) begin
      mem[888] <= N1006;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[887] <= 1'b0;
    end else if(N949) begin
      mem[887] <= N1005;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[886] <= 1'b0;
    end else if(N949) begin
      mem[886] <= N1004;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[885] <= 1'b0;
    end else if(N949) begin
      mem[885] <= N1003;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[884] <= 1'b0;
    end else if(N949) begin
      mem[884] <= N1002;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[883] <= 1'b0;
    end else if(N949) begin
      mem[883] <= N1001;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[882] <= 1'b0;
    end else if(N949) begin
      mem[882] <= N1000;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[881] <= 1'b0;
    end else if(N949) begin
      mem[881] <= N999;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[880] <= 1'b0;
    end else if(N949) begin
      mem[880] <= N998;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[879] <= 1'b0;
    end else if(N949) begin
      mem[879] <= N997;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[878] <= 1'b0;
    end else if(N949) begin
      mem[878] <= N996;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[877] <= 1'b0;
    end else if(N949) begin
      mem[877] <= N995;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[876] <= 1'b0;
    end else if(N949) begin
      mem[876] <= N994;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[875] <= 1'b0;
    end else if(N949) begin
      mem[875] <= N993;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[874] <= 1'b0;
    end else if(N949) begin
      mem[874] <= N992;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[873] <= 1'b0;
    end else if(N949) begin
      mem[873] <= N991;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[872] <= 1'b0;
    end else if(N949) begin
      mem[872] <= N990;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[871] <= 1'b0;
    end else if(N949) begin
      mem[871] <= N989;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[870] <= 1'b0;
    end else if(N949) begin
      mem[870] <= N988;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[869] <= 1'b0;
    end else if(N949) begin
      mem[869] <= N987;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[868] <= 1'b0;
    end else if(N949) begin
      mem[868] <= N986;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[867] <= 1'b0;
    end else if(N949) begin
      mem[867] <= N985;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[866] <= 1'b0;
    end else if(N949) begin
      mem[866] <= N984;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[865] <= 1'b0;
    end else if(N949) begin
      mem[865] <= N983;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[864] <= 1'b0;
    end else if(N949) begin
      mem[864] <= N982;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[863] <= 1'b0;
    end else if(N949) begin
      mem[863] <= N981;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[862] <= 1'b0;
    end else if(N949) begin
      mem[862] <= N980;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[861] <= 1'b0;
    end else if(N949) begin
      mem[861] <= N979;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[860] <= 1'b0;
    end else if(N949) begin
      mem[860] <= N978;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[859] <= 1'b0;
    end else if(N949) begin
      mem[859] <= N977;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[858] <= 1'b0;
    end else if(N949) begin
      mem[858] <= N976;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[857] <= 1'b0;
    end else if(N949) begin
      mem[857] <= N975;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[856] <= 1'b0;
    end else if(N949) begin
      mem[856] <= N974;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[855] <= 1'b0;
    end else if(N949) begin
      mem[855] <= N973;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[854] <= 1'b0;
    end else if(N949) begin
      mem[854] <= N972;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[853] <= 1'b0;
    end else if(N949) begin
      mem[853] <= N971;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[852] <= 1'b0;
    end else if(N949) begin
      mem[852] <= N970;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[851] <= 1'b0;
    end else if(N949) begin
      mem[851] <= N969;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[850] <= 1'b0;
    end else if(N949) begin
      mem[850] <= N968;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[849] <= 1'b0;
    end else if(N949) begin
      mem[849] <= N967;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[848] <= 1'b0;
    end else if(N949) begin
      mem[848] <= N966;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[847] <= 1'b0;
    end else if(N949) begin
      mem[847] <= N965;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[846] <= 1'b0;
    end else if(N949) begin
      mem[846] <= N964;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[845] <= 1'b0;
    end else if(N949) begin
      mem[845] <= N963;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[844] <= 1'b0;
    end else if(N949) begin
      mem[844] <= N962;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[843] <= 1'b0;
    end else if(N949) begin
      mem[843] <= N961;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[842] <= 1'b0;
    end else if(N949) begin
      mem[842] <= N960;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[841] <= 1'b0;
    end else if(N949) begin
      mem[841] <= N959;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[840] <= 1'b0;
    end else if(N949) begin
      mem[840] <= N958;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[839] <= 1'b0;
    end else if(N949) begin
      mem[839] <= N957;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[838] <= 1'b0;
    end else if(N949) begin
      mem[838] <= N956;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[837] <= 1'b0;
    end else if(N949) begin
      mem[837] <= N955;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[836] <= 1'b0;
    end else if(N949) begin
      mem[836] <= N954;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[835] <= 1'b0;
    end else if(N949) begin
      mem[835] <= N953;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[834] <= 1'b0;
    end else if(N949) begin
      mem[834] <= N952;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[833] <= 1'b0;
    end else if(N949) begin
      mem[833] <= N951;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[832] <= 1'b0;
    end else if(N949) begin
      mem[832] <= N950;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[831] <= 1'b0;
    end else if(N883) begin
      mem[831] <= N947;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[830] <= 1'b0;
    end else if(N883) begin
      mem[830] <= N946;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[829] <= 1'b0;
    end else if(N883) begin
      mem[829] <= N945;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[828] <= 1'b0;
    end else if(N883) begin
      mem[828] <= N944;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[827] <= 1'b0;
    end else if(N883) begin
      mem[827] <= N943;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[826] <= 1'b0;
    end else if(N883) begin
      mem[826] <= N942;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[825] <= 1'b0;
    end else if(N883) begin
      mem[825] <= N941;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[824] <= 1'b0;
    end else if(N883) begin
      mem[824] <= N940;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[823] <= 1'b0;
    end else if(N883) begin
      mem[823] <= N939;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[822] <= 1'b0;
    end else if(N883) begin
      mem[822] <= N938;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[821] <= 1'b0;
    end else if(N883) begin
      mem[821] <= N937;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[820] <= 1'b0;
    end else if(N883) begin
      mem[820] <= N936;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[819] <= 1'b0;
    end else if(N883) begin
      mem[819] <= N935;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[818] <= 1'b0;
    end else if(N883) begin
      mem[818] <= N934;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[817] <= 1'b0;
    end else if(N883) begin
      mem[817] <= N933;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[816] <= 1'b0;
    end else if(N883) begin
      mem[816] <= N932;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[815] <= 1'b0;
    end else if(N883) begin
      mem[815] <= N931;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[814] <= 1'b0;
    end else if(N883) begin
      mem[814] <= N930;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[813] <= 1'b0;
    end else if(N883) begin
      mem[813] <= N929;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[812] <= 1'b0;
    end else if(N883) begin
      mem[812] <= N928;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[811] <= 1'b0;
    end else if(N883) begin
      mem[811] <= N927;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[810] <= 1'b0;
    end else if(N883) begin
      mem[810] <= N926;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[809] <= 1'b0;
    end else if(N883) begin
      mem[809] <= N925;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[808] <= 1'b0;
    end else if(N883) begin
      mem[808] <= N924;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[807] <= 1'b0;
    end else if(N883) begin
      mem[807] <= N923;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[806] <= 1'b0;
    end else if(N883) begin
      mem[806] <= N922;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[805] <= 1'b0;
    end else if(N883) begin
      mem[805] <= N921;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[804] <= 1'b0;
    end else if(N883) begin
      mem[804] <= N920;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[803] <= 1'b0;
    end else if(N883) begin
      mem[803] <= N919;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[802] <= 1'b0;
    end else if(N883) begin
      mem[802] <= N918;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[801] <= 1'b0;
    end else if(N883) begin
      mem[801] <= N917;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[800] <= 1'b0;
    end else if(N883) begin
      mem[800] <= N916;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[799] <= 1'b0;
    end else if(N883) begin
      mem[799] <= N915;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[798] <= 1'b0;
    end else if(N883) begin
      mem[798] <= N914;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[797] <= 1'b0;
    end else if(N883) begin
      mem[797] <= N913;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[796] <= 1'b0;
    end else if(N883) begin
      mem[796] <= N912;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[795] <= 1'b0;
    end else if(N883) begin
      mem[795] <= N911;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[794] <= 1'b0;
    end else if(N883) begin
      mem[794] <= N910;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[793] <= 1'b0;
    end else if(N883) begin
      mem[793] <= N909;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[792] <= 1'b0;
    end else if(N883) begin
      mem[792] <= N908;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[791] <= 1'b0;
    end else if(N883) begin
      mem[791] <= N907;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[790] <= 1'b0;
    end else if(N883) begin
      mem[790] <= N906;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[789] <= 1'b0;
    end else if(N883) begin
      mem[789] <= N905;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[788] <= 1'b0;
    end else if(N883) begin
      mem[788] <= N904;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[787] <= 1'b0;
    end else if(N883) begin
      mem[787] <= N903;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[786] <= 1'b0;
    end else if(N883) begin
      mem[786] <= N902;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[785] <= 1'b0;
    end else if(N883) begin
      mem[785] <= N901;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[784] <= 1'b0;
    end else if(N883) begin
      mem[784] <= N900;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[783] <= 1'b0;
    end else if(N883) begin
      mem[783] <= N899;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[782] <= 1'b0;
    end else if(N883) begin
      mem[782] <= N898;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[781] <= 1'b0;
    end else if(N883) begin
      mem[781] <= N897;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[780] <= 1'b0;
    end else if(N883) begin
      mem[780] <= N896;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[779] <= 1'b0;
    end else if(N883) begin
      mem[779] <= N895;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[778] <= 1'b0;
    end else if(N883) begin
      mem[778] <= N894;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[777] <= 1'b0;
    end else if(N883) begin
      mem[777] <= N893;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[776] <= 1'b0;
    end else if(N883) begin
      mem[776] <= N892;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[775] <= 1'b0;
    end else if(N883) begin
      mem[775] <= N891;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[774] <= 1'b0;
    end else if(N883) begin
      mem[774] <= N890;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[773] <= 1'b0;
    end else if(N883) begin
      mem[773] <= N889;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[772] <= 1'b0;
    end else if(N883) begin
      mem[772] <= N888;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[771] <= 1'b0;
    end else if(N883) begin
      mem[771] <= N887;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[770] <= 1'b0;
    end else if(N883) begin
      mem[770] <= N886;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[769] <= 1'b0;
    end else if(N883) begin
      mem[769] <= N885;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[768] <= 1'b0;
    end else if(N883) begin
      mem[768] <= N884;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[767] <= 1'b0;
    end else if(N817) begin
      mem[767] <= N881;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[766] <= 1'b0;
    end else if(N817) begin
      mem[766] <= N880;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[765] <= 1'b0;
    end else if(N817) begin
      mem[765] <= N879;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[764] <= 1'b0;
    end else if(N817) begin
      mem[764] <= N878;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[763] <= 1'b0;
    end else if(N817) begin
      mem[763] <= N877;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[762] <= 1'b0;
    end else if(N817) begin
      mem[762] <= N876;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[761] <= 1'b0;
    end else if(N817) begin
      mem[761] <= N875;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[760] <= 1'b0;
    end else if(N817) begin
      mem[760] <= N874;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[759] <= 1'b0;
    end else if(N817) begin
      mem[759] <= N873;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[758] <= 1'b0;
    end else if(N817) begin
      mem[758] <= N872;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[757] <= 1'b0;
    end else if(N817) begin
      mem[757] <= N871;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[756] <= 1'b0;
    end else if(N817) begin
      mem[756] <= N870;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[755] <= 1'b0;
    end else if(N817) begin
      mem[755] <= N869;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[754] <= 1'b0;
    end else if(N817) begin
      mem[754] <= N868;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[753] <= 1'b0;
    end else if(N817) begin
      mem[753] <= N867;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[752] <= 1'b0;
    end else if(N817) begin
      mem[752] <= N866;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[751] <= 1'b0;
    end else if(N817) begin
      mem[751] <= N865;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[750] <= 1'b0;
    end else if(N817) begin
      mem[750] <= N864;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[749] <= 1'b0;
    end else if(N817) begin
      mem[749] <= N863;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[748] <= 1'b0;
    end else if(N817) begin
      mem[748] <= N862;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[747] <= 1'b0;
    end else if(N817) begin
      mem[747] <= N861;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[746] <= 1'b0;
    end else if(N817) begin
      mem[746] <= N860;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[745] <= 1'b0;
    end else if(N817) begin
      mem[745] <= N859;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[744] <= 1'b0;
    end else if(N817) begin
      mem[744] <= N858;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[743] <= 1'b0;
    end else if(N817) begin
      mem[743] <= N857;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[742] <= 1'b0;
    end else if(N817) begin
      mem[742] <= N856;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[741] <= 1'b0;
    end else if(N817) begin
      mem[741] <= N855;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[740] <= 1'b0;
    end else if(N817) begin
      mem[740] <= N854;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[739] <= 1'b0;
    end else if(N817) begin
      mem[739] <= N853;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[738] <= 1'b0;
    end else if(N817) begin
      mem[738] <= N852;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[737] <= 1'b0;
    end else if(N817) begin
      mem[737] <= N851;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[736] <= 1'b0;
    end else if(N817) begin
      mem[736] <= N850;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[735] <= 1'b0;
    end else if(N817) begin
      mem[735] <= N849;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[734] <= 1'b0;
    end else if(N817) begin
      mem[734] <= N848;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[733] <= 1'b0;
    end else if(N817) begin
      mem[733] <= N847;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[732] <= 1'b0;
    end else if(N817) begin
      mem[732] <= N846;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[731] <= 1'b0;
    end else if(N817) begin
      mem[731] <= N845;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[730] <= 1'b0;
    end else if(N817) begin
      mem[730] <= N844;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[729] <= 1'b0;
    end else if(N817) begin
      mem[729] <= N843;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[728] <= 1'b0;
    end else if(N817) begin
      mem[728] <= N842;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[727] <= 1'b0;
    end else if(N817) begin
      mem[727] <= N841;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[726] <= 1'b0;
    end else if(N817) begin
      mem[726] <= N840;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[725] <= 1'b0;
    end else if(N817) begin
      mem[725] <= N839;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[724] <= 1'b0;
    end else if(N817) begin
      mem[724] <= N838;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[723] <= 1'b0;
    end else if(N817) begin
      mem[723] <= N837;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[722] <= 1'b0;
    end else if(N817) begin
      mem[722] <= N836;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[721] <= 1'b0;
    end else if(N817) begin
      mem[721] <= N835;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[720] <= 1'b0;
    end else if(N817) begin
      mem[720] <= N834;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[719] <= 1'b0;
    end else if(N817) begin
      mem[719] <= N833;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[718] <= 1'b0;
    end else if(N817) begin
      mem[718] <= N832;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[717] <= 1'b0;
    end else if(N817) begin
      mem[717] <= N831;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[716] <= 1'b0;
    end else if(N817) begin
      mem[716] <= N830;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[715] <= 1'b0;
    end else if(N817) begin
      mem[715] <= N829;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[714] <= 1'b0;
    end else if(N817) begin
      mem[714] <= N828;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[713] <= 1'b0;
    end else if(N817) begin
      mem[713] <= N827;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[712] <= 1'b0;
    end else if(N817) begin
      mem[712] <= N826;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[711] <= 1'b0;
    end else if(N817) begin
      mem[711] <= N825;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[710] <= 1'b0;
    end else if(N817) begin
      mem[710] <= N824;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[709] <= 1'b0;
    end else if(N817) begin
      mem[709] <= N823;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[708] <= 1'b0;
    end else if(N817) begin
      mem[708] <= N822;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[707] <= 1'b0;
    end else if(N817) begin
      mem[707] <= N821;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[706] <= 1'b0;
    end else if(N817) begin
      mem[706] <= N820;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[705] <= 1'b0;
    end else if(N817) begin
      mem[705] <= N819;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[704] <= 1'b0;
    end else if(N817) begin
      mem[704] <= N818;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[703] <= 1'b0;
    end else if(N751) begin
      mem[703] <= N815;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[702] <= 1'b0;
    end else if(N751) begin
      mem[702] <= N814;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[701] <= 1'b0;
    end else if(N751) begin
      mem[701] <= N813;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[700] <= 1'b0;
    end else if(N751) begin
      mem[700] <= N812;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[699] <= 1'b0;
    end else if(N751) begin
      mem[699] <= N811;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[698] <= 1'b0;
    end else if(N751) begin
      mem[698] <= N810;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[697] <= 1'b0;
    end else if(N751) begin
      mem[697] <= N809;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[696] <= 1'b0;
    end else if(N751) begin
      mem[696] <= N808;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[695] <= 1'b0;
    end else if(N751) begin
      mem[695] <= N807;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[694] <= 1'b0;
    end else if(N751) begin
      mem[694] <= N806;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[693] <= 1'b0;
    end else if(N751) begin
      mem[693] <= N805;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[692] <= 1'b0;
    end else if(N751) begin
      mem[692] <= N804;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[691] <= 1'b0;
    end else if(N751) begin
      mem[691] <= N803;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[690] <= 1'b0;
    end else if(N751) begin
      mem[690] <= N802;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[689] <= 1'b0;
    end else if(N751) begin
      mem[689] <= N801;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[688] <= 1'b0;
    end else if(N751) begin
      mem[688] <= N800;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[687] <= 1'b0;
    end else if(N751) begin
      mem[687] <= N799;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[686] <= 1'b0;
    end else if(N751) begin
      mem[686] <= N798;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[685] <= 1'b0;
    end else if(N751) begin
      mem[685] <= N797;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[684] <= 1'b0;
    end else if(N751) begin
      mem[684] <= N796;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[683] <= 1'b0;
    end else if(N751) begin
      mem[683] <= N795;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[682] <= 1'b0;
    end else if(N751) begin
      mem[682] <= N794;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[681] <= 1'b0;
    end else if(N751) begin
      mem[681] <= N793;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[680] <= 1'b0;
    end else if(N751) begin
      mem[680] <= N792;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[679] <= 1'b0;
    end else if(N751) begin
      mem[679] <= N791;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[678] <= 1'b0;
    end else if(N751) begin
      mem[678] <= N790;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[677] <= 1'b0;
    end else if(N751) begin
      mem[677] <= N789;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[676] <= 1'b0;
    end else if(N751) begin
      mem[676] <= N788;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[675] <= 1'b0;
    end else if(N751) begin
      mem[675] <= N787;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[674] <= 1'b0;
    end else if(N751) begin
      mem[674] <= N786;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[673] <= 1'b0;
    end else if(N751) begin
      mem[673] <= N785;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[672] <= 1'b0;
    end else if(N751) begin
      mem[672] <= N784;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[671] <= 1'b0;
    end else if(N751) begin
      mem[671] <= N783;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[670] <= 1'b0;
    end else if(N751) begin
      mem[670] <= N782;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[669] <= 1'b0;
    end else if(N751) begin
      mem[669] <= N781;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[668] <= 1'b0;
    end else if(N751) begin
      mem[668] <= N780;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[667] <= 1'b0;
    end else if(N751) begin
      mem[667] <= N779;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[666] <= 1'b0;
    end else if(N751) begin
      mem[666] <= N778;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[665] <= 1'b0;
    end else if(N751) begin
      mem[665] <= N777;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[664] <= 1'b0;
    end else if(N751) begin
      mem[664] <= N776;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[663] <= 1'b0;
    end else if(N751) begin
      mem[663] <= N775;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[662] <= 1'b0;
    end else if(N751) begin
      mem[662] <= N774;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[661] <= 1'b0;
    end else if(N751) begin
      mem[661] <= N773;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[660] <= 1'b0;
    end else if(N751) begin
      mem[660] <= N772;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[659] <= 1'b0;
    end else if(N751) begin
      mem[659] <= N771;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[658] <= 1'b0;
    end else if(N751) begin
      mem[658] <= N770;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[657] <= 1'b0;
    end else if(N751) begin
      mem[657] <= N769;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[656] <= 1'b0;
    end else if(N751) begin
      mem[656] <= N768;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[655] <= 1'b0;
    end else if(N751) begin
      mem[655] <= N767;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[654] <= 1'b0;
    end else if(N751) begin
      mem[654] <= N766;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[653] <= 1'b0;
    end else if(N751) begin
      mem[653] <= N765;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[652] <= 1'b0;
    end else if(N751) begin
      mem[652] <= N764;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[651] <= 1'b0;
    end else if(N751) begin
      mem[651] <= N763;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[650] <= 1'b0;
    end else if(N751) begin
      mem[650] <= N762;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[649] <= 1'b0;
    end else if(N751) begin
      mem[649] <= N761;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[648] <= 1'b0;
    end else if(N751) begin
      mem[648] <= N760;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[647] <= 1'b0;
    end else if(N751) begin
      mem[647] <= N759;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[646] <= 1'b0;
    end else if(N751) begin
      mem[646] <= N758;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[645] <= 1'b0;
    end else if(N751) begin
      mem[645] <= N757;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[644] <= 1'b0;
    end else if(N751) begin
      mem[644] <= N756;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[643] <= 1'b0;
    end else if(N751) begin
      mem[643] <= N755;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[642] <= 1'b0;
    end else if(N751) begin
      mem[642] <= N754;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[641] <= 1'b0;
    end else if(N751) begin
      mem[641] <= N753;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[640] <= 1'b0;
    end else if(N751) begin
      mem[640] <= N752;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[639] <= 1'b0;
    end else if(N685) begin
      mem[639] <= N749;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[638] <= 1'b0;
    end else if(N685) begin
      mem[638] <= N748;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[637] <= 1'b0;
    end else if(N685) begin
      mem[637] <= N747;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[636] <= 1'b0;
    end else if(N685) begin
      mem[636] <= N746;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[635] <= 1'b0;
    end else if(N685) begin
      mem[635] <= N745;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[634] <= 1'b0;
    end else if(N685) begin
      mem[634] <= N744;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[633] <= 1'b0;
    end else if(N685) begin
      mem[633] <= N743;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[632] <= 1'b0;
    end else if(N685) begin
      mem[632] <= N742;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[631] <= 1'b0;
    end else if(N685) begin
      mem[631] <= N741;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[630] <= 1'b0;
    end else if(N685) begin
      mem[630] <= N740;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[629] <= 1'b0;
    end else if(N685) begin
      mem[629] <= N739;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[628] <= 1'b0;
    end else if(N685) begin
      mem[628] <= N738;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[627] <= 1'b0;
    end else if(N685) begin
      mem[627] <= N737;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[626] <= 1'b0;
    end else if(N685) begin
      mem[626] <= N736;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[625] <= 1'b0;
    end else if(N685) begin
      mem[625] <= N735;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[624] <= 1'b0;
    end else if(N685) begin
      mem[624] <= N734;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[623] <= 1'b0;
    end else if(N685) begin
      mem[623] <= N733;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[622] <= 1'b0;
    end else if(N685) begin
      mem[622] <= N732;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[621] <= 1'b0;
    end else if(N685) begin
      mem[621] <= N731;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[620] <= 1'b0;
    end else if(N685) begin
      mem[620] <= N730;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[619] <= 1'b0;
    end else if(N685) begin
      mem[619] <= N729;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[618] <= 1'b0;
    end else if(N685) begin
      mem[618] <= N728;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[617] <= 1'b0;
    end else if(N685) begin
      mem[617] <= N727;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[616] <= 1'b0;
    end else if(N685) begin
      mem[616] <= N726;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[615] <= 1'b0;
    end else if(N685) begin
      mem[615] <= N725;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[614] <= 1'b0;
    end else if(N685) begin
      mem[614] <= N724;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[613] <= 1'b0;
    end else if(N685) begin
      mem[613] <= N723;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[612] <= 1'b0;
    end else if(N685) begin
      mem[612] <= N722;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[611] <= 1'b0;
    end else if(N685) begin
      mem[611] <= N721;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[610] <= 1'b0;
    end else if(N685) begin
      mem[610] <= N720;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[609] <= 1'b0;
    end else if(N685) begin
      mem[609] <= N719;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[608] <= 1'b0;
    end else if(N685) begin
      mem[608] <= N718;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[607] <= 1'b0;
    end else if(N685) begin
      mem[607] <= N717;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[606] <= 1'b0;
    end else if(N685) begin
      mem[606] <= N716;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[605] <= 1'b0;
    end else if(N685) begin
      mem[605] <= N715;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[604] <= 1'b0;
    end else if(N685) begin
      mem[604] <= N714;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[603] <= 1'b0;
    end else if(N685) begin
      mem[603] <= N713;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[602] <= 1'b0;
    end else if(N685) begin
      mem[602] <= N712;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[601] <= 1'b0;
    end else if(N685) begin
      mem[601] <= N711;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[600] <= 1'b0;
    end else if(N685) begin
      mem[600] <= N710;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[599] <= 1'b0;
    end else if(N685) begin
      mem[599] <= N709;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[598] <= 1'b0;
    end else if(N685) begin
      mem[598] <= N708;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[597] <= 1'b0;
    end else if(N685) begin
      mem[597] <= N707;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[596] <= 1'b0;
    end else if(N685) begin
      mem[596] <= N706;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[595] <= 1'b0;
    end else if(N685) begin
      mem[595] <= N705;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[594] <= 1'b0;
    end else if(N685) begin
      mem[594] <= N704;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[593] <= 1'b0;
    end else if(N685) begin
      mem[593] <= N703;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[592] <= 1'b0;
    end else if(N685) begin
      mem[592] <= N702;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[591] <= 1'b0;
    end else if(N685) begin
      mem[591] <= N701;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[590] <= 1'b0;
    end else if(N685) begin
      mem[590] <= N700;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[589] <= 1'b0;
    end else if(N685) begin
      mem[589] <= N699;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[588] <= 1'b0;
    end else if(N685) begin
      mem[588] <= N698;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[587] <= 1'b0;
    end else if(N685) begin
      mem[587] <= N697;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[586] <= 1'b0;
    end else if(N685) begin
      mem[586] <= N696;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[585] <= 1'b0;
    end else if(N685) begin
      mem[585] <= N695;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[584] <= 1'b0;
    end else if(N685) begin
      mem[584] <= N694;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[583] <= 1'b0;
    end else if(N685) begin
      mem[583] <= N693;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[582] <= 1'b0;
    end else if(N685) begin
      mem[582] <= N692;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[581] <= 1'b0;
    end else if(N685) begin
      mem[581] <= N691;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[580] <= 1'b0;
    end else if(N685) begin
      mem[580] <= N690;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[579] <= 1'b0;
    end else if(N685) begin
      mem[579] <= N689;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[578] <= 1'b0;
    end else if(N685) begin
      mem[578] <= N688;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[577] <= 1'b0;
    end else if(N685) begin
      mem[577] <= N687;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[576] <= 1'b0;
    end else if(N685) begin
      mem[576] <= N686;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[575] <= 1'b0;
    end else if(N619) begin
      mem[575] <= N683;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[574] <= 1'b0;
    end else if(N619) begin
      mem[574] <= N682;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[573] <= 1'b0;
    end else if(N619) begin
      mem[573] <= N681;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[572] <= 1'b0;
    end else if(N619) begin
      mem[572] <= N680;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[571] <= 1'b0;
    end else if(N619) begin
      mem[571] <= N679;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[570] <= 1'b0;
    end else if(N619) begin
      mem[570] <= N678;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[569] <= 1'b0;
    end else if(N619) begin
      mem[569] <= N677;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[568] <= 1'b0;
    end else if(N619) begin
      mem[568] <= N676;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[567] <= 1'b0;
    end else if(N619) begin
      mem[567] <= N675;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[566] <= 1'b0;
    end else if(N619) begin
      mem[566] <= N674;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[565] <= 1'b0;
    end else if(N619) begin
      mem[565] <= N673;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[564] <= 1'b0;
    end else if(N619) begin
      mem[564] <= N672;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[563] <= 1'b0;
    end else if(N619) begin
      mem[563] <= N671;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[562] <= 1'b0;
    end else if(N619) begin
      mem[562] <= N670;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[561] <= 1'b0;
    end else if(N619) begin
      mem[561] <= N669;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[560] <= 1'b0;
    end else if(N619) begin
      mem[560] <= N668;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[559] <= 1'b0;
    end else if(N619) begin
      mem[559] <= N667;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[558] <= 1'b0;
    end else if(N619) begin
      mem[558] <= N666;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[557] <= 1'b0;
    end else if(N619) begin
      mem[557] <= N665;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[556] <= 1'b0;
    end else if(N619) begin
      mem[556] <= N664;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[555] <= 1'b0;
    end else if(N619) begin
      mem[555] <= N663;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[554] <= 1'b0;
    end else if(N619) begin
      mem[554] <= N662;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[553] <= 1'b0;
    end else if(N619) begin
      mem[553] <= N661;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[552] <= 1'b0;
    end else if(N619) begin
      mem[552] <= N660;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[551] <= 1'b0;
    end else if(N619) begin
      mem[551] <= N659;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[550] <= 1'b0;
    end else if(N619) begin
      mem[550] <= N658;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[549] <= 1'b0;
    end else if(N619) begin
      mem[549] <= N657;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[548] <= 1'b0;
    end else if(N619) begin
      mem[548] <= N656;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[547] <= 1'b0;
    end else if(N619) begin
      mem[547] <= N655;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[546] <= 1'b0;
    end else if(N619) begin
      mem[546] <= N654;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[545] <= 1'b0;
    end else if(N619) begin
      mem[545] <= N653;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[544] <= 1'b0;
    end else if(N619) begin
      mem[544] <= N652;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[543] <= 1'b0;
    end else if(N619) begin
      mem[543] <= N651;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[542] <= 1'b0;
    end else if(N619) begin
      mem[542] <= N650;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[541] <= 1'b0;
    end else if(N619) begin
      mem[541] <= N649;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[540] <= 1'b0;
    end else if(N619) begin
      mem[540] <= N648;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[539] <= 1'b0;
    end else if(N619) begin
      mem[539] <= N647;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[538] <= 1'b0;
    end else if(N619) begin
      mem[538] <= N646;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[537] <= 1'b0;
    end else if(N619) begin
      mem[537] <= N645;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[536] <= 1'b0;
    end else if(N619) begin
      mem[536] <= N644;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[535] <= 1'b0;
    end else if(N619) begin
      mem[535] <= N643;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[534] <= 1'b0;
    end else if(N619) begin
      mem[534] <= N642;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[533] <= 1'b0;
    end else if(N619) begin
      mem[533] <= N641;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[532] <= 1'b0;
    end else if(N619) begin
      mem[532] <= N640;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[531] <= 1'b0;
    end else if(N619) begin
      mem[531] <= N639;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[530] <= 1'b0;
    end else if(N619) begin
      mem[530] <= N638;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[529] <= 1'b0;
    end else if(N619) begin
      mem[529] <= N637;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[528] <= 1'b0;
    end else if(N619) begin
      mem[528] <= N636;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[527] <= 1'b0;
    end else if(N619) begin
      mem[527] <= N635;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[526] <= 1'b0;
    end else if(N619) begin
      mem[526] <= N634;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[525] <= 1'b0;
    end else if(N619) begin
      mem[525] <= N633;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[524] <= 1'b0;
    end else if(N619) begin
      mem[524] <= N632;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[523] <= 1'b0;
    end else if(N619) begin
      mem[523] <= N631;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[522] <= 1'b0;
    end else if(N619) begin
      mem[522] <= N630;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[521] <= 1'b0;
    end else if(N619) begin
      mem[521] <= N629;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[520] <= 1'b0;
    end else if(N619) begin
      mem[520] <= N628;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[519] <= 1'b0;
    end else if(N619) begin
      mem[519] <= N627;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[518] <= 1'b0;
    end else if(N619) begin
      mem[518] <= N626;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[517] <= 1'b0;
    end else if(N619) begin
      mem[517] <= N625;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[516] <= 1'b0;
    end else if(N619) begin
      mem[516] <= N624;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[515] <= 1'b0;
    end else if(N619) begin
      mem[515] <= N623;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[514] <= 1'b0;
    end else if(N619) begin
      mem[514] <= N622;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[513] <= 1'b0;
    end else if(N619) begin
      mem[513] <= N621;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[512] <= 1'b0;
    end else if(N619) begin
      mem[512] <= N620;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[511] <= 1'b0;
    end else if(N553) begin
      mem[511] <= N617;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[510] <= 1'b0;
    end else if(N553) begin
      mem[510] <= N616;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[509] <= 1'b0;
    end else if(N553) begin
      mem[509] <= N615;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[508] <= 1'b0;
    end else if(N553) begin
      mem[508] <= N614;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[507] <= 1'b0;
    end else if(N553) begin
      mem[507] <= N613;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[506] <= 1'b0;
    end else if(N553) begin
      mem[506] <= N612;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[505] <= 1'b0;
    end else if(N553) begin
      mem[505] <= N611;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[504] <= 1'b0;
    end else if(N553) begin
      mem[504] <= N610;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[503] <= 1'b0;
    end else if(N553) begin
      mem[503] <= N609;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[502] <= 1'b0;
    end else if(N553) begin
      mem[502] <= N608;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[501] <= 1'b0;
    end else if(N553) begin
      mem[501] <= N607;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[500] <= 1'b0;
    end else if(N553) begin
      mem[500] <= N606;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[499] <= 1'b0;
    end else if(N553) begin
      mem[499] <= N605;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[498] <= 1'b0;
    end else if(N553) begin
      mem[498] <= N604;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[497] <= 1'b0;
    end else if(N553) begin
      mem[497] <= N603;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[496] <= 1'b0;
    end else if(N553) begin
      mem[496] <= N602;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[495] <= 1'b0;
    end else if(N553) begin
      mem[495] <= N601;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[494] <= 1'b0;
    end else if(N553) begin
      mem[494] <= N600;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[493] <= 1'b0;
    end else if(N553) begin
      mem[493] <= N599;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[492] <= 1'b0;
    end else if(N553) begin
      mem[492] <= N598;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[491] <= 1'b0;
    end else if(N553) begin
      mem[491] <= N597;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[490] <= 1'b0;
    end else if(N553) begin
      mem[490] <= N596;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[489] <= 1'b0;
    end else if(N553) begin
      mem[489] <= N595;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[488] <= 1'b0;
    end else if(N553) begin
      mem[488] <= N594;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[487] <= 1'b0;
    end else if(N553) begin
      mem[487] <= N593;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[486] <= 1'b0;
    end else if(N553) begin
      mem[486] <= N592;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[485] <= 1'b0;
    end else if(N553) begin
      mem[485] <= N591;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[484] <= 1'b0;
    end else if(N553) begin
      mem[484] <= N590;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[483] <= 1'b0;
    end else if(N553) begin
      mem[483] <= N589;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[482] <= 1'b0;
    end else if(N553) begin
      mem[482] <= N588;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[481] <= 1'b0;
    end else if(N553) begin
      mem[481] <= N587;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[480] <= 1'b0;
    end else if(N553) begin
      mem[480] <= N586;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[479] <= 1'b0;
    end else if(N553) begin
      mem[479] <= N585;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[478] <= 1'b0;
    end else if(N553) begin
      mem[478] <= N584;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[477] <= 1'b0;
    end else if(N553) begin
      mem[477] <= N583;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[476] <= 1'b0;
    end else if(N553) begin
      mem[476] <= N582;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[475] <= 1'b0;
    end else if(N553) begin
      mem[475] <= N581;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[474] <= 1'b0;
    end else if(N553) begin
      mem[474] <= N580;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[473] <= 1'b0;
    end else if(N553) begin
      mem[473] <= N579;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[472] <= 1'b0;
    end else if(N553) begin
      mem[472] <= N578;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[471] <= 1'b0;
    end else if(N553) begin
      mem[471] <= N577;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[470] <= 1'b0;
    end else if(N553) begin
      mem[470] <= N576;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[469] <= 1'b0;
    end else if(N553) begin
      mem[469] <= N575;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[468] <= 1'b0;
    end else if(N553) begin
      mem[468] <= N574;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[467] <= 1'b0;
    end else if(N553) begin
      mem[467] <= N573;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[466] <= 1'b0;
    end else if(N553) begin
      mem[466] <= N572;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[465] <= 1'b0;
    end else if(N553) begin
      mem[465] <= N571;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[464] <= 1'b0;
    end else if(N553) begin
      mem[464] <= N570;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[463] <= 1'b0;
    end else if(N553) begin
      mem[463] <= N569;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[462] <= 1'b0;
    end else if(N553) begin
      mem[462] <= N568;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[461] <= 1'b0;
    end else if(N553) begin
      mem[461] <= N567;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[460] <= 1'b0;
    end else if(N553) begin
      mem[460] <= N566;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[459] <= 1'b0;
    end else if(N553) begin
      mem[459] <= N565;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[458] <= 1'b0;
    end else if(N553) begin
      mem[458] <= N564;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[457] <= 1'b0;
    end else if(N553) begin
      mem[457] <= N563;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[456] <= 1'b0;
    end else if(N553) begin
      mem[456] <= N562;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[455] <= 1'b0;
    end else if(N553) begin
      mem[455] <= N561;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[454] <= 1'b0;
    end else if(N553) begin
      mem[454] <= N560;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[453] <= 1'b0;
    end else if(N553) begin
      mem[453] <= N559;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[452] <= 1'b0;
    end else if(N553) begin
      mem[452] <= N558;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[451] <= 1'b0;
    end else if(N553) begin
      mem[451] <= N557;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[450] <= 1'b0;
    end else if(N553) begin
      mem[450] <= N556;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[449] <= 1'b0;
    end else if(N553) begin
      mem[449] <= N555;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[448] <= 1'b0;
    end else if(N553) begin
      mem[448] <= N554;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[447] <= 1'b0;
    end else if(N487) begin
      mem[447] <= N551;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[446] <= 1'b0;
    end else if(N487) begin
      mem[446] <= N550;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[445] <= 1'b0;
    end else if(N487) begin
      mem[445] <= N549;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[444] <= 1'b0;
    end else if(N487) begin
      mem[444] <= N548;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[443] <= 1'b0;
    end else if(N487) begin
      mem[443] <= N547;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[442] <= 1'b0;
    end else if(N487) begin
      mem[442] <= N546;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[441] <= 1'b0;
    end else if(N487) begin
      mem[441] <= N545;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[440] <= 1'b0;
    end else if(N487) begin
      mem[440] <= N544;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[439] <= 1'b0;
    end else if(N487) begin
      mem[439] <= N543;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[438] <= 1'b0;
    end else if(N487) begin
      mem[438] <= N542;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[437] <= 1'b0;
    end else if(N487) begin
      mem[437] <= N541;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[436] <= 1'b0;
    end else if(N487) begin
      mem[436] <= N540;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[435] <= 1'b0;
    end else if(N487) begin
      mem[435] <= N539;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[434] <= 1'b0;
    end else if(N487) begin
      mem[434] <= N538;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[433] <= 1'b0;
    end else if(N487) begin
      mem[433] <= N537;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[432] <= 1'b0;
    end else if(N487) begin
      mem[432] <= N536;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[431] <= 1'b0;
    end else if(N487) begin
      mem[431] <= N535;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[430] <= 1'b0;
    end else if(N487) begin
      mem[430] <= N534;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[429] <= 1'b0;
    end else if(N487) begin
      mem[429] <= N533;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[428] <= 1'b0;
    end else if(N487) begin
      mem[428] <= N532;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[427] <= 1'b0;
    end else if(N487) begin
      mem[427] <= N531;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[426] <= 1'b0;
    end else if(N487) begin
      mem[426] <= N530;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[425] <= 1'b0;
    end else if(N487) begin
      mem[425] <= N529;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[424] <= 1'b0;
    end else if(N487) begin
      mem[424] <= N528;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[423] <= 1'b0;
    end else if(N487) begin
      mem[423] <= N527;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[422] <= 1'b0;
    end else if(N487) begin
      mem[422] <= N526;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[421] <= 1'b0;
    end else if(N487) begin
      mem[421] <= N525;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[420] <= 1'b0;
    end else if(N487) begin
      mem[420] <= N524;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[419] <= 1'b0;
    end else if(N487) begin
      mem[419] <= N523;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[418] <= 1'b0;
    end else if(N487) begin
      mem[418] <= N522;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[417] <= 1'b0;
    end else if(N487) begin
      mem[417] <= N521;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[416] <= 1'b0;
    end else if(N487) begin
      mem[416] <= N520;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[415] <= 1'b0;
    end else if(N487) begin
      mem[415] <= N519;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[414] <= 1'b0;
    end else if(N487) begin
      mem[414] <= N518;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[413] <= 1'b0;
    end else if(N487) begin
      mem[413] <= N517;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[412] <= 1'b0;
    end else if(N487) begin
      mem[412] <= N516;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[411] <= 1'b0;
    end else if(N487) begin
      mem[411] <= N515;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[410] <= 1'b0;
    end else if(N487) begin
      mem[410] <= N514;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[409] <= 1'b0;
    end else if(N487) begin
      mem[409] <= N513;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[408] <= 1'b0;
    end else if(N487) begin
      mem[408] <= N512;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[407] <= 1'b0;
    end else if(N487) begin
      mem[407] <= N511;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[406] <= 1'b0;
    end else if(N487) begin
      mem[406] <= N510;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[405] <= 1'b0;
    end else if(N487) begin
      mem[405] <= N509;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[404] <= 1'b0;
    end else if(N487) begin
      mem[404] <= N508;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[403] <= 1'b0;
    end else if(N487) begin
      mem[403] <= N507;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[402] <= 1'b0;
    end else if(N487) begin
      mem[402] <= N506;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[401] <= 1'b0;
    end else if(N487) begin
      mem[401] <= N505;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[400] <= 1'b0;
    end else if(N487) begin
      mem[400] <= N504;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[399] <= 1'b0;
    end else if(N487) begin
      mem[399] <= N503;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[398] <= 1'b0;
    end else if(N487) begin
      mem[398] <= N502;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[397] <= 1'b0;
    end else if(N487) begin
      mem[397] <= N501;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[396] <= 1'b0;
    end else if(N487) begin
      mem[396] <= N500;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[395] <= 1'b0;
    end else if(N487) begin
      mem[395] <= N499;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[394] <= 1'b0;
    end else if(N487) begin
      mem[394] <= N498;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[393] <= 1'b0;
    end else if(N487) begin
      mem[393] <= N497;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[392] <= 1'b0;
    end else if(N487) begin
      mem[392] <= N496;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[391] <= 1'b0;
    end else if(N487) begin
      mem[391] <= N495;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[390] <= 1'b0;
    end else if(N487) begin
      mem[390] <= N494;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[389] <= 1'b0;
    end else if(N487) begin
      mem[389] <= N493;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[388] <= 1'b0;
    end else if(N487) begin
      mem[388] <= N492;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[387] <= 1'b0;
    end else if(N487) begin
      mem[387] <= N491;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[386] <= 1'b0;
    end else if(N487) begin
      mem[386] <= N490;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[385] <= 1'b0;
    end else if(N487) begin
      mem[385] <= N489;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[384] <= 1'b0;
    end else if(N487) begin
      mem[384] <= N488;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[383] <= 1'b0;
    end else if(N421) begin
      mem[383] <= N485;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[382] <= 1'b0;
    end else if(N421) begin
      mem[382] <= N484;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[381] <= 1'b0;
    end else if(N421) begin
      mem[381] <= N483;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[380] <= 1'b0;
    end else if(N421) begin
      mem[380] <= N482;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[379] <= 1'b0;
    end else if(N421) begin
      mem[379] <= N481;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[378] <= 1'b0;
    end else if(N421) begin
      mem[378] <= N480;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[377] <= 1'b0;
    end else if(N421) begin
      mem[377] <= N479;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[376] <= 1'b0;
    end else if(N421) begin
      mem[376] <= N478;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[375] <= 1'b0;
    end else if(N421) begin
      mem[375] <= N477;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[374] <= 1'b0;
    end else if(N421) begin
      mem[374] <= N476;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[373] <= 1'b0;
    end else if(N421) begin
      mem[373] <= N475;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[372] <= 1'b0;
    end else if(N421) begin
      mem[372] <= N474;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[371] <= 1'b0;
    end else if(N421) begin
      mem[371] <= N473;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[370] <= 1'b0;
    end else if(N421) begin
      mem[370] <= N472;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[369] <= 1'b0;
    end else if(N421) begin
      mem[369] <= N471;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[368] <= 1'b0;
    end else if(N421) begin
      mem[368] <= N470;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[367] <= 1'b0;
    end else if(N421) begin
      mem[367] <= N469;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[366] <= 1'b0;
    end else if(N421) begin
      mem[366] <= N468;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[365] <= 1'b0;
    end else if(N421) begin
      mem[365] <= N467;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[364] <= 1'b0;
    end else if(N421) begin
      mem[364] <= N466;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[363] <= 1'b0;
    end else if(N421) begin
      mem[363] <= N465;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[362] <= 1'b0;
    end else if(N421) begin
      mem[362] <= N464;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[361] <= 1'b0;
    end else if(N421) begin
      mem[361] <= N463;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[360] <= 1'b0;
    end else if(N421) begin
      mem[360] <= N462;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[359] <= 1'b0;
    end else if(N421) begin
      mem[359] <= N461;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[358] <= 1'b0;
    end else if(N421) begin
      mem[358] <= N460;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[357] <= 1'b0;
    end else if(N421) begin
      mem[357] <= N459;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[356] <= 1'b0;
    end else if(N421) begin
      mem[356] <= N458;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[355] <= 1'b0;
    end else if(N421) begin
      mem[355] <= N457;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[354] <= 1'b0;
    end else if(N421) begin
      mem[354] <= N456;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[353] <= 1'b0;
    end else if(N421) begin
      mem[353] <= N455;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[352] <= 1'b0;
    end else if(N421) begin
      mem[352] <= N454;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[351] <= 1'b0;
    end else if(N421) begin
      mem[351] <= N453;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[350] <= 1'b0;
    end else if(N421) begin
      mem[350] <= N452;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[349] <= 1'b0;
    end else if(N421) begin
      mem[349] <= N451;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[348] <= 1'b0;
    end else if(N421) begin
      mem[348] <= N450;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[347] <= 1'b0;
    end else if(N421) begin
      mem[347] <= N449;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[346] <= 1'b0;
    end else if(N421) begin
      mem[346] <= N448;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[345] <= 1'b0;
    end else if(N421) begin
      mem[345] <= N447;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[344] <= 1'b0;
    end else if(N421) begin
      mem[344] <= N446;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[343] <= 1'b0;
    end else if(N421) begin
      mem[343] <= N445;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[342] <= 1'b0;
    end else if(N421) begin
      mem[342] <= N444;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[341] <= 1'b0;
    end else if(N421) begin
      mem[341] <= N443;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[340] <= 1'b0;
    end else if(N421) begin
      mem[340] <= N442;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[339] <= 1'b0;
    end else if(N421) begin
      mem[339] <= N441;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[338] <= 1'b0;
    end else if(N421) begin
      mem[338] <= N440;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[337] <= 1'b0;
    end else if(N421) begin
      mem[337] <= N439;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[336] <= 1'b0;
    end else if(N421) begin
      mem[336] <= N438;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[335] <= 1'b0;
    end else if(N421) begin
      mem[335] <= N437;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[334] <= 1'b0;
    end else if(N421) begin
      mem[334] <= N436;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[333] <= 1'b0;
    end else if(N421) begin
      mem[333] <= N435;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[332] <= 1'b0;
    end else if(N421) begin
      mem[332] <= N434;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[331] <= 1'b0;
    end else if(N421) begin
      mem[331] <= N433;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[330] <= 1'b0;
    end else if(N421) begin
      mem[330] <= N432;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[329] <= 1'b0;
    end else if(N421) begin
      mem[329] <= N431;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[328] <= 1'b0;
    end else if(N421) begin
      mem[328] <= N430;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[327] <= 1'b0;
    end else if(N421) begin
      mem[327] <= N429;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[326] <= 1'b0;
    end else if(N421) begin
      mem[326] <= N428;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[325] <= 1'b0;
    end else if(N421) begin
      mem[325] <= N427;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[324] <= 1'b0;
    end else if(N421) begin
      mem[324] <= N426;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[323] <= 1'b0;
    end else if(N421) begin
      mem[323] <= N425;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[322] <= 1'b0;
    end else if(N421) begin
      mem[322] <= N424;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[321] <= 1'b0;
    end else if(N421) begin
      mem[321] <= N423;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[320] <= 1'b0;
    end else if(N421) begin
      mem[320] <= N422;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[319] <= 1'b0;
    end else if(N355) begin
      mem[319] <= N419;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[318] <= 1'b0;
    end else if(N355) begin
      mem[318] <= N418;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[317] <= 1'b0;
    end else if(N355) begin
      mem[317] <= N417;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[316] <= 1'b0;
    end else if(N355) begin
      mem[316] <= N416;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[315] <= 1'b0;
    end else if(N355) begin
      mem[315] <= N415;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[314] <= 1'b0;
    end else if(N355) begin
      mem[314] <= N414;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[313] <= 1'b0;
    end else if(N355) begin
      mem[313] <= N413;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[312] <= 1'b0;
    end else if(N355) begin
      mem[312] <= N412;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[311] <= 1'b0;
    end else if(N355) begin
      mem[311] <= N411;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[310] <= 1'b0;
    end else if(N355) begin
      mem[310] <= N410;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[309] <= 1'b0;
    end else if(N355) begin
      mem[309] <= N409;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[308] <= 1'b0;
    end else if(N355) begin
      mem[308] <= N408;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[307] <= 1'b0;
    end else if(N355) begin
      mem[307] <= N407;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[306] <= 1'b0;
    end else if(N355) begin
      mem[306] <= N406;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[305] <= 1'b0;
    end else if(N355) begin
      mem[305] <= N405;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[304] <= 1'b0;
    end else if(N355) begin
      mem[304] <= N404;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[303] <= 1'b0;
    end else if(N355) begin
      mem[303] <= N403;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[302] <= 1'b0;
    end else if(N355) begin
      mem[302] <= N402;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[301] <= 1'b0;
    end else if(N355) begin
      mem[301] <= N401;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[300] <= 1'b0;
    end else if(N355) begin
      mem[300] <= N400;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[299] <= 1'b0;
    end else if(N355) begin
      mem[299] <= N399;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[298] <= 1'b0;
    end else if(N355) begin
      mem[298] <= N398;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[297] <= 1'b0;
    end else if(N355) begin
      mem[297] <= N397;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[296] <= 1'b0;
    end else if(N355) begin
      mem[296] <= N396;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[295] <= 1'b0;
    end else if(N355) begin
      mem[295] <= N395;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[294] <= 1'b0;
    end else if(N355) begin
      mem[294] <= N394;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[293] <= 1'b0;
    end else if(N355) begin
      mem[293] <= N393;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[292] <= 1'b0;
    end else if(N355) begin
      mem[292] <= N392;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[291] <= 1'b0;
    end else if(N355) begin
      mem[291] <= N391;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[290] <= 1'b0;
    end else if(N355) begin
      mem[290] <= N390;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[289] <= 1'b0;
    end else if(N355) begin
      mem[289] <= N389;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[288] <= 1'b0;
    end else if(N355) begin
      mem[288] <= N388;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[287] <= 1'b0;
    end else if(N355) begin
      mem[287] <= N387;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[286] <= 1'b0;
    end else if(N355) begin
      mem[286] <= N386;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[285] <= 1'b0;
    end else if(N355) begin
      mem[285] <= N385;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[284] <= 1'b0;
    end else if(N355) begin
      mem[284] <= N384;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[283] <= 1'b0;
    end else if(N355) begin
      mem[283] <= N383;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[282] <= 1'b0;
    end else if(N355) begin
      mem[282] <= N382;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[281] <= 1'b0;
    end else if(N355) begin
      mem[281] <= N381;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[280] <= 1'b0;
    end else if(N355) begin
      mem[280] <= N380;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[279] <= 1'b0;
    end else if(N355) begin
      mem[279] <= N379;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[278] <= 1'b0;
    end else if(N355) begin
      mem[278] <= N378;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[277] <= 1'b0;
    end else if(N355) begin
      mem[277] <= N377;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[276] <= 1'b0;
    end else if(N355) begin
      mem[276] <= N376;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[275] <= 1'b0;
    end else if(N355) begin
      mem[275] <= N375;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[274] <= 1'b0;
    end else if(N355) begin
      mem[274] <= N374;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[273] <= 1'b0;
    end else if(N355) begin
      mem[273] <= N373;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[272] <= 1'b0;
    end else if(N355) begin
      mem[272] <= N372;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[271] <= 1'b0;
    end else if(N355) begin
      mem[271] <= N371;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[270] <= 1'b0;
    end else if(N355) begin
      mem[270] <= N370;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[269] <= 1'b0;
    end else if(N355) begin
      mem[269] <= N369;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[268] <= 1'b0;
    end else if(N355) begin
      mem[268] <= N368;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[267] <= 1'b0;
    end else if(N355) begin
      mem[267] <= N367;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[266] <= 1'b0;
    end else if(N355) begin
      mem[266] <= N366;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[265] <= 1'b0;
    end else if(N355) begin
      mem[265] <= N365;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[264] <= 1'b0;
    end else if(N355) begin
      mem[264] <= N364;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[263] <= 1'b0;
    end else if(N355) begin
      mem[263] <= N363;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[262] <= 1'b0;
    end else if(N355) begin
      mem[262] <= N362;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[261] <= 1'b0;
    end else if(N355) begin
      mem[261] <= N361;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[260] <= 1'b0;
    end else if(N355) begin
      mem[260] <= N360;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[259] <= 1'b0;
    end else if(N355) begin
      mem[259] <= N359;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[258] <= 1'b0;
    end else if(N355) begin
      mem[258] <= N358;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[257] <= 1'b0;
    end else if(N355) begin
      mem[257] <= N357;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[256] <= 1'b0;
    end else if(N355) begin
      mem[256] <= N356;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[255] <= 1'b0;
    end else if(N289) begin
      mem[255] <= N353;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[254] <= 1'b0;
    end else if(N289) begin
      mem[254] <= N352;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[253] <= 1'b0;
    end else if(N289) begin
      mem[253] <= N351;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[252] <= 1'b0;
    end else if(N289) begin
      mem[252] <= N350;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[251] <= 1'b0;
    end else if(N289) begin
      mem[251] <= N349;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[250] <= 1'b0;
    end else if(N289) begin
      mem[250] <= N348;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[249] <= 1'b0;
    end else if(N289) begin
      mem[249] <= N347;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[248] <= 1'b0;
    end else if(N289) begin
      mem[248] <= N346;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[247] <= 1'b0;
    end else if(N289) begin
      mem[247] <= N345;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[246] <= 1'b0;
    end else if(N289) begin
      mem[246] <= N344;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[245] <= 1'b0;
    end else if(N289) begin
      mem[245] <= N343;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[244] <= 1'b0;
    end else if(N289) begin
      mem[244] <= N342;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[243] <= 1'b0;
    end else if(N289) begin
      mem[243] <= N341;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[242] <= 1'b0;
    end else if(N289) begin
      mem[242] <= N340;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[241] <= 1'b0;
    end else if(N289) begin
      mem[241] <= N339;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[240] <= 1'b0;
    end else if(N289) begin
      mem[240] <= N338;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[239] <= 1'b0;
    end else if(N289) begin
      mem[239] <= N337;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[238] <= 1'b0;
    end else if(N289) begin
      mem[238] <= N336;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[237] <= 1'b0;
    end else if(N289) begin
      mem[237] <= N335;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[236] <= 1'b0;
    end else if(N289) begin
      mem[236] <= N334;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[235] <= 1'b0;
    end else if(N289) begin
      mem[235] <= N333;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[234] <= 1'b0;
    end else if(N289) begin
      mem[234] <= N332;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[233] <= 1'b0;
    end else if(N289) begin
      mem[233] <= N331;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[232] <= 1'b0;
    end else if(N289) begin
      mem[232] <= N330;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[231] <= 1'b0;
    end else if(N289) begin
      mem[231] <= N329;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[230] <= 1'b0;
    end else if(N289) begin
      mem[230] <= N328;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[229] <= 1'b0;
    end else if(N289) begin
      mem[229] <= N327;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[228] <= 1'b0;
    end else if(N289) begin
      mem[228] <= N326;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[227] <= 1'b0;
    end else if(N289) begin
      mem[227] <= N325;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[226] <= 1'b0;
    end else if(N289) begin
      mem[226] <= N324;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[225] <= 1'b0;
    end else if(N289) begin
      mem[225] <= N323;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[224] <= 1'b0;
    end else if(N289) begin
      mem[224] <= N322;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[223] <= 1'b0;
    end else if(N289) begin
      mem[223] <= N321;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[222] <= 1'b0;
    end else if(N289) begin
      mem[222] <= N320;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[221] <= 1'b0;
    end else if(N289) begin
      mem[221] <= N319;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[220] <= 1'b0;
    end else if(N289) begin
      mem[220] <= N318;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[219] <= 1'b0;
    end else if(N289) begin
      mem[219] <= N317;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[218] <= 1'b0;
    end else if(N289) begin
      mem[218] <= N316;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[217] <= 1'b0;
    end else if(N289) begin
      mem[217] <= N315;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[216] <= 1'b0;
    end else if(N289) begin
      mem[216] <= N314;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[215] <= 1'b0;
    end else if(N289) begin
      mem[215] <= N313;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[214] <= 1'b0;
    end else if(N289) begin
      mem[214] <= N312;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[213] <= 1'b0;
    end else if(N289) begin
      mem[213] <= N311;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[212] <= 1'b0;
    end else if(N289) begin
      mem[212] <= N310;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[211] <= 1'b0;
    end else if(N289) begin
      mem[211] <= N309;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[210] <= 1'b0;
    end else if(N289) begin
      mem[210] <= N308;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[209] <= 1'b0;
    end else if(N289) begin
      mem[209] <= N307;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[208] <= 1'b0;
    end else if(N289) begin
      mem[208] <= N306;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[207] <= 1'b0;
    end else if(N289) begin
      mem[207] <= N305;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[206] <= 1'b0;
    end else if(N289) begin
      mem[206] <= N304;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[205] <= 1'b0;
    end else if(N289) begin
      mem[205] <= N303;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[204] <= 1'b0;
    end else if(N289) begin
      mem[204] <= N302;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[203] <= 1'b0;
    end else if(N289) begin
      mem[203] <= N301;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[202] <= 1'b0;
    end else if(N289) begin
      mem[202] <= N300;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[201] <= 1'b0;
    end else if(N289) begin
      mem[201] <= N299;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[200] <= 1'b0;
    end else if(N289) begin
      mem[200] <= N298;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[199] <= 1'b0;
    end else if(N289) begin
      mem[199] <= N297;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[198] <= 1'b0;
    end else if(N289) begin
      mem[198] <= N296;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[197] <= 1'b0;
    end else if(N289) begin
      mem[197] <= N295;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[196] <= 1'b0;
    end else if(N289) begin
      mem[196] <= N294;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[195] <= 1'b0;
    end else if(N289) begin
      mem[195] <= N293;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[194] <= 1'b0;
    end else if(N289) begin
      mem[194] <= N292;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[193] <= 1'b0;
    end else if(N289) begin
      mem[193] <= N291;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[192] <= 1'b0;
    end else if(N289) begin
      mem[192] <= N290;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[191] <= 1'b0;
    end else if(N223) begin
      mem[191] <= N287;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[190] <= 1'b0;
    end else if(N223) begin
      mem[190] <= N286;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[189] <= 1'b0;
    end else if(N223) begin
      mem[189] <= N285;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[188] <= 1'b0;
    end else if(N223) begin
      mem[188] <= N284;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[187] <= 1'b0;
    end else if(N223) begin
      mem[187] <= N283;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[186] <= 1'b0;
    end else if(N223) begin
      mem[186] <= N282;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[185] <= 1'b0;
    end else if(N223) begin
      mem[185] <= N281;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[184] <= 1'b0;
    end else if(N223) begin
      mem[184] <= N280;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[183] <= 1'b0;
    end else if(N223) begin
      mem[183] <= N279;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[182] <= 1'b0;
    end else if(N223) begin
      mem[182] <= N278;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[181] <= 1'b0;
    end else if(N223) begin
      mem[181] <= N277;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[180] <= 1'b0;
    end else if(N223) begin
      mem[180] <= N276;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[179] <= 1'b0;
    end else if(N223) begin
      mem[179] <= N275;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[178] <= 1'b0;
    end else if(N223) begin
      mem[178] <= N274;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[177] <= 1'b0;
    end else if(N223) begin
      mem[177] <= N273;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[176] <= 1'b0;
    end else if(N223) begin
      mem[176] <= N272;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[175] <= 1'b0;
    end else if(N223) begin
      mem[175] <= N271;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[174] <= 1'b0;
    end else if(N223) begin
      mem[174] <= N270;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[173] <= 1'b0;
    end else if(N223) begin
      mem[173] <= N269;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[172] <= 1'b0;
    end else if(N223) begin
      mem[172] <= N268;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[171] <= 1'b0;
    end else if(N223) begin
      mem[171] <= N267;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[170] <= 1'b0;
    end else if(N223) begin
      mem[170] <= N266;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[169] <= 1'b0;
    end else if(N223) begin
      mem[169] <= N265;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[168] <= 1'b0;
    end else if(N223) begin
      mem[168] <= N264;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[167] <= 1'b0;
    end else if(N223) begin
      mem[167] <= N263;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[166] <= 1'b0;
    end else if(N223) begin
      mem[166] <= N262;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[165] <= 1'b0;
    end else if(N223) begin
      mem[165] <= N261;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[164] <= 1'b0;
    end else if(N223) begin
      mem[164] <= N260;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[163] <= 1'b0;
    end else if(N223) begin
      mem[163] <= N259;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[162] <= 1'b0;
    end else if(N223) begin
      mem[162] <= N258;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[161] <= 1'b0;
    end else if(N223) begin
      mem[161] <= N257;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[160] <= 1'b0;
    end else if(N223) begin
      mem[160] <= N256;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[159] <= 1'b0;
    end else if(N223) begin
      mem[159] <= N255;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[158] <= 1'b0;
    end else if(N223) begin
      mem[158] <= N254;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[157] <= 1'b0;
    end else if(N223) begin
      mem[157] <= N253;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[156] <= 1'b0;
    end else if(N223) begin
      mem[156] <= N252;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[155] <= 1'b0;
    end else if(N223) begin
      mem[155] <= N251;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[154] <= 1'b0;
    end else if(N223) begin
      mem[154] <= N250;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[153] <= 1'b0;
    end else if(N223) begin
      mem[153] <= N249;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[152] <= 1'b0;
    end else if(N223) begin
      mem[152] <= N248;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[151] <= 1'b0;
    end else if(N223) begin
      mem[151] <= N247;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[150] <= 1'b0;
    end else if(N223) begin
      mem[150] <= N246;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[149] <= 1'b0;
    end else if(N223) begin
      mem[149] <= N245;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[148] <= 1'b0;
    end else if(N223) begin
      mem[148] <= N244;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[147] <= 1'b0;
    end else if(N223) begin
      mem[147] <= N243;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[146] <= 1'b0;
    end else if(N223) begin
      mem[146] <= N242;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[145] <= 1'b0;
    end else if(N223) begin
      mem[145] <= N241;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[144] <= 1'b0;
    end else if(N223) begin
      mem[144] <= N240;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[143] <= 1'b0;
    end else if(N223) begin
      mem[143] <= N239;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[142] <= 1'b0;
    end else if(N223) begin
      mem[142] <= N238;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[141] <= 1'b0;
    end else if(N223) begin
      mem[141] <= N237;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[140] <= 1'b0;
    end else if(N223) begin
      mem[140] <= N236;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[139] <= 1'b0;
    end else if(N223) begin
      mem[139] <= N235;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[138] <= 1'b0;
    end else if(N223) begin
      mem[138] <= N234;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[137] <= 1'b0;
    end else if(N223) begin
      mem[137] <= N233;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[136] <= 1'b0;
    end else if(N223) begin
      mem[136] <= N232;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[135] <= 1'b0;
    end else if(N223) begin
      mem[135] <= N231;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[134] <= 1'b0;
    end else if(N223) begin
      mem[134] <= N230;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[133] <= 1'b0;
    end else if(N223) begin
      mem[133] <= N229;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[132] <= 1'b0;
    end else if(N223) begin
      mem[132] <= N228;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[131] <= 1'b0;
    end else if(N223) begin
      mem[131] <= N227;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[130] <= 1'b0;
    end else if(N223) begin
      mem[130] <= N226;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[129] <= 1'b0;
    end else if(N223) begin
      mem[129] <= N225;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[128] <= 1'b0;
    end else if(N223) begin
      mem[128] <= N224;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[127] <= 1'b0;
    end else if(N157) begin
      mem[127] <= N221;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[126] <= 1'b0;
    end else if(N157) begin
      mem[126] <= N220;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[125] <= 1'b0;
    end else if(N157) begin
      mem[125] <= N219;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[124] <= 1'b0;
    end else if(N157) begin
      mem[124] <= N218;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[123] <= 1'b0;
    end else if(N157) begin
      mem[123] <= N217;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[122] <= 1'b0;
    end else if(N157) begin
      mem[122] <= N216;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[121] <= 1'b0;
    end else if(N157) begin
      mem[121] <= N215;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[120] <= 1'b0;
    end else if(N157) begin
      mem[120] <= N214;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[119] <= 1'b0;
    end else if(N157) begin
      mem[119] <= N213;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[118] <= 1'b0;
    end else if(N157) begin
      mem[118] <= N212;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[117] <= 1'b0;
    end else if(N157) begin
      mem[117] <= N211;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[116] <= 1'b0;
    end else if(N157) begin
      mem[116] <= N210;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[115] <= 1'b0;
    end else if(N157) begin
      mem[115] <= N209;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[114] <= 1'b0;
    end else if(N157) begin
      mem[114] <= N208;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[113] <= 1'b0;
    end else if(N157) begin
      mem[113] <= N207;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[112] <= 1'b0;
    end else if(N157) begin
      mem[112] <= N206;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[111] <= 1'b0;
    end else if(N157) begin
      mem[111] <= N205;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[110] <= 1'b0;
    end else if(N157) begin
      mem[110] <= N204;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[109] <= 1'b0;
    end else if(N157) begin
      mem[109] <= N203;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[108] <= 1'b0;
    end else if(N157) begin
      mem[108] <= N202;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[107] <= 1'b0;
    end else if(N157) begin
      mem[107] <= N201;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[106] <= 1'b0;
    end else if(N157) begin
      mem[106] <= N200;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[105] <= 1'b0;
    end else if(N157) begin
      mem[105] <= N199;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[104] <= 1'b0;
    end else if(N157) begin
      mem[104] <= N198;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[103] <= 1'b0;
    end else if(N157) begin
      mem[103] <= N197;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[102] <= 1'b0;
    end else if(N157) begin
      mem[102] <= N196;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[101] <= 1'b0;
    end else if(N157) begin
      mem[101] <= N195;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[100] <= 1'b0;
    end else if(N157) begin
      mem[100] <= N194;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[99] <= 1'b0;
    end else if(N157) begin
      mem[99] <= N193;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[98] <= 1'b0;
    end else if(N157) begin
      mem[98] <= N192;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[97] <= 1'b0;
    end else if(N157) begin
      mem[97] <= N191;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[96] <= 1'b0;
    end else if(N157) begin
      mem[96] <= N190;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[95] <= 1'b0;
    end else if(N157) begin
      mem[95] <= N189;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[94] <= 1'b0;
    end else if(N157) begin
      mem[94] <= N188;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[93] <= 1'b0;
    end else if(N157) begin
      mem[93] <= N187;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[92] <= 1'b0;
    end else if(N157) begin
      mem[92] <= N186;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[91] <= 1'b0;
    end else if(N157) begin
      mem[91] <= N185;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[90] <= 1'b0;
    end else if(N157) begin
      mem[90] <= N184;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[89] <= 1'b0;
    end else if(N157) begin
      mem[89] <= N183;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[88] <= 1'b0;
    end else if(N157) begin
      mem[88] <= N182;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[87] <= 1'b0;
    end else if(N157) begin
      mem[87] <= N181;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[86] <= 1'b0;
    end else if(N157) begin
      mem[86] <= N180;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[85] <= 1'b0;
    end else if(N157) begin
      mem[85] <= N179;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[84] <= 1'b0;
    end else if(N157) begin
      mem[84] <= N178;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[83] <= 1'b0;
    end else if(N157) begin
      mem[83] <= N177;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[82] <= 1'b0;
    end else if(N157) begin
      mem[82] <= N176;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[81] <= 1'b0;
    end else if(N157) begin
      mem[81] <= N175;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[80] <= 1'b0;
    end else if(N157) begin
      mem[80] <= N174;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[79] <= 1'b0;
    end else if(N157) begin
      mem[79] <= N173;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[78] <= 1'b0;
    end else if(N157) begin
      mem[78] <= N172;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[77] <= 1'b0;
    end else if(N157) begin
      mem[77] <= N171;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[76] <= 1'b0;
    end else if(N157) begin
      mem[76] <= N170;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[75] <= 1'b0;
    end else if(N157) begin
      mem[75] <= N169;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[74] <= 1'b0;
    end else if(N157) begin
      mem[74] <= N168;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[73] <= 1'b0;
    end else if(N157) begin
      mem[73] <= N167;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[72] <= 1'b0;
    end else if(N157) begin
      mem[72] <= N166;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[71] <= 1'b0;
    end else if(N157) begin
      mem[71] <= N165;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[70] <= 1'b0;
    end else if(N157) begin
      mem[70] <= N164;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[69] <= 1'b0;
    end else if(N157) begin
      mem[69] <= N163;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[68] <= 1'b0;
    end else if(N157) begin
      mem[68] <= N162;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[67] <= 1'b0;
    end else if(N157) begin
      mem[67] <= N161;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[66] <= 1'b0;
    end else if(N157) begin
      mem[66] <= N160;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[65] <= 1'b0;
    end else if(N157) begin
      mem[65] <= N159;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[64] <= 1'b0;
    end else if(N157) begin
      mem[64] <= N158;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[63] <= 1'b0;
    end else if(1'b1) begin
      mem[63] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[62] <= 1'b0;
    end else if(1'b1) begin
      mem[62] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[61] <= 1'b0;
    end else if(1'b1) begin
      mem[61] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[60] <= 1'b0;
    end else if(1'b1) begin
      mem[60] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[59] <= 1'b0;
    end else if(1'b1) begin
      mem[59] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[58] <= 1'b0;
    end else if(1'b1) begin
      mem[58] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[57] <= 1'b0;
    end else if(1'b1) begin
      mem[57] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[56] <= 1'b0;
    end else if(1'b1) begin
      mem[56] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[55] <= 1'b0;
    end else if(1'b1) begin
      mem[55] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[54] <= 1'b0;
    end else if(1'b1) begin
      mem[54] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[53] <= 1'b0;
    end else if(1'b1) begin
      mem[53] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[52] <= 1'b0;
    end else if(1'b1) begin
      mem[52] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[51] <= 1'b0;
    end else if(1'b1) begin
      mem[51] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[50] <= 1'b0;
    end else if(1'b1) begin
      mem[50] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[49] <= 1'b0;
    end else if(1'b1) begin
      mem[49] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[48] <= 1'b0;
    end else if(1'b1) begin
      mem[48] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[47] <= 1'b0;
    end else if(1'b1) begin
      mem[47] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[46] <= 1'b0;
    end else if(1'b1) begin
      mem[46] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[45] <= 1'b0;
    end else if(1'b1) begin
      mem[45] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[44] <= 1'b0;
    end else if(1'b1) begin
      mem[44] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[43] <= 1'b0;
    end else if(1'b1) begin
      mem[43] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[42] <= 1'b0;
    end else if(1'b1) begin
      mem[42] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[41] <= 1'b0;
    end else if(1'b1) begin
      mem[41] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[40] <= 1'b0;
    end else if(1'b1) begin
      mem[40] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[39] <= 1'b0;
    end else if(1'b1) begin
      mem[39] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[38] <= 1'b0;
    end else if(1'b1) begin
      mem[38] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[37] <= 1'b0;
    end else if(1'b1) begin
      mem[37] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[36] <= 1'b0;
    end else if(1'b1) begin
      mem[36] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[35] <= 1'b0;
    end else if(1'b1) begin
      mem[35] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[34] <= 1'b0;
    end else if(1'b1) begin
      mem[34] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[33] <= 1'b0;
    end else if(1'b1) begin
      mem[33] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[32] <= 1'b0;
    end else if(1'b1) begin
      mem[32] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[31] <= 1'b0;
    end else if(1'b1) begin
      mem[31] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[30] <= 1'b0;
    end else if(1'b1) begin
      mem[30] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[29] <= 1'b0;
    end else if(1'b1) begin
      mem[29] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[28] <= 1'b0;
    end else if(1'b1) begin
      mem[28] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[27] <= 1'b0;
    end else if(1'b1) begin
      mem[27] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[26] <= 1'b0;
    end else if(1'b1) begin
      mem[26] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[25] <= 1'b0;
    end else if(1'b1) begin
      mem[25] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[24] <= 1'b0;
    end else if(1'b1) begin
      mem[24] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[23] <= 1'b0;
    end else if(1'b1) begin
      mem[23] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[22] <= 1'b0;
    end else if(1'b1) begin
      mem[22] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[21] <= 1'b0;
    end else if(1'b1) begin
      mem[21] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[20] <= 1'b0;
    end else if(1'b1) begin
      mem[20] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[19] <= 1'b0;
    end else if(1'b1) begin
      mem[19] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[18] <= 1'b0;
    end else if(1'b1) begin
      mem[18] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[17] <= 1'b0;
    end else if(1'b1) begin
      mem[17] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[16] <= 1'b0;
    end else if(1'b1) begin
      mem[16] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[15] <= 1'b0;
    end else if(1'b1) begin
      mem[15] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[14] <= 1'b0;
    end else if(1'b1) begin
      mem[14] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[13] <= 1'b0;
    end else if(1'b1) begin
      mem[13] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[12] <= 1'b0;
    end else if(1'b1) begin
      mem[12] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[11] <= 1'b0;
    end else if(1'b1) begin
      mem[11] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[10] <= 1'b0;
    end else if(1'b1) begin
      mem[10] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[9] <= 1'b0;
    end else if(1'b1) begin
      mem[9] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[8] <= 1'b0;
    end else if(1'b1) begin
      mem[8] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[7] <= 1'b0;
    end else if(1'b1) begin
      mem[7] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[6] <= 1'b0;
    end else if(1'b1) begin
      mem[6] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[5] <= 1'b0;
    end else if(1'b1) begin
      mem[5] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[4] <= 1'b0;
    end else if(1'b1) begin
      mem[4] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[3] <= 1'b0;
    end else if(1'b1) begin
      mem[3] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[2] <= 1'b0;
    end else if(1'b1) begin
      mem[2] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[1] <= 1'b0;
    end else if(1'b1) begin
      mem[1] <= 1'b0;
    end 
  end


  always @(posedge clk_i or posedge N155) begin
    if(N155) begin
      mem[0] <= 1'b0;
    end else if(1'b1) begin
      mem[0] <= 1'b0;
    end 
  end

  assign rdata_o[63] = (N2235)? mem[63] : 
                       (N2237)? mem[127] : 
                       (N2239)? mem[191] : 
                       (N2241)? mem[255] : 
                       (N2243)? mem[319] : 
                       (N2245)? mem[383] : 
                       (N2247)? mem[447] : 
                       (N2249)? mem[511] : 
                       (N2251)? mem[575] : 
                       (N2253)? mem[639] : 
                       (N2255)? mem[703] : 
                       (N2257)? mem[767] : 
                       (N2259)? mem[831] : 
                       (N2261)? mem[895] : 
                       (N2263)? mem[959] : 
                       (N2265)? mem[1023] : 
                       (N2236)? mem[1087] : 
                       (N2238)? mem[1151] : 
                       (N2240)? mem[1215] : 
                       (N2242)? mem[1279] : 
                       (N2244)? mem[1343] : 
                       (N2246)? mem[1407] : 
                       (N2248)? mem[1471] : 
                       (N2250)? mem[1535] : 
                       (N2252)? mem[1599] : 
                       (N2254)? mem[1663] : 
                       (N2256)? mem[1727] : 
                       (N2258)? mem[1791] : 
                       (N2260)? mem[1855] : 
                       (N2262)? mem[1919] : 
                       (N2264)? mem[1983] : 
                       (N2266)? mem[2047] : 1'b0;
  assign rdata_o[62] = (N2235)? mem[62] : 
                       (N2237)? mem[126] : 
                       (N2239)? mem[190] : 
                       (N2241)? mem[254] : 
                       (N2243)? mem[318] : 
                       (N2245)? mem[382] : 
                       (N2247)? mem[446] : 
                       (N2249)? mem[510] : 
                       (N2251)? mem[574] : 
                       (N2253)? mem[638] : 
                       (N2255)? mem[702] : 
                       (N2257)? mem[766] : 
                       (N2259)? mem[830] : 
                       (N2261)? mem[894] : 
                       (N2263)? mem[958] : 
                       (N2265)? mem[1022] : 
                       (N2236)? mem[1086] : 
                       (N2238)? mem[1150] : 
                       (N2240)? mem[1214] : 
                       (N2242)? mem[1278] : 
                       (N2244)? mem[1342] : 
                       (N2246)? mem[1406] : 
                       (N2248)? mem[1470] : 
                       (N2250)? mem[1534] : 
                       (N2252)? mem[1598] : 
                       (N2254)? mem[1662] : 
                       (N2256)? mem[1726] : 
                       (N2258)? mem[1790] : 
                       (N2260)? mem[1854] : 
                       (N2262)? mem[1918] : 
                       (N2264)? mem[1982] : 
                       (N2266)? mem[2046] : 1'b0;
  assign rdata_o[61] = (N2235)? mem[61] : 
                       (N2237)? mem[125] : 
                       (N2239)? mem[189] : 
                       (N2241)? mem[253] : 
                       (N2243)? mem[317] : 
                       (N2245)? mem[381] : 
                       (N2247)? mem[445] : 
                       (N2249)? mem[509] : 
                       (N2251)? mem[573] : 
                       (N2253)? mem[637] : 
                       (N2255)? mem[701] : 
                       (N2257)? mem[765] : 
                       (N2259)? mem[829] : 
                       (N2261)? mem[893] : 
                       (N2263)? mem[957] : 
                       (N2265)? mem[1021] : 
                       (N2236)? mem[1085] : 
                       (N2238)? mem[1149] : 
                       (N2240)? mem[1213] : 
                       (N2242)? mem[1277] : 
                       (N2244)? mem[1341] : 
                       (N2246)? mem[1405] : 
                       (N2248)? mem[1469] : 
                       (N2250)? mem[1533] : 
                       (N2252)? mem[1597] : 
                       (N2254)? mem[1661] : 
                       (N2256)? mem[1725] : 
                       (N2258)? mem[1789] : 
                       (N2260)? mem[1853] : 
                       (N2262)? mem[1917] : 
                       (N2264)? mem[1981] : 
                       (N2266)? mem[2045] : 1'b0;
  assign rdata_o[60] = (N2235)? mem[60] : 
                       (N2237)? mem[124] : 
                       (N2239)? mem[188] : 
                       (N2241)? mem[252] : 
                       (N2243)? mem[316] : 
                       (N2245)? mem[380] : 
                       (N2247)? mem[444] : 
                       (N2249)? mem[508] : 
                       (N2251)? mem[572] : 
                       (N2253)? mem[636] : 
                       (N2255)? mem[700] : 
                       (N2257)? mem[764] : 
                       (N2259)? mem[828] : 
                       (N2261)? mem[892] : 
                       (N2263)? mem[956] : 
                       (N2265)? mem[1020] : 
                       (N2236)? mem[1084] : 
                       (N2238)? mem[1148] : 
                       (N2240)? mem[1212] : 
                       (N2242)? mem[1276] : 
                       (N2244)? mem[1340] : 
                       (N2246)? mem[1404] : 
                       (N2248)? mem[1468] : 
                       (N2250)? mem[1532] : 
                       (N2252)? mem[1596] : 
                       (N2254)? mem[1660] : 
                       (N2256)? mem[1724] : 
                       (N2258)? mem[1788] : 
                       (N2260)? mem[1852] : 
                       (N2262)? mem[1916] : 
                       (N2264)? mem[1980] : 
                       (N2266)? mem[2044] : 1'b0;
  assign rdata_o[59] = (N2235)? mem[59] : 
                       (N2237)? mem[123] : 
                       (N2239)? mem[187] : 
                       (N2241)? mem[251] : 
                       (N2243)? mem[315] : 
                       (N2245)? mem[379] : 
                       (N2247)? mem[443] : 
                       (N2249)? mem[507] : 
                       (N2251)? mem[571] : 
                       (N2253)? mem[635] : 
                       (N2255)? mem[699] : 
                       (N2257)? mem[763] : 
                       (N2259)? mem[827] : 
                       (N2261)? mem[891] : 
                       (N2263)? mem[955] : 
                       (N2265)? mem[1019] : 
                       (N2236)? mem[1083] : 
                       (N2238)? mem[1147] : 
                       (N2240)? mem[1211] : 
                       (N2242)? mem[1275] : 
                       (N2244)? mem[1339] : 
                       (N2246)? mem[1403] : 
                       (N2248)? mem[1467] : 
                       (N2250)? mem[1531] : 
                       (N2252)? mem[1595] : 
                       (N2254)? mem[1659] : 
                       (N2256)? mem[1723] : 
                       (N2258)? mem[1787] : 
                       (N2260)? mem[1851] : 
                       (N2262)? mem[1915] : 
                       (N2264)? mem[1979] : 
                       (N2266)? mem[2043] : 1'b0;
  assign rdata_o[58] = (N2235)? mem[58] : 
                       (N2237)? mem[122] : 
                       (N2239)? mem[186] : 
                       (N2241)? mem[250] : 
                       (N2243)? mem[314] : 
                       (N2245)? mem[378] : 
                       (N2247)? mem[442] : 
                       (N2249)? mem[506] : 
                       (N2251)? mem[570] : 
                       (N2253)? mem[634] : 
                       (N2255)? mem[698] : 
                       (N2257)? mem[762] : 
                       (N2259)? mem[826] : 
                       (N2261)? mem[890] : 
                       (N2263)? mem[954] : 
                       (N2265)? mem[1018] : 
                       (N2236)? mem[1082] : 
                       (N2238)? mem[1146] : 
                       (N2240)? mem[1210] : 
                       (N2242)? mem[1274] : 
                       (N2244)? mem[1338] : 
                       (N2246)? mem[1402] : 
                       (N2248)? mem[1466] : 
                       (N2250)? mem[1530] : 
                       (N2252)? mem[1594] : 
                       (N2254)? mem[1658] : 
                       (N2256)? mem[1722] : 
                       (N2258)? mem[1786] : 
                       (N2260)? mem[1850] : 
                       (N2262)? mem[1914] : 
                       (N2264)? mem[1978] : 
                       (N2266)? mem[2042] : 1'b0;
  assign rdata_o[57] = (N2235)? mem[57] : 
                       (N2237)? mem[121] : 
                       (N2239)? mem[185] : 
                       (N2241)? mem[249] : 
                       (N2243)? mem[313] : 
                       (N2245)? mem[377] : 
                       (N2247)? mem[441] : 
                       (N2249)? mem[505] : 
                       (N2251)? mem[569] : 
                       (N2253)? mem[633] : 
                       (N2255)? mem[697] : 
                       (N2257)? mem[761] : 
                       (N2259)? mem[825] : 
                       (N2261)? mem[889] : 
                       (N2263)? mem[953] : 
                       (N2265)? mem[1017] : 
                       (N2236)? mem[1081] : 
                       (N2238)? mem[1145] : 
                       (N2240)? mem[1209] : 
                       (N2242)? mem[1273] : 
                       (N2244)? mem[1337] : 
                       (N2246)? mem[1401] : 
                       (N2248)? mem[1465] : 
                       (N2250)? mem[1529] : 
                       (N2252)? mem[1593] : 
                       (N2254)? mem[1657] : 
                       (N2256)? mem[1721] : 
                       (N2258)? mem[1785] : 
                       (N2260)? mem[1849] : 
                       (N2262)? mem[1913] : 
                       (N2264)? mem[1977] : 
                       (N2266)? mem[2041] : 1'b0;
  assign rdata_o[56] = (N2235)? mem[56] : 
                       (N2237)? mem[120] : 
                       (N2239)? mem[184] : 
                       (N2241)? mem[248] : 
                       (N2243)? mem[312] : 
                       (N2245)? mem[376] : 
                       (N2247)? mem[440] : 
                       (N2249)? mem[504] : 
                       (N2251)? mem[568] : 
                       (N2253)? mem[632] : 
                       (N2255)? mem[696] : 
                       (N2257)? mem[760] : 
                       (N2259)? mem[824] : 
                       (N2261)? mem[888] : 
                       (N2263)? mem[952] : 
                       (N2265)? mem[1016] : 
                       (N2236)? mem[1080] : 
                       (N2238)? mem[1144] : 
                       (N2240)? mem[1208] : 
                       (N2242)? mem[1272] : 
                       (N2244)? mem[1336] : 
                       (N2246)? mem[1400] : 
                       (N2248)? mem[1464] : 
                       (N2250)? mem[1528] : 
                       (N2252)? mem[1592] : 
                       (N2254)? mem[1656] : 
                       (N2256)? mem[1720] : 
                       (N2258)? mem[1784] : 
                       (N2260)? mem[1848] : 
                       (N2262)? mem[1912] : 
                       (N2264)? mem[1976] : 
                       (N2266)? mem[2040] : 1'b0;
  assign rdata_o[55] = (N2235)? mem[55] : 
                       (N2237)? mem[119] : 
                       (N2239)? mem[183] : 
                       (N2241)? mem[247] : 
                       (N2243)? mem[311] : 
                       (N2245)? mem[375] : 
                       (N2247)? mem[439] : 
                       (N2249)? mem[503] : 
                       (N2251)? mem[567] : 
                       (N2253)? mem[631] : 
                       (N2255)? mem[695] : 
                       (N2257)? mem[759] : 
                       (N2259)? mem[823] : 
                       (N2261)? mem[887] : 
                       (N2263)? mem[951] : 
                       (N2265)? mem[1015] : 
                       (N2236)? mem[1079] : 
                       (N2238)? mem[1143] : 
                       (N2240)? mem[1207] : 
                       (N2242)? mem[1271] : 
                       (N2244)? mem[1335] : 
                       (N2246)? mem[1399] : 
                       (N2248)? mem[1463] : 
                       (N2250)? mem[1527] : 
                       (N2252)? mem[1591] : 
                       (N2254)? mem[1655] : 
                       (N2256)? mem[1719] : 
                       (N2258)? mem[1783] : 
                       (N2260)? mem[1847] : 
                       (N2262)? mem[1911] : 
                       (N2264)? mem[1975] : 
                       (N2266)? mem[2039] : 1'b0;
  assign rdata_o[54] = (N2235)? mem[54] : 
                       (N2237)? mem[118] : 
                       (N2239)? mem[182] : 
                       (N2241)? mem[246] : 
                       (N2243)? mem[310] : 
                       (N2245)? mem[374] : 
                       (N2247)? mem[438] : 
                       (N2249)? mem[502] : 
                       (N2251)? mem[566] : 
                       (N2253)? mem[630] : 
                       (N2255)? mem[694] : 
                       (N2257)? mem[758] : 
                       (N2259)? mem[822] : 
                       (N2261)? mem[886] : 
                       (N2263)? mem[950] : 
                       (N2265)? mem[1014] : 
                       (N2236)? mem[1078] : 
                       (N2238)? mem[1142] : 
                       (N2240)? mem[1206] : 
                       (N2242)? mem[1270] : 
                       (N2244)? mem[1334] : 
                       (N2246)? mem[1398] : 
                       (N2248)? mem[1462] : 
                       (N2250)? mem[1526] : 
                       (N2252)? mem[1590] : 
                       (N2254)? mem[1654] : 
                       (N2256)? mem[1718] : 
                       (N2258)? mem[1782] : 
                       (N2260)? mem[1846] : 
                       (N2262)? mem[1910] : 
                       (N2264)? mem[1974] : 
                       (N2266)? mem[2038] : 1'b0;
  assign rdata_o[53] = (N2235)? mem[53] : 
                       (N2237)? mem[117] : 
                       (N2239)? mem[181] : 
                       (N2241)? mem[245] : 
                       (N2243)? mem[309] : 
                       (N2245)? mem[373] : 
                       (N2247)? mem[437] : 
                       (N2249)? mem[501] : 
                       (N2251)? mem[565] : 
                       (N2253)? mem[629] : 
                       (N2255)? mem[693] : 
                       (N2257)? mem[757] : 
                       (N2259)? mem[821] : 
                       (N2261)? mem[885] : 
                       (N2263)? mem[949] : 
                       (N2265)? mem[1013] : 
                       (N2236)? mem[1077] : 
                       (N2238)? mem[1141] : 
                       (N2240)? mem[1205] : 
                       (N2242)? mem[1269] : 
                       (N2244)? mem[1333] : 
                       (N2246)? mem[1397] : 
                       (N2248)? mem[1461] : 
                       (N2250)? mem[1525] : 
                       (N2252)? mem[1589] : 
                       (N2254)? mem[1653] : 
                       (N2256)? mem[1717] : 
                       (N2258)? mem[1781] : 
                       (N2260)? mem[1845] : 
                       (N2262)? mem[1909] : 
                       (N2264)? mem[1973] : 
                       (N2266)? mem[2037] : 1'b0;
  assign rdata_o[52] = (N2235)? mem[52] : 
                       (N2237)? mem[116] : 
                       (N2239)? mem[180] : 
                       (N2241)? mem[244] : 
                       (N2243)? mem[308] : 
                       (N2245)? mem[372] : 
                       (N2247)? mem[436] : 
                       (N2249)? mem[500] : 
                       (N2251)? mem[564] : 
                       (N2253)? mem[628] : 
                       (N2255)? mem[692] : 
                       (N2257)? mem[756] : 
                       (N2259)? mem[820] : 
                       (N2261)? mem[884] : 
                       (N2263)? mem[948] : 
                       (N2265)? mem[1012] : 
                       (N2236)? mem[1076] : 
                       (N2238)? mem[1140] : 
                       (N2240)? mem[1204] : 
                       (N2242)? mem[1268] : 
                       (N2244)? mem[1332] : 
                       (N2246)? mem[1396] : 
                       (N2248)? mem[1460] : 
                       (N2250)? mem[1524] : 
                       (N2252)? mem[1588] : 
                       (N2254)? mem[1652] : 
                       (N2256)? mem[1716] : 
                       (N2258)? mem[1780] : 
                       (N2260)? mem[1844] : 
                       (N2262)? mem[1908] : 
                       (N2264)? mem[1972] : 
                       (N2266)? mem[2036] : 1'b0;
  assign rdata_o[51] = (N2235)? mem[51] : 
                       (N2237)? mem[115] : 
                       (N2239)? mem[179] : 
                       (N2241)? mem[243] : 
                       (N2243)? mem[307] : 
                       (N2245)? mem[371] : 
                       (N2247)? mem[435] : 
                       (N2249)? mem[499] : 
                       (N2251)? mem[563] : 
                       (N2253)? mem[627] : 
                       (N2255)? mem[691] : 
                       (N2257)? mem[755] : 
                       (N2259)? mem[819] : 
                       (N2261)? mem[883] : 
                       (N2263)? mem[947] : 
                       (N2265)? mem[1011] : 
                       (N2236)? mem[1075] : 
                       (N2238)? mem[1139] : 
                       (N2240)? mem[1203] : 
                       (N2242)? mem[1267] : 
                       (N2244)? mem[1331] : 
                       (N2246)? mem[1395] : 
                       (N2248)? mem[1459] : 
                       (N2250)? mem[1523] : 
                       (N2252)? mem[1587] : 
                       (N2254)? mem[1651] : 
                       (N2256)? mem[1715] : 
                       (N2258)? mem[1779] : 
                       (N2260)? mem[1843] : 
                       (N2262)? mem[1907] : 
                       (N2264)? mem[1971] : 
                       (N2266)? mem[2035] : 1'b0;
  assign rdata_o[50] = (N2235)? mem[50] : 
                       (N2237)? mem[114] : 
                       (N2239)? mem[178] : 
                       (N2241)? mem[242] : 
                       (N2243)? mem[306] : 
                       (N2245)? mem[370] : 
                       (N2247)? mem[434] : 
                       (N2249)? mem[498] : 
                       (N2251)? mem[562] : 
                       (N2253)? mem[626] : 
                       (N2255)? mem[690] : 
                       (N2257)? mem[754] : 
                       (N2259)? mem[818] : 
                       (N2261)? mem[882] : 
                       (N2263)? mem[946] : 
                       (N2265)? mem[1010] : 
                       (N2236)? mem[1074] : 
                       (N2238)? mem[1138] : 
                       (N2240)? mem[1202] : 
                       (N2242)? mem[1266] : 
                       (N2244)? mem[1330] : 
                       (N2246)? mem[1394] : 
                       (N2248)? mem[1458] : 
                       (N2250)? mem[1522] : 
                       (N2252)? mem[1586] : 
                       (N2254)? mem[1650] : 
                       (N2256)? mem[1714] : 
                       (N2258)? mem[1778] : 
                       (N2260)? mem[1842] : 
                       (N2262)? mem[1906] : 
                       (N2264)? mem[1970] : 
                       (N2266)? mem[2034] : 1'b0;
  assign rdata_o[49] = (N2235)? mem[49] : 
                       (N2237)? mem[113] : 
                       (N2239)? mem[177] : 
                       (N2241)? mem[241] : 
                       (N2243)? mem[305] : 
                       (N2245)? mem[369] : 
                       (N2247)? mem[433] : 
                       (N2249)? mem[497] : 
                       (N2251)? mem[561] : 
                       (N2253)? mem[625] : 
                       (N2255)? mem[689] : 
                       (N2257)? mem[753] : 
                       (N2259)? mem[817] : 
                       (N2261)? mem[881] : 
                       (N2263)? mem[945] : 
                       (N2265)? mem[1009] : 
                       (N2236)? mem[1073] : 
                       (N2238)? mem[1137] : 
                       (N2240)? mem[1201] : 
                       (N2242)? mem[1265] : 
                       (N2244)? mem[1329] : 
                       (N2246)? mem[1393] : 
                       (N2248)? mem[1457] : 
                       (N2250)? mem[1521] : 
                       (N2252)? mem[1585] : 
                       (N2254)? mem[1649] : 
                       (N2256)? mem[1713] : 
                       (N2258)? mem[1777] : 
                       (N2260)? mem[1841] : 
                       (N2262)? mem[1905] : 
                       (N2264)? mem[1969] : 
                       (N2266)? mem[2033] : 1'b0;
  assign rdata_o[48] = (N2235)? mem[48] : 
                       (N2237)? mem[112] : 
                       (N2239)? mem[176] : 
                       (N2241)? mem[240] : 
                       (N2243)? mem[304] : 
                       (N2245)? mem[368] : 
                       (N2247)? mem[432] : 
                       (N2249)? mem[496] : 
                       (N2251)? mem[560] : 
                       (N2253)? mem[624] : 
                       (N2255)? mem[688] : 
                       (N2257)? mem[752] : 
                       (N2259)? mem[816] : 
                       (N2261)? mem[880] : 
                       (N2263)? mem[944] : 
                       (N2265)? mem[1008] : 
                       (N2236)? mem[1072] : 
                       (N2238)? mem[1136] : 
                       (N2240)? mem[1200] : 
                       (N2242)? mem[1264] : 
                       (N2244)? mem[1328] : 
                       (N2246)? mem[1392] : 
                       (N2248)? mem[1456] : 
                       (N2250)? mem[1520] : 
                       (N2252)? mem[1584] : 
                       (N2254)? mem[1648] : 
                       (N2256)? mem[1712] : 
                       (N2258)? mem[1776] : 
                       (N2260)? mem[1840] : 
                       (N2262)? mem[1904] : 
                       (N2264)? mem[1968] : 
                       (N2266)? mem[2032] : 1'b0;
  assign rdata_o[47] = (N2235)? mem[47] : 
                       (N2237)? mem[111] : 
                       (N2239)? mem[175] : 
                       (N2241)? mem[239] : 
                       (N2243)? mem[303] : 
                       (N2245)? mem[367] : 
                       (N2247)? mem[431] : 
                       (N2249)? mem[495] : 
                       (N2251)? mem[559] : 
                       (N2253)? mem[623] : 
                       (N2255)? mem[687] : 
                       (N2257)? mem[751] : 
                       (N2259)? mem[815] : 
                       (N2261)? mem[879] : 
                       (N2263)? mem[943] : 
                       (N2265)? mem[1007] : 
                       (N2236)? mem[1071] : 
                       (N2238)? mem[1135] : 
                       (N2240)? mem[1199] : 
                       (N2242)? mem[1263] : 
                       (N2244)? mem[1327] : 
                       (N2246)? mem[1391] : 
                       (N2248)? mem[1455] : 
                       (N2250)? mem[1519] : 
                       (N2252)? mem[1583] : 
                       (N2254)? mem[1647] : 
                       (N2256)? mem[1711] : 
                       (N2258)? mem[1775] : 
                       (N2260)? mem[1839] : 
                       (N2262)? mem[1903] : 
                       (N2264)? mem[1967] : 
                       (N2266)? mem[2031] : 1'b0;
  assign rdata_o[46] = (N2235)? mem[46] : 
                       (N2237)? mem[110] : 
                       (N2239)? mem[174] : 
                       (N2241)? mem[238] : 
                       (N2243)? mem[302] : 
                       (N2245)? mem[366] : 
                       (N2247)? mem[430] : 
                       (N2249)? mem[494] : 
                       (N2251)? mem[558] : 
                       (N2253)? mem[622] : 
                       (N2255)? mem[686] : 
                       (N2257)? mem[750] : 
                       (N2259)? mem[814] : 
                       (N2261)? mem[878] : 
                       (N2263)? mem[942] : 
                       (N2265)? mem[1006] : 
                       (N2236)? mem[1070] : 
                       (N2238)? mem[1134] : 
                       (N2240)? mem[1198] : 
                       (N2242)? mem[1262] : 
                       (N2244)? mem[1326] : 
                       (N2246)? mem[1390] : 
                       (N2248)? mem[1454] : 
                       (N2250)? mem[1518] : 
                       (N2252)? mem[1582] : 
                       (N2254)? mem[1646] : 
                       (N2256)? mem[1710] : 
                       (N2258)? mem[1774] : 
                       (N2260)? mem[1838] : 
                       (N2262)? mem[1902] : 
                       (N2264)? mem[1966] : 
                       (N2266)? mem[2030] : 1'b0;
  assign rdata_o[45] = (N2235)? mem[45] : 
                       (N2237)? mem[109] : 
                       (N2239)? mem[173] : 
                       (N2241)? mem[237] : 
                       (N2243)? mem[301] : 
                       (N2245)? mem[365] : 
                       (N2247)? mem[429] : 
                       (N2249)? mem[493] : 
                       (N2251)? mem[557] : 
                       (N2253)? mem[621] : 
                       (N2255)? mem[685] : 
                       (N2257)? mem[749] : 
                       (N2259)? mem[813] : 
                       (N2261)? mem[877] : 
                       (N2263)? mem[941] : 
                       (N2265)? mem[1005] : 
                       (N2236)? mem[1069] : 
                       (N2238)? mem[1133] : 
                       (N2240)? mem[1197] : 
                       (N2242)? mem[1261] : 
                       (N2244)? mem[1325] : 
                       (N2246)? mem[1389] : 
                       (N2248)? mem[1453] : 
                       (N2250)? mem[1517] : 
                       (N2252)? mem[1581] : 
                       (N2254)? mem[1645] : 
                       (N2256)? mem[1709] : 
                       (N2258)? mem[1773] : 
                       (N2260)? mem[1837] : 
                       (N2262)? mem[1901] : 
                       (N2264)? mem[1965] : 
                       (N2266)? mem[2029] : 1'b0;
  assign rdata_o[44] = (N2235)? mem[44] : 
                       (N2237)? mem[108] : 
                       (N2239)? mem[172] : 
                       (N2241)? mem[236] : 
                       (N2243)? mem[300] : 
                       (N2245)? mem[364] : 
                       (N2247)? mem[428] : 
                       (N2249)? mem[492] : 
                       (N2251)? mem[556] : 
                       (N2253)? mem[620] : 
                       (N2255)? mem[684] : 
                       (N2257)? mem[748] : 
                       (N2259)? mem[812] : 
                       (N2261)? mem[876] : 
                       (N2263)? mem[940] : 
                       (N2265)? mem[1004] : 
                       (N2236)? mem[1068] : 
                       (N2238)? mem[1132] : 
                       (N2240)? mem[1196] : 
                       (N2242)? mem[1260] : 
                       (N2244)? mem[1324] : 
                       (N2246)? mem[1388] : 
                       (N2248)? mem[1452] : 
                       (N2250)? mem[1516] : 
                       (N2252)? mem[1580] : 
                       (N2254)? mem[1644] : 
                       (N2256)? mem[1708] : 
                       (N2258)? mem[1772] : 
                       (N2260)? mem[1836] : 
                       (N2262)? mem[1900] : 
                       (N2264)? mem[1964] : 
                       (N2266)? mem[2028] : 1'b0;
  assign rdata_o[43] = (N2235)? mem[43] : 
                       (N2237)? mem[107] : 
                       (N2239)? mem[171] : 
                       (N2241)? mem[235] : 
                       (N2243)? mem[299] : 
                       (N2245)? mem[363] : 
                       (N2247)? mem[427] : 
                       (N2249)? mem[491] : 
                       (N2251)? mem[555] : 
                       (N2253)? mem[619] : 
                       (N2255)? mem[683] : 
                       (N2257)? mem[747] : 
                       (N2259)? mem[811] : 
                       (N2261)? mem[875] : 
                       (N2263)? mem[939] : 
                       (N2265)? mem[1003] : 
                       (N2236)? mem[1067] : 
                       (N2238)? mem[1131] : 
                       (N2240)? mem[1195] : 
                       (N2242)? mem[1259] : 
                       (N2244)? mem[1323] : 
                       (N2246)? mem[1387] : 
                       (N2248)? mem[1451] : 
                       (N2250)? mem[1515] : 
                       (N2252)? mem[1579] : 
                       (N2254)? mem[1643] : 
                       (N2256)? mem[1707] : 
                       (N2258)? mem[1771] : 
                       (N2260)? mem[1835] : 
                       (N2262)? mem[1899] : 
                       (N2264)? mem[1963] : 
                       (N2266)? mem[2027] : 1'b0;
  assign rdata_o[42] = (N2235)? mem[42] : 
                       (N2237)? mem[106] : 
                       (N2239)? mem[170] : 
                       (N2241)? mem[234] : 
                       (N2243)? mem[298] : 
                       (N2245)? mem[362] : 
                       (N2247)? mem[426] : 
                       (N2249)? mem[490] : 
                       (N2251)? mem[554] : 
                       (N2253)? mem[618] : 
                       (N2255)? mem[682] : 
                       (N2257)? mem[746] : 
                       (N2259)? mem[810] : 
                       (N2261)? mem[874] : 
                       (N2263)? mem[938] : 
                       (N2265)? mem[1002] : 
                       (N2236)? mem[1066] : 
                       (N2238)? mem[1130] : 
                       (N2240)? mem[1194] : 
                       (N2242)? mem[1258] : 
                       (N2244)? mem[1322] : 
                       (N2246)? mem[1386] : 
                       (N2248)? mem[1450] : 
                       (N2250)? mem[1514] : 
                       (N2252)? mem[1578] : 
                       (N2254)? mem[1642] : 
                       (N2256)? mem[1706] : 
                       (N2258)? mem[1770] : 
                       (N2260)? mem[1834] : 
                       (N2262)? mem[1898] : 
                       (N2264)? mem[1962] : 
                       (N2266)? mem[2026] : 1'b0;
  assign rdata_o[41] = (N2235)? mem[41] : 
                       (N2237)? mem[105] : 
                       (N2239)? mem[169] : 
                       (N2241)? mem[233] : 
                       (N2243)? mem[297] : 
                       (N2245)? mem[361] : 
                       (N2247)? mem[425] : 
                       (N2249)? mem[489] : 
                       (N2251)? mem[553] : 
                       (N2253)? mem[617] : 
                       (N2255)? mem[681] : 
                       (N2257)? mem[745] : 
                       (N2259)? mem[809] : 
                       (N2261)? mem[873] : 
                       (N2263)? mem[937] : 
                       (N2265)? mem[1001] : 
                       (N2236)? mem[1065] : 
                       (N2238)? mem[1129] : 
                       (N2240)? mem[1193] : 
                       (N2242)? mem[1257] : 
                       (N2244)? mem[1321] : 
                       (N2246)? mem[1385] : 
                       (N2248)? mem[1449] : 
                       (N2250)? mem[1513] : 
                       (N2252)? mem[1577] : 
                       (N2254)? mem[1641] : 
                       (N2256)? mem[1705] : 
                       (N2258)? mem[1769] : 
                       (N2260)? mem[1833] : 
                       (N2262)? mem[1897] : 
                       (N2264)? mem[1961] : 
                       (N2266)? mem[2025] : 1'b0;
  assign rdata_o[40] = (N2235)? mem[40] : 
                       (N2237)? mem[104] : 
                       (N2239)? mem[168] : 
                       (N2241)? mem[232] : 
                       (N2243)? mem[296] : 
                       (N2245)? mem[360] : 
                       (N2247)? mem[424] : 
                       (N2249)? mem[488] : 
                       (N2251)? mem[552] : 
                       (N2253)? mem[616] : 
                       (N2255)? mem[680] : 
                       (N2257)? mem[744] : 
                       (N2259)? mem[808] : 
                       (N2261)? mem[872] : 
                       (N2263)? mem[936] : 
                       (N2265)? mem[1000] : 
                       (N2236)? mem[1064] : 
                       (N2238)? mem[1128] : 
                       (N2240)? mem[1192] : 
                       (N2242)? mem[1256] : 
                       (N2244)? mem[1320] : 
                       (N2246)? mem[1384] : 
                       (N2248)? mem[1448] : 
                       (N2250)? mem[1512] : 
                       (N2252)? mem[1576] : 
                       (N2254)? mem[1640] : 
                       (N2256)? mem[1704] : 
                       (N2258)? mem[1768] : 
                       (N2260)? mem[1832] : 
                       (N2262)? mem[1896] : 
                       (N2264)? mem[1960] : 
                       (N2266)? mem[2024] : 1'b0;
  assign rdata_o[39] = (N2235)? mem[39] : 
                       (N2237)? mem[103] : 
                       (N2239)? mem[167] : 
                       (N2241)? mem[231] : 
                       (N2243)? mem[295] : 
                       (N2245)? mem[359] : 
                       (N2247)? mem[423] : 
                       (N2249)? mem[487] : 
                       (N2251)? mem[551] : 
                       (N2253)? mem[615] : 
                       (N2255)? mem[679] : 
                       (N2257)? mem[743] : 
                       (N2259)? mem[807] : 
                       (N2261)? mem[871] : 
                       (N2263)? mem[935] : 
                       (N2265)? mem[999] : 
                       (N2236)? mem[1063] : 
                       (N2238)? mem[1127] : 
                       (N2240)? mem[1191] : 
                       (N2242)? mem[1255] : 
                       (N2244)? mem[1319] : 
                       (N2246)? mem[1383] : 
                       (N2248)? mem[1447] : 
                       (N2250)? mem[1511] : 
                       (N2252)? mem[1575] : 
                       (N2254)? mem[1639] : 
                       (N2256)? mem[1703] : 
                       (N2258)? mem[1767] : 
                       (N2260)? mem[1831] : 
                       (N2262)? mem[1895] : 
                       (N2264)? mem[1959] : 
                       (N2266)? mem[2023] : 1'b0;
  assign rdata_o[38] = (N2235)? mem[38] : 
                       (N2237)? mem[102] : 
                       (N2239)? mem[166] : 
                       (N2241)? mem[230] : 
                       (N2243)? mem[294] : 
                       (N2245)? mem[358] : 
                       (N2247)? mem[422] : 
                       (N2249)? mem[486] : 
                       (N2251)? mem[550] : 
                       (N2253)? mem[614] : 
                       (N2255)? mem[678] : 
                       (N2257)? mem[742] : 
                       (N2259)? mem[806] : 
                       (N2261)? mem[870] : 
                       (N2263)? mem[934] : 
                       (N2265)? mem[998] : 
                       (N2236)? mem[1062] : 
                       (N2238)? mem[1126] : 
                       (N2240)? mem[1190] : 
                       (N2242)? mem[1254] : 
                       (N2244)? mem[1318] : 
                       (N2246)? mem[1382] : 
                       (N2248)? mem[1446] : 
                       (N2250)? mem[1510] : 
                       (N2252)? mem[1574] : 
                       (N2254)? mem[1638] : 
                       (N2256)? mem[1702] : 
                       (N2258)? mem[1766] : 
                       (N2260)? mem[1830] : 
                       (N2262)? mem[1894] : 
                       (N2264)? mem[1958] : 
                       (N2266)? mem[2022] : 1'b0;
  assign rdata_o[37] = (N2235)? mem[37] : 
                       (N2237)? mem[101] : 
                       (N2239)? mem[165] : 
                       (N2241)? mem[229] : 
                       (N2243)? mem[293] : 
                       (N2245)? mem[357] : 
                       (N2247)? mem[421] : 
                       (N2249)? mem[485] : 
                       (N2251)? mem[549] : 
                       (N2253)? mem[613] : 
                       (N2255)? mem[677] : 
                       (N2257)? mem[741] : 
                       (N2259)? mem[805] : 
                       (N2261)? mem[869] : 
                       (N2263)? mem[933] : 
                       (N2265)? mem[997] : 
                       (N2236)? mem[1061] : 
                       (N2238)? mem[1125] : 
                       (N2240)? mem[1189] : 
                       (N2242)? mem[1253] : 
                       (N2244)? mem[1317] : 
                       (N2246)? mem[1381] : 
                       (N2248)? mem[1445] : 
                       (N2250)? mem[1509] : 
                       (N2252)? mem[1573] : 
                       (N2254)? mem[1637] : 
                       (N2256)? mem[1701] : 
                       (N2258)? mem[1765] : 
                       (N2260)? mem[1829] : 
                       (N2262)? mem[1893] : 
                       (N2264)? mem[1957] : 
                       (N2266)? mem[2021] : 1'b0;
  assign rdata_o[36] = (N2235)? mem[36] : 
                       (N2237)? mem[100] : 
                       (N2239)? mem[164] : 
                       (N2241)? mem[228] : 
                       (N2243)? mem[292] : 
                       (N2245)? mem[356] : 
                       (N2247)? mem[420] : 
                       (N2249)? mem[484] : 
                       (N2251)? mem[548] : 
                       (N2253)? mem[612] : 
                       (N2255)? mem[676] : 
                       (N2257)? mem[740] : 
                       (N2259)? mem[804] : 
                       (N2261)? mem[868] : 
                       (N2263)? mem[932] : 
                       (N2265)? mem[996] : 
                       (N2236)? mem[1060] : 
                       (N2238)? mem[1124] : 
                       (N2240)? mem[1188] : 
                       (N2242)? mem[1252] : 
                       (N2244)? mem[1316] : 
                       (N2246)? mem[1380] : 
                       (N2248)? mem[1444] : 
                       (N2250)? mem[1508] : 
                       (N2252)? mem[1572] : 
                       (N2254)? mem[1636] : 
                       (N2256)? mem[1700] : 
                       (N2258)? mem[1764] : 
                       (N2260)? mem[1828] : 
                       (N2262)? mem[1892] : 
                       (N2264)? mem[1956] : 
                       (N2266)? mem[2020] : 1'b0;
  assign rdata_o[35] = (N2235)? mem[35] : 
                       (N2237)? mem[99] : 
                       (N2239)? mem[163] : 
                       (N2241)? mem[227] : 
                       (N2243)? mem[291] : 
                       (N2245)? mem[355] : 
                       (N2247)? mem[419] : 
                       (N2249)? mem[483] : 
                       (N2251)? mem[547] : 
                       (N2253)? mem[611] : 
                       (N2255)? mem[675] : 
                       (N2257)? mem[739] : 
                       (N2259)? mem[803] : 
                       (N2261)? mem[867] : 
                       (N2263)? mem[931] : 
                       (N2265)? mem[995] : 
                       (N2236)? mem[1059] : 
                       (N2238)? mem[1123] : 
                       (N2240)? mem[1187] : 
                       (N2242)? mem[1251] : 
                       (N2244)? mem[1315] : 
                       (N2246)? mem[1379] : 
                       (N2248)? mem[1443] : 
                       (N2250)? mem[1507] : 
                       (N2252)? mem[1571] : 
                       (N2254)? mem[1635] : 
                       (N2256)? mem[1699] : 
                       (N2258)? mem[1763] : 
                       (N2260)? mem[1827] : 
                       (N2262)? mem[1891] : 
                       (N2264)? mem[1955] : 
                       (N2266)? mem[2019] : 1'b0;
  assign rdata_o[34] = (N2235)? mem[34] : 
                       (N2237)? mem[98] : 
                       (N2239)? mem[162] : 
                       (N2241)? mem[226] : 
                       (N2243)? mem[290] : 
                       (N2245)? mem[354] : 
                       (N2247)? mem[418] : 
                       (N2249)? mem[482] : 
                       (N2251)? mem[546] : 
                       (N2253)? mem[610] : 
                       (N2255)? mem[674] : 
                       (N2257)? mem[738] : 
                       (N2259)? mem[802] : 
                       (N2261)? mem[866] : 
                       (N2263)? mem[930] : 
                       (N2265)? mem[994] : 
                       (N2236)? mem[1058] : 
                       (N2238)? mem[1122] : 
                       (N2240)? mem[1186] : 
                       (N2242)? mem[1250] : 
                       (N2244)? mem[1314] : 
                       (N2246)? mem[1378] : 
                       (N2248)? mem[1442] : 
                       (N2250)? mem[1506] : 
                       (N2252)? mem[1570] : 
                       (N2254)? mem[1634] : 
                       (N2256)? mem[1698] : 
                       (N2258)? mem[1762] : 
                       (N2260)? mem[1826] : 
                       (N2262)? mem[1890] : 
                       (N2264)? mem[1954] : 
                       (N2266)? mem[2018] : 1'b0;
  assign rdata_o[33] = (N2235)? mem[33] : 
                       (N2237)? mem[97] : 
                       (N2239)? mem[161] : 
                       (N2241)? mem[225] : 
                       (N2243)? mem[289] : 
                       (N2245)? mem[353] : 
                       (N2247)? mem[417] : 
                       (N2249)? mem[481] : 
                       (N2251)? mem[545] : 
                       (N2253)? mem[609] : 
                       (N2255)? mem[673] : 
                       (N2257)? mem[737] : 
                       (N2259)? mem[801] : 
                       (N2261)? mem[865] : 
                       (N2263)? mem[929] : 
                       (N2265)? mem[993] : 
                       (N2236)? mem[1057] : 
                       (N2238)? mem[1121] : 
                       (N2240)? mem[1185] : 
                       (N2242)? mem[1249] : 
                       (N2244)? mem[1313] : 
                       (N2246)? mem[1377] : 
                       (N2248)? mem[1441] : 
                       (N2250)? mem[1505] : 
                       (N2252)? mem[1569] : 
                       (N2254)? mem[1633] : 
                       (N2256)? mem[1697] : 
                       (N2258)? mem[1761] : 
                       (N2260)? mem[1825] : 
                       (N2262)? mem[1889] : 
                       (N2264)? mem[1953] : 
                       (N2266)? mem[2017] : 1'b0;
  assign rdata_o[32] = (N2235)? mem[32] : 
                       (N2237)? mem[96] : 
                       (N2239)? mem[160] : 
                       (N2241)? mem[224] : 
                       (N2243)? mem[288] : 
                       (N2245)? mem[352] : 
                       (N2247)? mem[416] : 
                       (N2249)? mem[480] : 
                       (N2251)? mem[544] : 
                       (N2253)? mem[608] : 
                       (N2255)? mem[672] : 
                       (N2257)? mem[736] : 
                       (N2259)? mem[800] : 
                       (N2261)? mem[864] : 
                       (N2263)? mem[928] : 
                       (N2265)? mem[992] : 
                       (N2236)? mem[1056] : 
                       (N2238)? mem[1120] : 
                       (N2240)? mem[1184] : 
                       (N2242)? mem[1248] : 
                       (N2244)? mem[1312] : 
                       (N2246)? mem[1376] : 
                       (N2248)? mem[1440] : 
                       (N2250)? mem[1504] : 
                       (N2252)? mem[1568] : 
                       (N2254)? mem[1632] : 
                       (N2256)? mem[1696] : 
                       (N2258)? mem[1760] : 
                       (N2260)? mem[1824] : 
                       (N2262)? mem[1888] : 
                       (N2264)? mem[1952] : 
                       (N2266)? mem[2016] : 1'b0;
  assign rdata_o[31] = (N2235)? mem[31] : 
                       (N2237)? mem[95] : 
                       (N2239)? mem[159] : 
                       (N2241)? mem[223] : 
                       (N2243)? mem[287] : 
                       (N2245)? mem[351] : 
                       (N2247)? mem[415] : 
                       (N2249)? mem[479] : 
                       (N2251)? mem[543] : 
                       (N2253)? mem[607] : 
                       (N2255)? mem[671] : 
                       (N2257)? mem[735] : 
                       (N2259)? mem[799] : 
                       (N2261)? mem[863] : 
                       (N2263)? mem[927] : 
                       (N2265)? mem[991] : 
                       (N2236)? mem[1055] : 
                       (N2238)? mem[1119] : 
                       (N2240)? mem[1183] : 
                       (N2242)? mem[1247] : 
                       (N2244)? mem[1311] : 
                       (N2246)? mem[1375] : 
                       (N2248)? mem[1439] : 
                       (N2250)? mem[1503] : 
                       (N2252)? mem[1567] : 
                       (N2254)? mem[1631] : 
                       (N2256)? mem[1695] : 
                       (N2258)? mem[1759] : 
                       (N2260)? mem[1823] : 
                       (N2262)? mem[1887] : 
                       (N2264)? mem[1951] : 
                       (N2266)? mem[2015] : 1'b0;
  assign rdata_o[30] = (N2235)? mem[30] : 
                       (N2237)? mem[94] : 
                       (N2239)? mem[158] : 
                       (N2241)? mem[222] : 
                       (N2243)? mem[286] : 
                       (N2245)? mem[350] : 
                       (N2247)? mem[414] : 
                       (N2249)? mem[478] : 
                       (N2251)? mem[542] : 
                       (N2253)? mem[606] : 
                       (N2255)? mem[670] : 
                       (N2257)? mem[734] : 
                       (N2259)? mem[798] : 
                       (N2261)? mem[862] : 
                       (N2263)? mem[926] : 
                       (N2265)? mem[990] : 
                       (N2236)? mem[1054] : 
                       (N2238)? mem[1118] : 
                       (N2240)? mem[1182] : 
                       (N2242)? mem[1246] : 
                       (N2244)? mem[1310] : 
                       (N2246)? mem[1374] : 
                       (N2248)? mem[1438] : 
                       (N2250)? mem[1502] : 
                       (N2252)? mem[1566] : 
                       (N2254)? mem[1630] : 
                       (N2256)? mem[1694] : 
                       (N2258)? mem[1758] : 
                       (N2260)? mem[1822] : 
                       (N2262)? mem[1886] : 
                       (N2264)? mem[1950] : 
                       (N2266)? mem[2014] : 1'b0;
  assign rdata_o[29] = (N2235)? mem[29] : 
                       (N2237)? mem[93] : 
                       (N2239)? mem[157] : 
                       (N2241)? mem[221] : 
                       (N2243)? mem[285] : 
                       (N2245)? mem[349] : 
                       (N2247)? mem[413] : 
                       (N2249)? mem[477] : 
                       (N2251)? mem[541] : 
                       (N2253)? mem[605] : 
                       (N2255)? mem[669] : 
                       (N2257)? mem[733] : 
                       (N2259)? mem[797] : 
                       (N2261)? mem[861] : 
                       (N2263)? mem[925] : 
                       (N2265)? mem[989] : 
                       (N2236)? mem[1053] : 
                       (N2238)? mem[1117] : 
                       (N2240)? mem[1181] : 
                       (N2242)? mem[1245] : 
                       (N2244)? mem[1309] : 
                       (N2246)? mem[1373] : 
                       (N2248)? mem[1437] : 
                       (N2250)? mem[1501] : 
                       (N2252)? mem[1565] : 
                       (N2254)? mem[1629] : 
                       (N2256)? mem[1693] : 
                       (N2258)? mem[1757] : 
                       (N2260)? mem[1821] : 
                       (N2262)? mem[1885] : 
                       (N2264)? mem[1949] : 
                       (N2266)? mem[2013] : 1'b0;
  assign rdata_o[28] = (N2235)? mem[28] : 
                       (N2237)? mem[92] : 
                       (N2239)? mem[156] : 
                       (N2241)? mem[220] : 
                       (N2243)? mem[284] : 
                       (N2245)? mem[348] : 
                       (N2247)? mem[412] : 
                       (N2249)? mem[476] : 
                       (N2251)? mem[540] : 
                       (N2253)? mem[604] : 
                       (N2255)? mem[668] : 
                       (N2257)? mem[732] : 
                       (N2259)? mem[796] : 
                       (N2261)? mem[860] : 
                       (N2263)? mem[924] : 
                       (N2265)? mem[988] : 
                       (N2236)? mem[1052] : 
                       (N2238)? mem[1116] : 
                       (N2240)? mem[1180] : 
                       (N2242)? mem[1244] : 
                       (N2244)? mem[1308] : 
                       (N2246)? mem[1372] : 
                       (N2248)? mem[1436] : 
                       (N2250)? mem[1500] : 
                       (N2252)? mem[1564] : 
                       (N2254)? mem[1628] : 
                       (N2256)? mem[1692] : 
                       (N2258)? mem[1756] : 
                       (N2260)? mem[1820] : 
                       (N2262)? mem[1884] : 
                       (N2264)? mem[1948] : 
                       (N2266)? mem[2012] : 1'b0;
  assign rdata_o[27] = (N2235)? mem[27] : 
                       (N2237)? mem[91] : 
                       (N2239)? mem[155] : 
                       (N2241)? mem[219] : 
                       (N2243)? mem[283] : 
                       (N2245)? mem[347] : 
                       (N2247)? mem[411] : 
                       (N2249)? mem[475] : 
                       (N2251)? mem[539] : 
                       (N2253)? mem[603] : 
                       (N2255)? mem[667] : 
                       (N2257)? mem[731] : 
                       (N2259)? mem[795] : 
                       (N2261)? mem[859] : 
                       (N2263)? mem[923] : 
                       (N2265)? mem[987] : 
                       (N2236)? mem[1051] : 
                       (N2238)? mem[1115] : 
                       (N2240)? mem[1179] : 
                       (N2242)? mem[1243] : 
                       (N2244)? mem[1307] : 
                       (N2246)? mem[1371] : 
                       (N2248)? mem[1435] : 
                       (N2250)? mem[1499] : 
                       (N2252)? mem[1563] : 
                       (N2254)? mem[1627] : 
                       (N2256)? mem[1691] : 
                       (N2258)? mem[1755] : 
                       (N2260)? mem[1819] : 
                       (N2262)? mem[1883] : 
                       (N2264)? mem[1947] : 
                       (N2266)? mem[2011] : 1'b0;
  assign rdata_o[26] = (N2235)? mem[26] : 
                       (N2237)? mem[90] : 
                       (N2239)? mem[154] : 
                       (N2241)? mem[218] : 
                       (N2243)? mem[282] : 
                       (N2245)? mem[346] : 
                       (N2247)? mem[410] : 
                       (N2249)? mem[474] : 
                       (N2251)? mem[538] : 
                       (N2253)? mem[602] : 
                       (N2255)? mem[666] : 
                       (N2257)? mem[730] : 
                       (N2259)? mem[794] : 
                       (N2261)? mem[858] : 
                       (N2263)? mem[922] : 
                       (N2265)? mem[986] : 
                       (N2236)? mem[1050] : 
                       (N2238)? mem[1114] : 
                       (N2240)? mem[1178] : 
                       (N2242)? mem[1242] : 
                       (N2244)? mem[1306] : 
                       (N2246)? mem[1370] : 
                       (N2248)? mem[1434] : 
                       (N2250)? mem[1498] : 
                       (N2252)? mem[1562] : 
                       (N2254)? mem[1626] : 
                       (N2256)? mem[1690] : 
                       (N2258)? mem[1754] : 
                       (N2260)? mem[1818] : 
                       (N2262)? mem[1882] : 
                       (N2264)? mem[1946] : 
                       (N2266)? mem[2010] : 1'b0;
  assign rdata_o[25] = (N2235)? mem[25] : 
                       (N2237)? mem[89] : 
                       (N2239)? mem[153] : 
                       (N2241)? mem[217] : 
                       (N2243)? mem[281] : 
                       (N2245)? mem[345] : 
                       (N2247)? mem[409] : 
                       (N2249)? mem[473] : 
                       (N2251)? mem[537] : 
                       (N2253)? mem[601] : 
                       (N2255)? mem[665] : 
                       (N2257)? mem[729] : 
                       (N2259)? mem[793] : 
                       (N2261)? mem[857] : 
                       (N2263)? mem[921] : 
                       (N2265)? mem[985] : 
                       (N2236)? mem[1049] : 
                       (N2238)? mem[1113] : 
                       (N2240)? mem[1177] : 
                       (N2242)? mem[1241] : 
                       (N2244)? mem[1305] : 
                       (N2246)? mem[1369] : 
                       (N2248)? mem[1433] : 
                       (N2250)? mem[1497] : 
                       (N2252)? mem[1561] : 
                       (N2254)? mem[1625] : 
                       (N2256)? mem[1689] : 
                       (N2258)? mem[1753] : 
                       (N2260)? mem[1817] : 
                       (N2262)? mem[1881] : 
                       (N2264)? mem[1945] : 
                       (N2266)? mem[2009] : 1'b0;
  assign rdata_o[24] = (N2235)? mem[24] : 
                       (N2237)? mem[88] : 
                       (N2239)? mem[152] : 
                       (N2241)? mem[216] : 
                       (N2243)? mem[280] : 
                       (N2245)? mem[344] : 
                       (N2247)? mem[408] : 
                       (N2249)? mem[472] : 
                       (N2251)? mem[536] : 
                       (N2253)? mem[600] : 
                       (N2255)? mem[664] : 
                       (N2257)? mem[728] : 
                       (N2259)? mem[792] : 
                       (N2261)? mem[856] : 
                       (N2263)? mem[920] : 
                       (N2265)? mem[984] : 
                       (N2236)? mem[1048] : 
                       (N2238)? mem[1112] : 
                       (N2240)? mem[1176] : 
                       (N2242)? mem[1240] : 
                       (N2244)? mem[1304] : 
                       (N2246)? mem[1368] : 
                       (N2248)? mem[1432] : 
                       (N2250)? mem[1496] : 
                       (N2252)? mem[1560] : 
                       (N2254)? mem[1624] : 
                       (N2256)? mem[1688] : 
                       (N2258)? mem[1752] : 
                       (N2260)? mem[1816] : 
                       (N2262)? mem[1880] : 
                       (N2264)? mem[1944] : 
                       (N2266)? mem[2008] : 1'b0;
  assign rdata_o[23] = (N2235)? mem[23] : 
                       (N2237)? mem[87] : 
                       (N2239)? mem[151] : 
                       (N2241)? mem[215] : 
                       (N2243)? mem[279] : 
                       (N2245)? mem[343] : 
                       (N2247)? mem[407] : 
                       (N2249)? mem[471] : 
                       (N2251)? mem[535] : 
                       (N2253)? mem[599] : 
                       (N2255)? mem[663] : 
                       (N2257)? mem[727] : 
                       (N2259)? mem[791] : 
                       (N2261)? mem[855] : 
                       (N2263)? mem[919] : 
                       (N2265)? mem[983] : 
                       (N2236)? mem[1047] : 
                       (N2238)? mem[1111] : 
                       (N2240)? mem[1175] : 
                       (N2242)? mem[1239] : 
                       (N2244)? mem[1303] : 
                       (N2246)? mem[1367] : 
                       (N2248)? mem[1431] : 
                       (N2250)? mem[1495] : 
                       (N2252)? mem[1559] : 
                       (N2254)? mem[1623] : 
                       (N2256)? mem[1687] : 
                       (N2258)? mem[1751] : 
                       (N2260)? mem[1815] : 
                       (N2262)? mem[1879] : 
                       (N2264)? mem[1943] : 
                       (N2266)? mem[2007] : 1'b0;
  assign rdata_o[22] = (N2235)? mem[22] : 
                       (N2237)? mem[86] : 
                       (N2239)? mem[150] : 
                       (N2241)? mem[214] : 
                       (N2243)? mem[278] : 
                       (N2245)? mem[342] : 
                       (N2247)? mem[406] : 
                       (N2249)? mem[470] : 
                       (N2251)? mem[534] : 
                       (N2253)? mem[598] : 
                       (N2255)? mem[662] : 
                       (N2257)? mem[726] : 
                       (N2259)? mem[790] : 
                       (N2261)? mem[854] : 
                       (N2263)? mem[918] : 
                       (N2265)? mem[982] : 
                       (N2236)? mem[1046] : 
                       (N2238)? mem[1110] : 
                       (N2240)? mem[1174] : 
                       (N2242)? mem[1238] : 
                       (N2244)? mem[1302] : 
                       (N2246)? mem[1366] : 
                       (N2248)? mem[1430] : 
                       (N2250)? mem[1494] : 
                       (N2252)? mem[1558] : 
                       (N2254)? mem[1622] : 
                       (N2256)? mem[1686] : 
                       (N2258)? mem[1750] : 
                       (N2260)? mem[1814] : 
                       (N2262)? mem[1878] : 
                       (N2264)? mem[1942] : 
                       (N2266)? mem[2006] : 1'b0;
  assign rdata_o[21] = (N2235)? mem[21] : 
                       (N2237)? mem[85] : 
                       (N2239)? mem[149] : 
                       (N2241)? mem[213] : 
                       (N2243)? mem[277] : 
                       (N2245)? mem[341] : 
                       (N2247)? mem[405] : 
                       (N2249)? mem[469] : 
                       (N2251)? mem[533] : 
                       (N2253)? mem[597] : 
                       (N2255)? mem[661] : 
                       (N2257)? mem[725] : 
                       (N2259)? mem[789] : 
                       (N2261)? mem[853] : 
                       (N2263)? mem[917] : 
                       (N2265)? mem[981] : 
                       (N2236)? mem[1045] : 
                       (N2238)? mem[1109] : 
                       (N2240)? mem[1173] : 
                       (N2242)? mem[1237] : 
                       (N2244)? mem[1301] : 
                       (N2246)? mem[1365] : 
                       (N2248)? mem[1429] : 
                       (N2250)? mem[1493] : 
                       (N2252)? mem[1557] : 
                       (N2254)? mem[1621] : 
                       (N2256)? mem[1685] : 
                       (N2258)? mem[1749] : 
                       (N2260)? mem[1813] : 
                       (N2262)? mem[1877] : 
                       (N2264)? mem[1941] : 
                       (N2266)? mem[2005] : 1'b0;
  assign rdata_o[20] = (N2235)? mem[20] : 
                       (N2237)? mem[84] : 
                       (N2239)? mem[148] : 
                       (N2241)? mem[212] : 
                       (N2243)? mem[276] : 
                       (N2245)? mem[340] : 
                       (N2247)? mem[404] : 
                       (N2249)? mem[468] : 
                       (N2251)? mem[532] : 
                       (N2253)? mem[596] : 
                       (N2255)? mem[660] : 
                       (N2257)? mem[724] : 
                       (N2259)? mem[788] : 
                       (N2261)? mem[852] : 
                       (N2263)? mem[916] : 
                       (N2265)? mem[980] : 
                       (N2236)? mem[1044] : 
                       (N2238)? mem[1108] : 
                       (N2240)? mem[1172] : 
                       (N2242)? mem[1236] : 
                       (N2244)? mem[1300] : 
                       (N2246)? mem[1364] : 
                       (N2248)? mem[1428] : 
                       (N2250)? mem[1492] : 
                       (N2252)? mem[1556] : 
                       (N2254)? mem[1620] : 
                       (N2256)? mem[1684] : 
                       (N2258)? mem[1748] : 
                       (N2260)? mem[1812] : 
                       (N2262)? mem[1876] : 
                       (N2264)? mem[1940] : 
                       (N2266)? mem[2004] : 1'b0;
  assign rdata_o[19] = (N2235)? mem[19] : 
                       (N2237)? mem[83] : 
                       (N2239)? mem[147] : 
                       (N2241)? mem[211] : 
                       (N2243)? mem[275] : 
                       (N2245)? mem[339] : 
                       (N2247)? mem[403] : 
                       (N2249)? mem[467] : 
                       (N2251)? mem[531] : 
                       (N2253)? mem[595] : 
                       (N2255)? mem[659] : 
                       (N2257)? mem[723] : 
                       (N2259)? mem[787] : 
                       (N2261)? mem[851] : 
                       (N2263)? mem[915] : 
                       (N2265)? mem[979] : 
                       (N2236)? mem[1043] : 
                       (N2238)? mem[1107] : 
                       (N2240)? mem[1171] : 
                       (N2242)? mem[1235] : 
                       (N2244)? mem[1299] : 
                       (N2246)? mem[1363] : 
                       (N2248)? mem[1427] : 
                       (N2250)? mem[1491] : 
                       (N2252)? mem[1555] : 
                       (N2254)? mem[1619] : 
                       (N2256)? mem[1683] : 
                       (N2258)? mem[1747] : 
                       (N2260)? mem[1811] : 
                       (N2262)? mem[1875] : 
                       (N2264)? mem[1939] : 
                       (N2266)? mem[2003] : 1'b0;
  assign rdata_o[18] = (N2235)? mem[18] : 
                       (N2237)? mem[82] : 
                       (N2239)? mem[146] : 
                       (N2241)? mem[210] : 
                       (N2243)? mem[274] : 
                       (N2245)? mem[338] : 
                       (N2247)? mem[402] : 
                       (N2249)? mem[466] : 
                       (N2251)? mem[530] : 
                       (N2253)? mem[594] : 
                       (N2255)? mem[658] : 
                       (N2257)? mem[722] : 
                       (N2259)? mem[786] : 
                       (N2261)? mem[850] : 
                       (N2263)? mem[914] : 
                       (N2265)? mem[978] : 
                       (N2236)? mem[1042] : 
                       (N2238)? mem[1106] : 
                       (N2240)? mem[1170] : 
                       (N2242)? mem[1234] : 
                       (N2244)? mem[1298] : 
                       (N2246)? mem[1362] : 
                       (N2248)? mem[1426] : 
                       (N2250)? mem[1490] : 
                       (N2252)? mem[1554] : 
                       (N2254)? mem[1618] : 
                       (N2256)? mem[1682] : 
                       (N2258)? mem[1746] : 
                       (N2260)? mem[1810] : 
                       (N2262)? mem[1874] : 
                       (N2264)? mem[1938] : 
                       (N2266)? mem[2002] : 1'b0;
  assign rdata_o[17] = (N2235)? mem[17] : 
                       (N2237)? mem[81] : 
                       (N2239)? mem[145] : 
                       (N2241)? mem[209] : 
                       (N2243)? mem[273] : 
                       (N2245)? mem[337] : 
                       (N2247)? mem[401] : 
                       (N2249)? mem[465] : 
                       (N2251)? mem[529] : 
                       (N2253)? mem[593] : 
                       (N2255)? mem[657] : 
                       (N2257)? mem[721] : 
                       (N2259)? mem[785] : 
                       (N2261)? mem[849] : 
                       (N2263)? mem[913] : 
                       (N2265)? mem[977] : 
                       (N2236)? mem[1041] : 
                       (N2238)? mem[1105] : 
                       (N2240)? mem[1169] : 
                       (N2242)? mem[1233] : 
                       (N2244)? mem[1297] : 
                       (N2246)? mem[1361] : 
                       (N2248)? mem[1425] : 
                       (N2250)? mem[1489] : 
                       (N2252)? mem[1553] : 
                       (N2254)? mem[1617] : 
                       (N2256)? mem[1681] : 
                       (N2258)? mem[1745] : 
                       (N2260)? mem[1809] : 
                       (N2262)? mem[1873] : 
                       (N2264)? mem[1937] : 
                       (N2266)? mem[2001] : 1'b0;
  assign rdata_o[16] = (N2235)? mem[16] : 
                       (N2237)? mem[80] : 
                       (N2239)? mem[144] : 
                       (N2241)? mem[208] : 
                       (N2243)? mem[272] : 
                       (N2245)? mem[336] : 
                       (N2247)? mem[400] : 
                       (N2249)? mem[464] : 
                       (N2251)? mem[528] : 
                       (N2253)? mem[592] : 
                       (N2255)? mem[656] : 
                       (N2257)? mem[720] : 
                       (N2259)? mem[784] : 
                       (N2261)? mem[848] : 
                       (N2263)? mem[912] : 
                       (N2265)? mem[976] : 
                       (N2236)? mem[1040] : 
                       (N2238)? mem[1104] : 
                       (N2240)? mem[1168] : 
                       (N2242)? mem[1232] : 
                       (N2244)? mem[1296] : 
                       (N2246)? mem[1360] : 
                       (N2248)? mem[1424] : 
                       (N2250)? mem[1488] : 
                       (N2252)? mem[1552] : 
                       (N2254)? mem[1616] : 
                       (N2256)? mem[1680] : 
                       (N2258)? mem[1744] : 
                       (N2260)? mem[1808] : 
                       (N2262)? mem[1872] : 
                       (N2264)? mem[1936] : 
                       (N2266)? mem[2000] : 1'b0;
  assign rdata_o[15] = (N2235)? mem[15] : 
                       (N2237)? mem[79] : 
                       (N2239)? mem[143] : 
                       (N2241)? mem[207] : 
                       (N2243)? mem[271] : 
                       (N2245)? mem[335] : 
                       (N2247)? mem[399] : 
                       (N2249)? mem[463] : 
                       (N2251)? mem[527] : 
                       (N2253)? mem[591] : 
                       (N2255)? mem[655] : 
                       (N2257)? mem[719] : 
                       (N2259)? mem[783] : 
                       (N2261)? mem[847] : 
                       (N2263)? mem[911] : 
                       (N2265)? mem[975] : 
                       (N2236)? mem[1039] : 
                       (N2238)? mem[1103] : 
                       (N2240)? mem[1167] : 
                       (N2242)? mem[1231] : 
                       (N2244)? mem[1295] : 
                       (N2246)? mem[1359] : 
                       (N2248)? mem[1423] : 
                       (N2250)? mem[1487] : 
                       (N2252)? mem[1551] : 
                       (N2254)? mem[1615] : 
                       (N2256)? mem[1679] : 
                       (N2258)? mem[1743] : 
                       (N2260)? mem[1807] : 
                       (N2262)? mem[1871] : 
                       (N2264)? mem[1935] : 
                       (N2266)? mem[1999] : 1'b0;
  assign rdata_o[14] = (N2235)? mem[14] : 
                       (N2237)? mem[78] : 
                       (N2239)? mem[142] : 
                       (N2241)? mem[206] : 
                       (N2243)? mem[270] : 
                       (N2245)? mem[334] : 
                       (N2247)? mem[398] : 
                       (N2249)? mem[462] : 
                       (N2251)? mem[526] : 
                       (N2253)? mem[590] : 
                       (N2255)? mem[654] : 
                       (N2257)? mem[718] : 
                       (N2259)? mem[782] : 
                       (N2261)? mem[846] : 
                       (N2263)? mem[910] : 
                       (N2265)? mem[974] : 
                       (N2236)? mem[1038] : 
                       (N2238)? mem[1102] : 
                       (N2240)? mem[1166] : 
                       (N2242)? mem[1230] : 
                       (N2244)? mem[1294] : 
                       (N2246)? mem[1358] : 
                       (N2248)? mem[1422] : 
                       (N2250)? mem[1486] : 
                       (N2252)? mem[1550] : 
                       (N2254)? mem[1614] : 
                       (N2256)? mem[1678] : 
                       (N2258)? mem[1742] : 
                       (N2260)? mem[1806] : 
                       (N2262)? mem[1870] : 
                       (N2264)? mem[1934] : 
                       (N2266)? mem[1998] : 1'b0;
  assign rdata_o[13] = (N2235)? mem[13] : 
                       (N2237)? mem[77] : 
                       (N2239)? mem[141] : 
                       (N2241)? mem[205] : 
                       (N2243)? mem[269] : 
                       (N2245)? mem[333] : 
                       (N2247)? mem[397] : 
                       (N2249)? mem[461] : 
                       (N2251)? mem[525] : 
                       (N2253)? mem[589] : 
                       (N2255)? mem[653] : 
                       (N2257)? mem[717] : 
                       (N2259)? mem[781] : 
                       (N2261)? mem[845] : 
                       (N2263)? mem[909] : 
                       (N2265)? mem[973] : 
                       (N2236)? mem[1037] : 
                       (N2238)? mem[1101] : 
                       (N2240)? mem[1165] : 
                       (N2242)? mem[1229] : 
                       (N2244)? mem[1293] : 
                       (N2246)? mem[1357] : 
                       (N2248)? mem[1421] : 
                       (N2250)? mem[1485] : 
                       (N2252)? mem[1549] : 
                       (N2254)? mem[1613] : 
                       (N2256)? mem[1677] : 
                       (N2258)? mem[1741] : 
                       (N2260)? mem[1805] : 
                       (N2262)? mem[1869] : 
                       (N2264)? mem[1933] : 
                       (N2266)? mem[1997] : 1'b0;
  assign rdata_o[12] = (N2235)? mem[12] : 
                       (N2237)? mem[76] : 
                       (N2239)? mem[140] : 
                       (N2241)? mem[204] : 
                       (N2243)? mem[268] : 
                       (N2245)? mem[332] : 
                       (N2247)? mem[396] : 
                       (N2249)? mem[460] : 
                       (N2251)? mem[524] : 
                       (N2253)? mem[588] : 
                       (N2255)? mem[652] : 
                       (N2257)? mem[716] : 
                       (N2259)? mem[780] : 
                       (N2261)? mem[844] : 
                       (N2263)? mem[908] : 
                       (N2265)? mem[972] : 
                       (N2236)? mem[1036] : 
                       (N2238)? mem[1100] : 
                       (N2240)? mem[1164] : 
                       (N2242)? mem[1228] : 
                       (N2244)? mem[1292] : 
                       (N2246)? mem[1356] : 
                       (N2248)? mem[1420] : 
                       (N2250)? mem[1484] : 
                       (N2252)? mem[1548] : 
                       (N2254)? mem[1612] : 
                       (N2256)? mem[1676] : 
                       (N2258)? mem[1740] : 
                       (N2260)? mem[1804] : 
                       (N2262)? mem[1868] : 
                       (N2264)? mem[1932] : 
                       (N2266)? mem[1996] : 1'b0;
  assign rdata_o[11] = (N2235)? mem[11] : 
                       (N2237)? mem[75] : 
                       (N2239)? mem[139] : 
                       (N2241)? mem[203] : 
                       (N2243)? mem[267] : 
                       (N2245)? mem[331] : 
                       (N2247)? mem[395] : 
                       (N2249)? mem[459] : 
                       (N2251)? mem[523] : 
                       (N2253)? mem[587] : 
                       (N2255)? mem[651] : 
                       (N2257)? mem[715] : 
                       (N2259)? mem[779] : 
                       (N2261)? mem[843] : 
                       (N2263)? mem[907] : 
                       (N2265)? mem[971] : 
                       (N2236)? mem[1035] : 
                       (N2238)? mem[1099] : 
                       (N2240)? mem[1163] : 
                       (N2242)? mem[1227] : 
                       (N2244)? mem[1291] : 
                       (N2246)? mem[1355] : 
                       (N2248)? mem[1419] : 
                       (N2250)? mem[1483] : 
                       (N2252)? mem[1547] : 
                       (N2254)? mem[1611] : 
                       (N2256)? mem[1675] : 
                       (N2258)? mem[1739] : 
                       (N2260)? mem[1803] : 
                       (N2262)? mem[1867] : 
                       (N2264)? mem[1931] : 
                       (N2266)? mem[1995] : 1'b0;
  assign rdata_o[10] = (N2235)? mem[10] : 
                       (N2237)? mem[74] : 
                       (N2239)? mem[138] : 
                       (N2241)? mem[202] : 
                       (N2243)? mem[266] : 
                       (N2245)? mem[330] : 
                       (N2247)? mem[394] : 
                       (N2249)? mem[458] : 
                       (N2251)? mem[522] : 
                       (N2253)? mem[586] : 
                       (N2255)? mem[650] : 
                       (N2257)? mem[714] : 
                       (N2259)? mem[778] : 
                       (N2261)? mem[842] : 
                       (N2263)? mem[906] : 
                       (N2265)? mem[970] : 
                       (N2236)? mem[1034] : 
                       (N2238)? mem[1098] : 
                       (N2240)? mem[1162] : 
                       (N2242)? mem[1226] : 
                       (N2244)? mem[1290] : 
                       (N2246)? mem[1354] : 
                       (N2248)? mem[1418] : 
                       (N2250)? mem[1482] : 
                       (N2252)? mem[1546] : 
                       (N2254)? mem[1610] : 
                       (N2256)? mem[1674] : 
                       (N2258)? mem[1738] : 
                       (N2260)? mem[1802] : 
                       (N2262)? mem[1866] : 
                       (N2264)? mem[1930] : 
                       (N2266)? mem[1994] : 1'b0;
  assign rdata_o[9] = (N2235)? mem[9] : 
                      (N2237)? mem[73] : 
                      (N2239)? mem[137] : 
                      (N2241)? mem[201] : 
                      (N2243)? mem[265] : 
                      (N2245)? mem[329] : 
                      (N2247)? mem[393] : 
                      (N2249)? mem[457] : 
                      (N2251)? mem[521] : 
                      (N2253)? mem[585] : 
                      (N2255)? mem[649] : 
                      (N2257)? mem[713] : 
                      (N2259)? mem[777] : 
                      (N2261)? mem[841] : 
                      (N2263)? mem[905] : 
                      (N2265)? mem[969] : 
                      (N2236)? mem[1033] : 
                      (N2238)? mem[1097] : 
                      (N2240)? mem[1161] : 
                      (N2242)? mem[1225] : 
                      (N2244)? mem[1289] : 
                      (N2246)? mem[1353] : 
                      (N2248)? mem[1417] : 
                      (N2250)? mem[1481] : 
                      (N2252)? mem[1545] : 
                      (N2254)? mem[1609] : 
                      (N2256)? mem[1673] : 
                      (N2258)? mem[1737] : 
                      (N2260)? mem[1801] : 
                      (N2262)? mem[1865] : 
                      (N2264)? mem[1929] : 
                      (N2266)? mem[1993] : 1'b0;
  assign rdata_o[8] = (N2235)? mem[8] : 
                      (N2237)? mem[72] : 
                      (N2239)? mem[136] : 
                      (N2241)? mem[200] : 
                      (N2243)? mem[264] : 
                      (N2245)? mem[328] : 
                      (N2247)? mem[392] : 
                      (N2249)? mem[456] : 
                      (N2251)? mem[520] : 
                      (N2253)? mem[584] : 
                      (N2255)? mem[648] : 
                      (N2257)? mem[712] : 
                      (N2259)? mem[776] : 
                      (N2261)? mem[840] : 
                      (N2263)? mem[904] : 
                      (N2265)? mem[968] : 
                      (N2236)? mem[1032] : 
                      (N2238)? mem[1096] : 
                      (N2240)? mem[1160] : 
                      (N2242)? mem[1224] : 
                      (N2244)? mem[1288] : 
                      (N2246)? mem[1352] : 
                      (N2248)? mem[1416] : 
                      (N2250)? mem[1480] : 
                      (N2252)? mem[1544] : 
                      (N2254)? mem[1608] : 
                      (N2256)? mem[1672] : 
                      (N2258)? mem[1736] : 
                      (N2260)? mem[1800] : 
                      (N2262)? mem[1864] : 
                      (N2264)? mem[1928] : 
                      (N2266)? mem[1992] : 1'b0;
  assign rdata_o[7] = (N2235)? mem[7] : 
                      (N2237)? mem[71] : 
                      (N2239)? mem[135] : 
                      (N2241)? mem[199] : 
                      (N2243)? mem[263] : 
                      (N2245)? mem[327] : 
                      (N2247)? mem[391] : 
                      (N2249)? mem[455] : 
                      (N2251)? mem[519] : 
                      (N2253)? mem[583] : 
                      (N2255)? mem[647] : 
                      (N2257)? mem[711] : 
                      (N2259)? mem[775] : 
                      (N2261)? mem[839] : 
                      (N2263)? mem[903] : 
                      (N2265)? mem[967] : 
                      (N2236)? mem[1031] : 
                      (N2238)? mem[1095] : 
                      (N2240)? mem[1159] : 
                      (N2242)? mem[1223] : 
                      (N2244)? mem[1287] : 
                      (N2246)? mem[1351] : 
                      (N2248)? mem[1415] : 
                      (N2250)? mem[1479] : 
                      (N2252)? mem[1543] : 
                      (N2254)? mem[1607] : 
                      (N2256)? mem[1671] : 
                      (N2258)? mem[1735] : 
                      (N2260)? mem[1799] : 
                      (N2262)? mem[1863] : 
                      (N2264)? mem[1927] : 
                      (N2266)? mem[1991] : 1'b0;
  assign rdata_o[6] = (N2235)? mem[6] : 
                      (N2237)? mem[70] : 
                      (N2239)? mem[134] : 
                      (N2241)? mem[198] : 
                      (N2243)? mem[262] : 
                      (N2245)? mem[326] : 
                      (N2247)? mem[390] : 
                      (N2249)? mem[454] : 
                      (N2251)? mem[518] : 
                      (N2253)? mem[582] : 
                      (N2255)? mem[646] : 
                      (N2257)? mem[710] : 
                      (N2259)? mem[774] : 
                      (N2261)? mem[838] : 
                      (N2263)? mem[902] : 
                      (N2265)? mem[966] : 
                      (N2236)? mem[1030] : 
                      (N2238)? mem[1094] : 
                      (N2240)? mem[1158] : 
                      (N2242)? mem[1222] : 
                      (N2244)? mem[1286] : 
                      (N2246)? mem[1350] : 
                      (N2248)? mem[1414] : 
                      (N2250)? mem[1478] : 
                      (N2252)? mem[1542] : 
                      (N2254)? mem[1606] : 
                      (N2256)? mem[1670] : 
                      (N2258)? mem[1734] : 
                      (N2260)? mem[1798] : 
                      (N2262)? mem[1862] : 
                      (N2264)? mem[1926] : 
                      (N2266)? mem[1990] : 1'b0;
  assign rdata_o[5] = (N2235)? mem[5] : 
                      (N2237)? mem[69] : 
                      (N2239)? mem[133] : 
                      (N2241)? mem[197] : 
                      (N2243)? mem[261] : 
                      (N2245)? mem[325] : 
                      (N2247)? mem[389] : 
                      (N2249)? mem[453] : 
                      (N2251)? mem[517] : 
                      (N2253)? mem[581] : 
                      (N2255)? mem[645] : 
                      (N2257)? mem[709] : 
                      (N2259)? mem[773] : 
                      (N2261)? mem[837] : 
                      (N2263)? mem[901] : 
                      (N2265)? mem[965] : 
                      (N2236)? mem[1029] : 
                      (N2238)? mem[1093] : 
                      (N2240)? mem[1157] : 
                      (N2242)? mem[1221] : 
                      (N2244)? mem[1285] : 
                      (N2246)? mem[1349] : 
                      (N2248)? mem[1413] : 
                      (N2250)? mem[1477] : 
                      (N2252)? mem[1541] : 
                      (N2254)? mem[1605] : 
                      (N2256)? mem[1669] : 
                      (N2258)? mem[1733] : 
                      (N2260)? mem[1797] : 
                      (N2262)? mem[1861] : 
                      (N2264)? mem[1925] : 
                      (N2266)? mem[1989] : 1'b0;
  assign rdata_o[4] = (N2235)? mem[4] : 
                      (N2237)? mem[68] : 
                      (N2239)? mem[132] : 
                      (N2241)? mem[196] : 
                      (N2243)? mem[260] : 
                      (N2245)? mem[324] : 
                      (N2247)? mem[388] : 
                      (N2249)? mem[452] : 
                      (N2251)? mem[516] : 
                      (N2253)? mem[580] : 
                      (N2255)? mem[644] : 
                      (N2257)? mem[708] : 
                      (N2259)? mem[772] : 
                      (N2261)? mem[836] : 
                      (N2263)? mem[900] : 
                      (N2265)? mem[964] : 
                      (N2236)? mem[1028] : 
                      (N2238)? mem[1092] : 
                      (N2240)? mem[1156] : 
                      (N2242)? mem[1220] : 
                      (N2244)? mem[1284] : 
                      (N2246)? mem[1348] : 
                      (N2248)? mem[1412] : 
                      (N2250)? mem[1476] : 
                      (N2252)? mem[1540] : 
                      (N2254)? mem[1604] : 
                      (N2256)? mem[1668] : 
                      (N2258)? mem[1732] : 
                      (N2260)? mem[1796] : 
                      (N2262)? mem[1860] : 
                      (N2264)? mem[1924] : 
                      (N2266)? mem[1988] : 1'b0;
  assign rdata_o[3] = (N2235)? mem[3] : 
                      (N2237)? mem[67] : 
                      (N2239)? mem[131] : 
                      (N2241)? mem[195] : 
                      (N2243)? mem[259] : 
                      (N2245)? mem[323] : 
                      (N2247)? mem[387] : 
                      (N2249)? mem[451] : 
                      (N2251)? mem[515] : 
                      (N2253)? mem[579] : 
                      (N2255)? mem[643] : 
                      (N2257)? mem[707] : 
                      (N2259)? mem[771] : 
                      (N2261)? mem[835] : 
                      (N2263)? mem[899] : 
                      (N2265)? mem[963] : 
                      (N2236)? mem[1027] : 
                      (N2238)? mem[1091] : 
                      (N2240)? mem[1155] : 
                      (N2242)? mem[1219] : 
                      (N2244)? mem[1283] : 
                      (N2246)? mem[1347] : 
                      (N2248)? mem[1411] : 
                      (N2250)? mem[1475] : 
                      (N2252)? mem[1539] : 
                      (N2254)? mem[1603] : 
                      (N2256)? mem[1667] : 
                      (N2258)? mem[1731] : 
                      (N2260)? mem[1795] : 
                      (N2262)? mem[1859] : 
                      (N2264)? mem[1923] : 
                      (N2266)? mem[1987] : 1'b0;
  assign rdata_o[2] = (N2235)? mem[2] : 
                      (N2237)? mem[66] : 
                      (N2239)? mem[130] : 
                      (N2241)? mem[194] : 
                      (N2243)? mem[258] : 
                      (N2245)? mem[322] : 
                      (N2247)? mem[386] : 
                      (N2249)? mem[450] : 
                      (N2251)? mem[514] : 
                      (N2253)? mem[578] : 
                      (N2255)? mem[642] : 
                      (N2257)? mem[706] : 
                      (N2259)? mem[770] : 
                      (N2261)? mem[834] : 
                      (N2263)? mem[898] : 
                      (N2265)? mem[962] : 
                      (N2236)? mem[1026] : 
                      (N2238)? mem[1090] : 
                      (N2240)? mem[1154] : 
                      (N2242)? mem[1218] : 
                      (N2244)? mem[1282] : 
                      (N2246)? mem[1346] : 
                      (N2248)? mem[1410] : 
                      (N2250)? mem[1474] : 
                      (N2252)? mem[1538] : 
                      (N2254)? mem[1602] : 
                      (N2256)? mem[1666] : 
                      (N2258)? mem[1730] : 
                      (N2260)? mem[1794] : 
                      (N2262)? mem[1858] : 
                      (N2264)? mem[1922] : 
                      (N2266)? mem[1986] : 1'b0;
  assign rdata_o[1] = (N2235)? mem[1] : 
                      (N2237)? mem[65] : 
                      (N2239)? mem[129] : 
                      (N2241)? mem[193] : 
                      (N2243)? mem[257] : 
                      (N2245)? mem[321] : 
                      (N2247)? mem[385] : 
                      (N2249)? mem[449] : 
                      (N2251)? mem[513] : 
                      (N2253)? mem[577] : 
                      (N2255)? mem[641] : 
                      (N2257)? mem[705] : 
                      (N2259)? mem[769] : 
                      (N2261)? mem[833] : 
                      (N2263)? mem[897] : 
                      (N2265)? mem[961] : 
                      (N2236)? mem[1025] : 
                      (N2238)? mem[1089] : 
                      (N2240)? mem[1153] : 
                      (N2242)? mem[1217] : 
                      (N2244)? mem[1281] : 
                      (N2246)? mem[1345] : 
                      (N2248)? mem[1409] : 
                      (N2250)? mem[1473] : 
                      (N2252)? mem[1537] : 
                      (N2254)? mem[1601] : 
                      (N2256)? mem[1665] : 
                      (N2258)? mem[1729] : 
                      (N2260)? mem[1793] : 
                      (N2262)? mem[1857] : 
                      (N2264)? mem[1921] : 
                      (N2266)? mem[1985] : 1'b0;
  assign rdata_o[0] = (N2235)? mem[0] : 
                      (N2237)? mem[64] : 
                      (N2239)? mem[128] : 
                      (N2241)? mem[192] : 
                      (N2243)? mem[256] : 
                      (N2245)? mem[320] : 
                      (N2247)? mem[384] : 
                      (N2249)? mem[448] : 
                      (N2251)? mem[512] : 
                      (N2253)? mem[576] : 
                      (N2255)? mem[640] : 
                      (N2257)? mem[704] : 
                      (N2259)? mem[768] : 
                      (N2261)? mem[832] : 
                      (N2263)? mem[896] : 
                      (N2265)? mem[960] : 
                      (N2236)? mem[1024] : 
                      (N2238)? mem[1088] : 
                      (N2240)? mem[1152] : 
                      (N2242)? mem[1216] : 
                      (N2244)? mem[1280] : 
                      (N2246)? mem[1344] : 
                      (N2248)? mem[1408] : 
                      (N2250)? mem[1472] : 
                      (N2252)? mem[1536] : 
                      (N2254)? mem[1600] : 
                      (N2256)? mem[1664] : 
                      (N2258)? mem[1728] : 
                      (N2260)? mem[1792] : 
                      (N2262)? mem[1856] : 
                      (N2264)? mem[1920] : 
                      (N2266)? mem[1984] : 1'b0;
  assign rdata_o[127] = (N2300)? mem[63] : 
                        (N2302)? mem[127] : 
                        (N2304)? mem[191] : 
                        (N2306)? mem[255] : 
                        (N2308)? mem[319] : 
                        (N2310)? mem[383] : 
                        (N2312)? mem[447] : 
                        (N2314)? mem[511] : 
                        (N2316)? mem[575] : 
                        (N2318)? mem[639] : 
                        (N2320)? mem[703] : 
                        (N2322)? mem[767] : 
                        (N2324)? mem[831] : 
                        (N2326)? mem[895] : 
                        (N2328)? mem[959] : 
                        (N2330)? mem[1023] : 
                        (N2301)? mem[1087] : 
                        (N2303)? mem[1151] : 
                        (N2305)? mem[1215] : 
                        (N2307)? mem[1279] : 
                        (N2309)? mem[1343] : 
                        (N2311)? mem[1407] : 
                        (N2313)? mem[1471] : 
                        (N2315)? mem[1535] : 
                        (N2317)? mem[1599] : 
                        (N2319)? mem[1663] : 
                        (N2321)? mem[1727] : 
                        (N2323)? mem[1791] : 
                        (N2325)? mem[1855] : 
                        (N2327)? mem[1919] : 
                        (N2329)? mem[1983] : 
                        (N2331)? mem[2047] : 1'b0;
  assign rdata_o[126] = (N2300)? mem[62] : 
                        (N2302)? mem[126] : 
                        (N2304)? mem[190] : 
                        (N2306)? mem[254] : 
                        (N2308)? mem[318] : 
                        (N2310)? mem[382] : 
                        (N2312)? mem[446] : 
                        (N2314)? mem[510] : 
                        (N2316)? mem[574] : 
                        (N2318)? mem[638] : 
                        (N2320)? mem[702] : 
                        (N2322)? mem[766] : 
                        (N2324)? mem[830] : 
                        (N2326)? mem[894] : 
                        (N2328)? mem[958] : 
                        (N2330)? mem[1022] : 
                        (N2301)? mem[1086] : 
                        (N2303)? mem[1150] : 
                        (N2305)? mem[1214] : 
                        (N2307)? mem[1278] : 
                        (N2309)? mem[1342] : 
                        (N2311)? mem[1406] : 
                        (N2313)? mem[1470] : 
                        (N2315)? mem[1534] : 
                        (N2317)? mem[1598] : 
                        (N2319)? mem[1662] : 
                        (N2321)? mem[1726] : 
                        (N2323)? mem[1790] : 
                        (N2325)? mem[1854] : 
                        (N2327)? mem[1918] : 
                        (N2329)? mem[1982] : 
                        (N2331)? mem[2046] : 1'b0;
  assign rdata_o[125] = (N2300)? mem[61] : 
                        (N2302)? mem[125] : 
                        (N2304)? mem[189] : 
                        (N2306)? mem[253] : 
                        (N2308)? mem[317] : 
                        (N2310)? mem[381] : 
                        (N2312)? mem[445] : 
                        (N2314)? mem[509] : 
                        (N2316)? mem[573] : 
                        (N2318)? mem[637] : 
                        (N2320)? mem[701] : 
                        (N2322)? mem[765] : 
                        (N2324)? mem[829] : 
                        (N2326)? mem[893] : 
                        (N2328)? mem[957] : 
                        (N2330)? mem[1021] : 
                        (N2301)? mem[1085] : 
                        (N2303)? mem[1149] : 
                        (N2305)? mem[1213] : 
                        (N2307)? mem[1277] : 
                        (N2309)? mem[1341] : 
                        (N2311)? mem[1405] : 
                        (N2313)? mem[1469] : 
                        (N2315)? mem[1533] : 
                        (N2317)? mem[1597] : 
                        (N2319)? mem[1661] : 
                        (N2321)? mem[1725] : 
                        (N2323)? mem[1789] : 
                        (N2325)? mem[1853] : 
                        (N2327)? mem[1917] : 
                        (N2329)? mem[1981] : 
                        (N2331)? mem[2045] : 1'b0;
  assign rdata_o[124] = (N2300)? mem[60] : 
                        (N2302)? mem[124] : 
                        (N2304)? mem[188] : 
                        (N2306)? mem[252] : 
                        (N2308)? mem[316] : 
                        (N2310)? mem[380] : 
                        (N2312)? mem[444] : 
                        (N2314)? mem[508] : 
                        (N2316)? mem[572] : 
                        (N2318)? mem[636] : 
                        (N2320)? mem[700] : 
                        (N2322)? mem[764] : 
                        (N2324)? mem[828] : 
                        (N2326)? mem[892] : 
                        (N2328)? mem[956] : 
                        (N2330)? mem[1020] : 
                        (N2301)? mem[1084] : 
                        (N2303)? mem[1148] : 
                        (N2305)? mem[1212] : 
                        (N2307)? mem[1276] : 
                        (N2309)? mem[1340] : 
                        (N2311)? mem[1404] : 
                        (N2313)? mem[1468] : 
                        (N2315)? mem[1532] : 
                        (N2317)? mem[1596] : 
                        (N2319)? mem[1660] : 
                        (N2321)? mem[1724] : 
                        (N2323)? mem[1788] : 
                        (N2325)? mem[1852] : 
                        (N2327)? mem[1916] : 
                        (N2329)? mem[1980] : 
                        (N2331)? mem[2044] : 1'b0;
  assign rdata_o[123] = (N2300)? mem[59] : 
                        (N2302)? mem[123] : 
                        (N2304)? mem[187] : 
                        (N2306)? mem[251] : 
                        (N2308)? mem[315] : 
                        (N2310)? mem[379] : 
                        (N2312)? mem[443] : 
                        (N2314)? mem[507] : 
                        (N2316)? mem[571] : 
                        (N2318)? mem[635] : 
                        (N2320)? mem[699] : 
                        (N2322)? mem[763] : 
                        (N2324)? mem[827] : 
                        (N2326)? mem[891] : 
                        (N2328)? mem[955] : 
                        (N2330)? mem[1019] : 
                        (N2301)? mem[1083] : 
                        (N2303)? mem[1147] : 
                        (N2305)? mem[1211] : 
                        (N2307)? mem[1275] : 
                        (N2309)? mem[1339] : 
                        (N2311)? mem[1403] : 
                        (N2313)? mem[1467] : 
                        (N2315)? mem[1531] : 
                        (N2317)? mem[1595] : 
                        (N2319)? mem[1659] : 
                        (N2321)? mem[1723] : 
                        (N2323)? mem[1787] : 
                        (N2325)? mem[1851] : 
                        (N2327)? mem[1915] : 
                        (N2329)? mem[1979] : 
                        (N2331)? mem[2043] : 1'b0;
  assign rdata_o[122] = (N2300)? mem[58] : 
                        (N2302)? mem[122] : 
                        (N2304)? mem[186] : 
                        (N2306)? mem[250] : 
                        (N2308)? mem[314] : 
                        (N2310)? mem[378] : 
                        (N2312)? mem[442] : 
                        (N2314)? mem[506] : 
                        (N2316)? mem[570] : 
                        (N2318)? mem[634] : 
                        (N2320)? mem[698] : 
                        (N2322)? mem[762] : 
                        (N2324)? mem[826] : 
                        (N2326)? mem[890] : 
                        (N2328)? mem[954] : 
                        (N2330)? mem[1018] : 
                        (N2301)? mem[1082] : 
                        (N2303)? mem[1146] : 
                        (N2305)? mem[1210] : 
                        (N2307)? mem[1274] : 
                        (N2309)? mem[1338] : 
                        (N2311)? mem[1402] : 
                        (N2313)? mem[1466] : 
                        (N2315)? mem[1530] : 
                        (N2317)? mem[1594] : 
                        (N2319)? mem[1658] : 
                        (N2321)? mem[1722] : 
                        (N2323)? mem[1786] : 
                        (N2325)? mem[1850] : 
                        (N2327)? mem[1914] : 
                        (N2329)? mem[1978] : 
                        (N2331)? mem[2042] : 1'b0;
  assign rdata_o[121] = (N2300)? mem[57] : 
                        (N2302)? mem[121] : 
                        (N2304)? mem[185] : 
                        (N2306)? mem[249] : 
                        (N2308)? mem[313] : 
                        (N2310)? mem[377] : 
                        (N2312)? mem[441] : 
                        (N2314)? mem[505] : 
                        (N2316)? mem[569] : 
                        (N2318)? mem[633] : 
                        (N2320)? mem[697] : 
                        (N2322)? mem[761] : 
                        (N2324)? mem[825] : 
                        (N2326)? mem[889] : 
                        (N2328)? mem[953] : 
                        (N2330)? mem[1017] : 
                        (N2301)? mem[1081] : 
                        (N2303)? mem[1145] : 
                        (N2305)? mem[1209] : 
                        (N2307)? mem[1273] : 
                        (N2309)? mem[1337] : 
                        (N2311)? mem[1401] : 
                        (N2313)? mem[1465] : 
                        (N2315)? mem[1529] : 
                        (N2317)? mem[1593] : 
                        (N2319)? mem[1657] : 
                        (N2321)? mem[1721] : 
                        (N2323)? mem[1785] : 
                        (N2325)? mem[1849] : 
                        (N2327)? mem[1913] : 
                        (N2329)? mem[1977] : 
                        (N2331)? mem[2041] : 1'b0;
  assign rdata_o[120] = (N2300)? mem[56] : 
                        (N2302)? mem[120] : 
                        (N2304)? mem[184] : 
                        (N2306)? mem[248] : 
                        (N2308)? mem[312] : 
                        (N2310)? mem[376] : 
                        (N2312)? mem[440] : 
                        (N2314)? mem[504] : 
                        (N2316)? mem[568] : 
                        (N2318)? mem[632] : 
                        (N2320)? mem[696] : 
                        (N2322)? mem[760] : 
                        (N2324)? mem[824] : 
                        (N2326)? mem[888] : 
                        (N2328)? mem[952] : 
                        (N2330)? mem[1016] : 
                        (N2301)? mem[1080] : 
                        (N2303)? mem[1144] : 
                        (N2305)? mem[1208] : 
                        (N2307)? mem[1272] : 
                        (N2309)? mem[1336] : 
                        (N2311)? mem[1400] : 
                        (N2313)? mem[1464] : 
                        (N2315)? mem[1528] : 
                        (N2317)? mem[1592] : 
                        (N2319)? mem[1656] : 
                        (N2321)? mem[1720] : 
                        (N2323)? mem[1784] : 
                        (N2325)? mem[1848] : 
                        (N2327)? mem[1912] : 
                        (N2329)? mem[1976] : 
                        (N2331)? mem[2040] : 1'b0;
  assign rdata_o[119] = (N2300)? mem[55] : 
                        (N2302)? mem[119] : 
                        (N2304)? mem[183] : 
                        (N2306)? mem[247] : 
                        (N2308)? mem[311] : 
                        (N2310)? mem[375] : 
                        (N2312)? mem[439] : 
                        (N2314)? mem[503] : 
                        (N2316)? mem[567] : 
                        (N2318)? mem[631] : 
                        (N2320)? mem[695] : 
                        (N2322)? mem[759] : 
                        (N2324)? mem[823] : 
                        (N2326)? mem[887] : 
                        (N2328)? mem[951] : 
                        (N2330)? mem[1015] : 
                        (N2301)? mem[1079] : 
                        (N2303)? mem[1143] : 
                        (N2305)? mem[1207] : 
                        (N2307)? mem[1271] : 
                        (N2309)? mem[1335] : 
                        (N2311)? mem[1399] : 
                        (N2313)? mem[1463] : 
                        (N2315)? mem[1527] : 
                        (N2317)? mem[1591] : 
                        (N2319)? mem[1655] : 
                        (N2321)? mem[1719] : 
                        (N2323)? mem[1783] : 
                        (N2325)? mem[1847] : 
                        (N2327)? mem[1911] : 
                        (N2329)? mem[1975] : 
                        (N2331)? mem[2039] : 1'b0;
  assign rdata_o[118] = (N2300)? mem[54] : 
                        (N2302)? mem[118] : 
                        (N2304)? mem[182] : 
                        (N2306)? mem[246] : 
                        (N2308)? mem[310] : 
                        (N2310)? mem[374] : 
                        (N2312)? mem[438] : 
                        (N2314)? mem[502] : 
                        (N2316)? mem[566] : 
                        (N2318)? mem[630] : 
                        (N2320)? mem[694] : 
                        (N2322)? mem[758] : 
                        (N2324)? mem[822] : 
                        (N2326)? mem[886] : 
                        (N2328)? mem[950] : 
                        (N2330)? mem[1014] : 
                        (N2301)? mem[1078] : 
                        (N2303)? mem[1142] : 
                        (N2305)? mem[1206] : 
                        (N2307)? mem[1270] : 
                        (N2309)? mem[1334] : 
                        (N2311)? mem[1398] : 
                        (N2313)? mem[1462] : 
                        (N2315)? mem[1526] : 
                        (N2317)? mem[1590] : 
                        (N2319)? mem[1654] : 
                        (N2321)? mem[1718] : 
                        (N2323)? mem[1782] : 
                        (N2325)? mem[1846] : 
                        (N2327)? mem[1910] : 
                        (N2329)? mem[1974] : 
                        (N2331)? mem[2038] : 1'b0;
  assign rdata_o[117] = (N2300)? mem[53] : 
                        (N2302)? mem[117] : 
                        (N2304)? mem[181] : 
                        (N2306)? mem[245] : 
                        (N2308)? mem[309] : 
                        (N2310)? mem[373] : 
                        (N2312)? mem[437] : 
                        (N2314)? mem[501] : 
                        (N2316)? mem[565] : 
                        (N2318)? mem[629] : 
                        (N2320)? mem[693] : 
                        (N2322)? mem[757] : 
                        (N2324)? mem[821] : 
                        (N2326)? mem[885] : 
                        (N2328)? mem[949] : 
                        (N2330)? mem[1013] : 
                        (N2301)? mem[1077] : 
                        (N2303)? mem[1141] : 
                        (N2305)? mem[1205] : 
                        (N2307)? mem[1269] : 
                        (N2309)? mem[1333] : 
                        (N2311)? mem[1397] : 
                        (N2313)? mem[1461] : 
                        (N2315)? mem[1525] : 
                        (N2317)? mem[1589] : 
                        (N2319)? mem[1653] : 
                        (N2321)? mem[1717] : 
                        (N2323)? mem[1781] : 
                        (N2325)? mem[1845] : 
                        (N2327)? mem[1909] : 
                        (N2329)? mem[1973] : 
                        (N2331)? mem[2037] : 1'b0;
  assign rdata_o[116] = (N2300)? mem[52] : 
                        (N2302)? mem[116] : 
                        (N2304)? mem[180] : 
                        (N2306)? mem[244] : 
                        (N2308)? mem[308] : 
                        (N2310)? mem[372] : 
                        (N2312)? mem[436] : 
                        (N2314)? mem[500] : 
                        (N2316)? mem[564] : 
                        (N2318)? mem[628] : 
                        (N2320)? mem[692] : 
                        (N2322)? mem[756] : 
                        (N2324)? mem[820] : 
                        (N2326)? mem[884] : 
                        (N2328)? mem[948] : 
                        (N2330)? mem[1012] : 
                        (N2301)? mem[1076] : 
                        (N2303)? mem[1140] : 
                        (N2305)? mem[1204] : 
                        (N2307)? mem[1268] : 
                        (N2309)? mem[1332] : 
                        (N2311)? mem[1396] : 
                        (N2313)? mem[1460] : 
                        (N2315)? mem[1524] : 
                        (N2317)? mem[1588] : 
                        (N2319)? mem[1652] : 
                        (N2321)? mem[1716] : 
                        (N2323)? mem[1780] : 
                        (N2325)? mem[1844] : 
                        (N2327)? mem[1908] : 
                        (N2329)? mem[1972] : 
                        (N2331)? mem[2036] : 1'b0;
  assign rdata_o[115] = (N2300)? mem[51] : 
                        (N2302)? mem[115] : 
                        (N2304)? mem[179] : 
                        (N2306)? mem[243] : 
                        (N2308)? mem[307] : 
                        (N2310)? mem[371] : 
                        (N2312)? mem[435] : 
                        (N2314)? mem[499] : 
                        (N2316)? mem[563] : 
                        (N2318)? mem[627] : 
                        (N2320)? mem[691] : 
                        (N2322)? mem[755] : 
                        (N2324)? mem[819] : 
                        (N2326)? mem[883] : 
                        (N2328)? mem[947] : 
                        (N2330)? mem[1011] : 
                        (N2301)? mem[1075] : 
                        (N2303)? mem[1139] : 
                        (N2305)? mem[1203] : 
                        (N2307)? mem[1267] : 
                        (N2309)? mem[1331] : 
                        (N2311)? mem[1395] : 
                        (N2313)? mem[1459] : 
                        (N2315)? mem[1523] : 
                        (N2317)? mem[1587] : 
                        (N2319)? mem[1651] : 
                        (N2321)? mem[1715] : 
                        (N2323)? mem[1779] : 
                        (N2325)? mem[1843] : 
                        (N2327)? mem[1907] : 
                        (N2329)? mem[1971] : 
                        (N2331)? mem[2035] : 1'b0;
  assign rdata_o[114] = (N2300)? mem[50] : 
                        (N2302)? mem[114] : 
                        (N2304)? mem[178] : 
                        (N2306)? mem[242] : 
                        (N2308)? mem[306] : 
                        (N2310)? mem[370] : 
                        (N2312)? mem[434] : 
                        (N2314)? mem[498] : 
                        (N2316)? mem[562] : 
                        (N2318)? mem[626] : 
                        (N2320)? mem[690] : 
                        (N2322)? mem[754] : 
                        (N2324)? mem[818] : 
                        (N2326)? mem[882] : 
                        (N2328)? mem[946] : 
                        (N2330)? mem[1010] : 
                        (N2301)? mem[1074] : 
                        (N2303)? mem[1138] : 
                        (N2305)? mem[1202] : 
                        (N2307)? mem[1266] : 
                        (N2309)? mem[1330] : 
                        (N2311)? mem[1394] : 
                        (N2313)? mem[1458] : 
                        (N2315)? mem[1522] : 
                        (N2317)? mem[1586] : 
                        (N2319)? mem[1650] : 
                        (N2321)? mem[1714] : 
                        (N2323)? mem[1778] : 
                        (N2325)? mem[1842] : 
                        (N2327)? mem[1906] : 
                        (N2329)? mem[1970] : 
                        (N2331)? mem[2034] : 1'b0;
  assign rdata_o[113] = (N2300)? mem[49] : 
                        (N2302)? mem[113] : 
                        (N2304)? mem[177] : 
                        (N2306)? mem[241] : 
                        (N2308)? mem[305] : 
                        (N2310)? mem[369] : 
                        (N2312)? mem[433] : 
                        (N2314)? mem[497] : 
                        (N2316)? mem[561] : 
                        (N2318)? mem[625] : 
                        (N2320)? mem[689] : 
                        (N2322)? mem[753] : 
                        (N2324)? mem[817] : 
                        (N2326)? mem[881] : 
                        (N2328)? mem[945] : 
                        (N2330)? mem[1009] : 
                        (N2301)? mem[1073] : 
                        (N2303)? mem[1137] : 
                        (N2305)? mem[1201] : 
                        (N2307)? mem[1265] : 
                        (N2309)? mem[1329] : 
                        (N2311)? mem[1393] : 
                        (N2313)? mem[1457] : 
                        (N2315)? mem[1521] : 
                        (N2317)? mem[1585] : 
                        (N2319)? mem[1649] : 
                        (N2321)? mem[1713] : 
                        (N2323)? mem[1777] : 
                        (N2325)? mem[1841] : 
                        (N2327)? mem[1905] : 
                        (N2329)? mem[1969] : 
                        (N2331)? mem[2033] : 1'b0;
  assign rdata_o[112] = (N2300)? mem[48] : 
                        (N2302)? mem[112] : 
                        (N2304)? mem[176] : 
                        (N2306)? mem[240] : 
                        (N2308)? mem[304] : 
                        (N2310)? mem[368] : 
                        (N2312)? mem[432] : 
                        (N2314)? mem[496] : 
                        (N2316)? mem[560] : 
                        (N2318)? mem[624] : 
                        (N2320)? mem[688] : 
                        (N2322)? mem[752] : 
                        (N2324)? mem[816] : 
                        (N2326)? mem[880] : 
                        (N2328)? mem[944] : 
                        (N2330)? mem[1008] : 
                        (N2301)? mem[1072] : 
                        (N2303)? mem[1136] : 
                        (N2305)? mem[1200] : 
                        (N2307)? mem[1264] : 
                        (N2309)? mem[1328] : 
                        (N2311)? mem[1392] : 
                        (N2313)? mem[1456] : 
                        (N2315)? mem[1520] : 
                        (N2317)? mem[1584] : 
                        (N2319)? mem[1648] : 
                        (N2321)? mem[1712] : 
                        (N2323)? mem[1776] : 
                        (N2325)? mem[1840] : 
                        (N2327)? mem[1904] : 
                        (N2329)? mem[1968] : 
                        (N2331)? mem[2032] : 1'b0;
  assign rdata_o[111] = (N2300)? mem[47] : 
                        (N2302)? mem[111] : 
                        (N2304)? mem[175] : 
                        (N2306)? mem[239] : 
                        (N2308)? mem[303] : 
                        (N2310)? mem[367] : 
                        (N2312)? mem[431] : 
                        (N2314)? mem[495] : 
                        (N2316)? mem[559] : 
                        (N2318)? mem[623] : 
                        (N2320)? mem[687] : 
                        (N2322)? mem[751] : 
                        (N2324)? mem[815] : 
                        (N2326)? mem[879] : 
                        (N2328)? mem[943] : 
                        (N2330)? mem[1007] : 
                        (N2301)? mem[1071] : 
                        (N2303)? mem[1135] : 
                        (N2305)? mem[1199] : 
                        (N2307)? mem[1263] : 
                        (N2309)? mem[1327] : 
                        (N2311)? mem[1391] : 
                        (N2313)? mem[1455] : 
                        (N2315)? mem[1519] : 
                        (N2317)? mem[1583] : 
                        (N2319)? mem[1647] : 
                        (N2321)? mem[1711] : 
                        (N2323)? mem[1775] : 
                        (N2325)? mem[1839] : 
                        (N2327)? mem[1903] : 
                        (N2329)? mem[1967] : 
                        (N2331)? mem[2031] : 1'b0;
  assign rdata_o[110] = (N2300)? mem[46] : 
                        (N2302)? mem[110] : 
                        (N2304)? mem[174] : 
                        (N2306)? mem[238] : 
                        (N2308)? mem[302] : 
                        (N2310)? mem[366] : 
                        (N2312)? mem[430] : 
                        (N2314)? mem[494] : 
                        (N2316)? mem[558] : 
                        (N2318)? mem[622] : 
                        (N2320)? mem[686] : 
                        (N2322)? mem[750] : 
                        (N2324)? mem[814] : 
                        (N2326)? mem[878] : 
                        (N2328)? mem[942] : 
                        (N2330)? mem[1006] : 
                        (N2301)? mem[1070] : 
                        (N2303)? mem[1134] : 
                        (N2305)? mem[1198] : 
                        (N2307)? mem[1262] : 
                        (N2309)? mem[1326] : 
                        (N2311)? mem[1390] : 
                        (N2313)? mem[1454] : 
                        (N2315)? mem[1518] : 
                        (N2317)? mem[1582] : 
                        (N2319)? mem[1646] : 
                        (N2321)? mem[1710] : 
                        (N2323)? mem[1774] : 
                        (N2325)? mem[1838] : 
                        (N2327)? mem[1902] : 
                        (N2329)? mem[1966] : 
                        (N2331)? mem[2030] : 1'b0;
  assign rdata_o[109] = (N2300)? mem[45] : 
                        (N2302)? mem[109] : 
                        (N2304)? mem[173] : 
                        (N2306)? mem[237] : 
                        (N2308)? mem[301] : 
                        (N2310)? mem[365] : 
                        (N2312)? mem[429] : 
                        (N2314)? mem[493] : 
                        (N2316)? mem[557] : 
                        (N2318)? mem[621] : 
                        (N2320)? mem[685] : 
                        (N2322)? mem[749] : 
                        (N2324)? mem[813] : 
                        (N2326)? mem[877] : 
                        (N2328)? mem[941] : 
                        (N2330)? mem[1005] : 
                        (N2301)? mem[1069] : 
                        (N2303)? mem[1133] : 
                        (N2305)? mem[1197] : 
                        (N2307)? mem[1261] : 
                        (N2309)? mem[1325] : 
                        (N2311)? mem[1389] : 
                        (N2313)? mem[1453] : 
                        (N2315)? mem[1517] : 
                        (N2317)? mem[1581] : 
                        (N2319)? mem[1645] : 
                        (N2321)? mem[1709] : 
                        (N2323)? mem[1773] : 
                        (N2325)? mem[1837] : 
                        (N2327)? mem[1901] : 
                        (N2329)? mem[1965] : 
                        (N2331)? mem[2029] : 1'b0;
  assign rdata_o[108] = (N2300)? mem[44] : 
                        (N2302)? mem[108] : 
                        (N2304)? mem[172] : 
                        (N2306)? mem[236] : 
                        (N2308)? mem[300] : 
                        (N2310)? mem[364] : 
                        (N2312)? mem[428] : 
                        (N2314)? mem[492] : 
                        (N2316)? mem[556] : 
                        (N2318)? mem[620] : 
                        (N2320)? mem[684] : 
                        (N2322)? mem[748] : 
                        (N2324)? mem[812] : 
                        (N2326)? mem[876] : 
                        (N2328)? mem[940] : 
                        (N2330)? mem[1004] : 
                        (N2301)? mem[1068] : 
                        (N2303)? mem[1132] : 
                        (N2305)? mem[1196] : 
                        (N2307)? mem[1260] : 
                        (N2309)? mem[1324] : 
                        (N2311)? mem[1388] : 
                        (N2313)? mem[1452] : 
                        (N2315)? mem[1516] : 
                        (N2317)? mem[1580] : 
                        (N2319)? mem[1644] : 
                        (N2321)? mem[1708] : 
                        (N2323)? mem[1772] : 
                        (N2325)? mem[1836] : 
                        (N2327)? mem[1900] : 
                        (N2329)? mem[1964] : 
                        (N2331)? mem[2028] : 1'b0;
  assign rdata_o[107] = (N2300)? mem[43] : 
                        (N2302)? mem[107] : 
                        (N2304)? mem[171] : 
                        (N2306)? mem[235] : 
                        (N2308)? mem[299] : 
                        (N2310)? mem[363] : 
                        (N2312)? mem[427] : 
                        (N2314)? mem[491] : 
                        (N2316)? mem[555] : 
                        (N2318)? mem[619] : 
                        (N2320)? mem[683] : 
                        (N2322)? mem[747] : 
                        (N2324)? mem[811] : 
                        (N2326)? mem[875] : 
                        (N2328)? mem[939] : 
                        (N2330)? mem[1003] : 
                        (N2301)? mem[1067] : 
                        (N2303)? mem[1131] : 
                        (N2305)? mem[1195] : 
                        (N2307)? mem[1259] : 
                        (N2309)? mem[1323] : 
                        (N2311)? mem[1387] : 
                        (N2313)? mem[1451] : 
                        (N2315)? mem[1515] : 
                        (N2317)? mem[1579] : 
                        (N2319)? mem[1643] : 
                        (N2321)? mem[1707] : 
                        (N2323)? mem[1771] : 
                        (N2325)? mem[1835] : 
                        (N2327)? mem[1899] : 
                        (N2329)? mem[1963] : 
                        (N2331)? mem[2027] : 1'b0;
  assign rdata_o[106] = (N2300)? mem[42] : 
                        (N2302)? mem[106] : 
                        (N2304)? mem[170] : 
                        (N2306)? mem[234] : 
                        (N2308)? mem[298] : 
                        (N2310)? mem[362] : 
                        (N2312)? mem[426] : 
                        (N2314)? mem[490] : 
                        (N2316)? mem[554] : 
                        (N2318)? mem[618] : 
                        (N2320)? mem[682] : 
                        (N2322)? mem[746] : 
                        (N2324)? mem[810] : 
                        (N2326)? mem[874] : 
                        (N2328)? mem[938] : 
                        (N2330)? mem[1002] : 
                        (N2301)? mem[1066] : 
                        (N2303)? mem[1130] : 
                        (N2305)? mem[1194] : 
                        (N2307)? mem[1258] : 
                        (N2309)? mem[1322] : 
                        (N2311)? mem[1386] : 
                        (N2313)? mem[1450] : 
                        (N2315)? mem[1514] : 
                        (N2317)? mem[1578] : 
                        (N2319)? mem[1642] : 
                        (N2321)? mem[1706] : 
                        (N2323)? mem[1770] : 
                        (N2325)? mem[1834] : 
                        (N2327)? mem[1898] : 
                        (N2329)? mem[1962] : 
                        (N2331)? mem[2026] : 1'b0;
  assign rdata_o[105] = (N2300)? mem[41] : 
                        (N2302)? mem[105] : 
                        (N2304)? mem[169] : 
                        (N2306)? mem[233] : 
                        (N2308)? mem[297] : 
                        (N2310)? mem[361] : 
                        (N2312)? mem[425] : 
                        (N2314)? mem[489] : 
                        (N2316)? mem[553] : 
                        (N2318)? mem[617] : 
                        (N2320)? mem[681] : 
                        (N2322)? mem[745] : 
                        (N2324)? mem[809] : 
                        (N2326)? mem[873] : 
                        (N2328)? mem[937] : 
                        (N2330)? mem[1001] : 
                        (N2301)? mem[1065] : 
                        (N2303)? mem[1129] : 
                        (N2305)? mem[1193] : 
                        (N2307)? mem[1257] : 
                        (N2309)? mem[1321] : 
                        (N2311)? mem[1385] : 
                        (N2313)? mem[1449] : 
                        (N2315)? mem[1513] : 
                        (N2317)? mem[1577] : 
                        (N2319)? mem[1641] : 
                        (N2321)? mem[1705] : 
                        (N2323)? mem[1769] : 
                        (N2325)? mem[1833] : 
                        (N2327)? mem[1897] : 
                        (N2329)? mem[1961] : 
                        (N2331)? mem[2025] : 1'b0;
  assign rdata_o[104] = (N2300)? mem[40] : 
                        (N2302)? mem[104] : 
                        (N2304)? mem[168] : 
                        (N2306)? mem[232] : 
                        (N2308)? mem[296] : 
                        (N2310)? mem[360] : 
                        (N2312)? mem[424] : 
                        (N2314)? mem[488] : 
                        (N2316)? mem[552] : 
                        (N2318)? mem[616] : 
                        (N2320)? mem[680] : 
                        (N2322)? mem[744] : 
                        (N2324)? mem[808] : 
                        (N2326)? mem[872] : 
                        (N2328)? mem[936] : 
                        (N2330)? mem[1000] : 
                        (N2301)? mem[1064] : 
                        (N2303)? mem[1128] : 
                        (N2305)? mem[1192] : 
                        (N2307)? mem[1256] : 
                        (N2309)? mem[1320] : 
                        (N2311)? mem[1384] : 
                        (N2313)? mem[1448] : 
                        (N2315)? mem[1512] : 
                        (N2317)? mem[1576] : 
                        (N2319)? mem[1640] : 
                        (N2321)? mem[1704] : 
                        (N2323)? mem[1768] : 
                        (N2325)? mem[1832] : 
                        (N2327)? mem[1896] : 
                        (N2329)? mem[1960] : 
                        (N2331)? mem[2024] : 1'b0;
  assign rdata_o[103] = (N2300)? mem[39] : 
                        (N2302)? mem[103] : 
                        (N2304)? mem[167] : 
                        (N2306)? mem[231] : 
                        (N2308)? mem[295] : 
                        (N2310)? mem[359] : 
                        (N2312)? mem[423] : 
                        (N2314)? mem[487] : 
                        (N2316)? mem[551] : 
                        (N2318)? mem[615] : 
                        (N2320)? mem[679] : 
                        (N2322)? mem[743] : 
                        (N2324)? mem[807] : 
                        (N2326)? mem[871] : 
                        (N2328)? mem[935] : 
                        (N2330)? mem[999] : 
                        (N2301)? mem[1063] : 
                        (N2303)? mem[1127] : 
                        (N2305)? mem[1191] : 
                        (N2307)? mem[1255] : 
                        (N2309)? mem[1319] : 
                        (N2311)? mem[1383] : 
                        (N2313)? mem[1447] : 
                        (N2315)? mem[1511] : 
                        (N2317)? mem[1575] : 
                        (N2319)? mem[1639] : 
                        (N2321)? mem[1703] : 
                        (N2323)? mem[1767] : 
                        (N2325)? mem[1831] : 
                        (N2327)? mem[1895] : 
                        (N2329)? mem[1959] : 
                        (N2331)? mem[2023] : 1'b0;
  assign rdata_o[102] = (N2300)? mem[38] : 
                        (N2302)? mem[102] : 
                        (N2304)? mem[166] : 
                        (N2306)? mem[230] : 
                        (N2308)? mem[294] : 
                        (N2310)? mem[358] : 
                        (N2312)? mem[422] : 
                        (N2314)? mem[486] : 
                        (N2316)? mem[550] : 
                        (N2318)? mem[614] : 
                        (N2320)? mem[678] : 
                        (N2322)? mem[742] : 
                        (N2324)? mem[806] : 
                        (N2326)? mem[870] : 
                        (N2328)? mem[934] : 
                        (N2330)? mem[998] : 
                        (N2301)? mem[1062] : 
                        (N2303)? mem[1126] : 
                        (N2305)? mem[1190] : 
                        (N2307)? mem[1254] : 
                        (N2309)? mem[1318] : 
                        (N2311)? mem[1382] : 
                        (N2313)? mem[1446] : 
                        (N2315)? mem[1510] : 
                        (N2317)? mem[1574] : 
                        (N2319)? mem[1638] : 
                        (N2321)? mem[1702] : 
                        (N2323)? mem[1766] : 
                        (N2325)? mem[1830] : 
                        (N2327)? mem[1894] : 
                        (N2329)? mem[1958] : 
                        (N2331)? mem[2022] : 1'b0;
  assign rdata_o[101] = (N2300)? mem[37] : 
                        (N2302)? mem[101] : 
                        (N2304)? mem[165] : 
                        (N2306)? mem[229] : 
                        (N2308)? mem[293] : 
                        (N2310)? mem[357] : 
                        (N2312)? mem[421] : 
                        (N2314)? mem[485] : 
                        (N2316)? mem[549] : 
                        (N2318)? mem[613] : 
                        (N2320)? mem[677] : 
                        (N2322)? mem[741] : 
                        (N2324)? mem[805] : 
                        (N2326)? mem[869] : 
                        (N2328)? mem[933] : 
                        (N2330)? mem[997] : 
                        (N2301)? mem[1061] : 
                        (N2303)? mem[1125] : 
                        (N2305)? mem[1189] : 
                        (N2307)? mem[1253] : 
                        (N2309)? mem[1317] : 
                        (N2311)? mem[1381] : 
                        (N2313)? mem[1445] : 
                        (N2315)? mem[1509] : 
                        (N2317)? mem[1573] : 
                        (N2319)? mem[1637] : 
                        (N2321)? mem[1701] : 
                        (N2323)? mem[1765] : 
                        (N2325)? mem[1829] : 
                        (N2327)? mem[1893] : 
                        (N2329)? mem[1957] : 
                        (N2331)? mem[2021] : 1'b0;
  assign rdata_o[100] = (N2300)? mem[36] : 
                        (N2302)? mem[100] : 
                        (N2304)? mem[164] : 
                        (N2306)? mem[228] : 
                        (N2308)? mem[292] : 
                        (N2310)? mem[356] : 
                        (N2312)? mem[420] : 
                        (N2314)? mem[484] : 
                        (N2316)? mem[548] : 
                        (N2318)? mem[612] : 
                        (N2320)? mem[676] : 
                        (N2322)? mem[740] : 
                        (N2324)? mem[804] : 
                        (N2326)? mem[868] : 
                        (N2328)? mem[932] : 
                        (N2330)? mem[996] : 
                        (N2301)? mem[1060] : 
                        (N2303)? mem[1124] : 
                        (N2305)? mem[1188] : 
                        (N2307)? mem[1252] : 
                        (N2309)? mem[1316] : 
                        (N2311)? mem[1380] : 
                        (N2313)? mem[1444] : 
                        (N2315)? mem[1508] : 
                        (N2317)? mem[1572] : 
                        (N2319)? mem[1636] : 
                        (N2321)? mem[1700] : 
                        (N2323)? mem[1764] : 
                        (N2325)? mem[1828] : 
                        (N2327)? mem[1892] : 
                        (N2329)? mem[1956] : 
                        (N2331)? mem[2020] : 1'b0;
  assign rdata_o[99] = (N2300)? mem[35] : 
                       (N2302)? mem[99] : 
                       (N2304)? mem[163] : 
                       (N2306)? mem[227] : 
                       (N2308)? mem[291] : 
                       (N2310)? mem[355] : 
                       (N2312)? mem[419] : 
                       (N2314)? mem[483] : 
                       (N2316)? mem[547] : 
                       (N2318)? mem[611] : 
                       (N2320)? mem[675] : 
                       (N2322)? mem[739] : 
                       (N2324)? mem[803] : 
                       (N2326)? mem[867] : 
                       (N2328)? mem[931] : 
                       (N2330)? mem[995] : 
                       (N2301)? mem[1059] : 
                       (N2303)? mem[1123] : 
                       (N2305)? mem[1187] : 
                       (N2307)? mem[1251] : 
                       (N2309)? mem[1315] : 
                       (N2311)? mem[1379] : 
                       (N2313)? mem[1443] : 
                       (N2315)? mem[1507] : 
                       (N2317)? mem[1571] : 
                       (N2319)? mem[1635] : 
                       (N2321)? mem[1699] : 
                       (N2323)? mem[1763] : 
                       (N2325)? mem[1827] : 
                       (N2327)? mem[1891] : 
                       (N2329)? mem[1955] : 
                       (N2331)? mem[2019] : 1'b0;
  assign rdata_o[98] = (N2300)? mem[34] : 
                       (N2302)? mem[98] : 
                       (N2304)? mem[162] : 
                       (N2306)? mem[226] : 
                       (N2308)? mem[290] : 
                       (N2310)? mem[354] : 
                       (N2312)? mem[418] : 
                       (N2314)? mem[482] : 
                       (N2316)? mem[546] : 
                       (N2318)? mem[610] : 
                       (N2320)? mem[674] : 
                       (N2322)? mem[738] : 
                       (N2324)? mem[802] : 
                       (N2326)? mem[866] : 
                       (N2328)? mem[930] : 
                       (N2330)? mem[994] : 
                       (N2301)? mem[1058] : 
                       (N2303)? mem[1122] : 
                       (N2305)? mem[1186] : 
                       (N2307)? mem[1250] : 
                       (N2309)? mem[1314] : 
                       (N2311)? mem[1378] : 
                       (N2313)? mem[1442] : 
                       (N2315)? mem[1506] : 
                       (N2317)? mem[1570] : 
                       (N2319)? mem[1634] : 
                       (N2321)? mem[1698] : 
                       (N2323)? mem[1762] : 
                       (N2325)? mem[1826] : 
                       (N2327)? mem[1890] : 
                       (N2329)? mem[1954] : 
                       (N2331)? mem[2018] : 1'b0;
  assign rdata_o[97] = (N2300)? mem[33] : 
                       (N2302)? mem[97] : 
                       (N2304)? mem[161] : 
                       (N2306)? mem[225] : 
                       (N2308)? mem[289] : 
                       (N2310)? mem[353] : 
                       (N2312)? mem[417] : 
                       (N2314)? mem[481] : 
                       (N2316)? mem[545] : 
                       (N2318)? mem[609] : 
                       (N2320)? mem[673] : 
                       (N2322)? mem[737] : 
                       (N2324)? mem[801] : 
                       (N2326)? mem[865] : 
                       (N2328)? mem[929] : 
                       (N2330)? mem[993] : 
                       (N2301)? mem[1057] : 
                       (N2303)? mem[1121] : 
                       (N2305)? mem[1185] : 
                       (N2307)? mem[1249] : 
                       (N2309)? mem[1313] : 
                       (N2311)? mem[1377] : 
                       (N2313)? mem[1441] : 
                       (N2315)? mem[1505] : 
                       (N2317)? mem[1569] : 
                       (N2319)? mem[1633] : 
                       (N2321)? mem[1697] : 
                       (N2323)? mem[1761] : 
                       (N2325)? mem[1825] : 
                       (N2327)? mem[1889] : 
                       (N2329)? mem[1953] : 
                       (N2331)? mem[2017] : 1'b0;
  assign rdata_o[96] = (N2300)? mem[32] : 
                       (N2302)? mem[96] : 
                       (N2304)? mem[160] : 
                       (N2306)? mem[224] : 
                       (N2308)? mem[288] : 
                       (N2310)? mem[352] : 
                       (N2312)? mem[416] : 
                       (N2314)? mem[480] : 
                       (N2316)? mem[544] : 
                       (N2318)? mem[608] : 
                       (N2320)? mem[672] : 
                       (N2322)? mem[736] : 
                       (N2324)? mem[800] : 
                       (N2326)? mem[864] : 
                       (N2328)? mem[928] : 
                       (N2330)? mem[992] : 
                       (N2301)? mem[1056] : 
                       (N2303)? mem[1120] : 
                       (N2305)? mem[1184] : 
                       (N2307)? mem[1248] : 
                       (N2309)? mem[1312] : 
                       (N2311)? mem[1376] : 
                       (N2313)? mem[1440] : 
                       (N2315)? mem[1504] : 
                       (N2317)? mem[1568] : 
                       (N2319)? mem[1632] : 
                       (N2321)? mem[1696] : 
                       (N2323)? mem[1760] : 
                       (N2325)? mem[1824] : 
                       (N2327)? mem[1888] : 
                       (N2329)? mem[1952] : 
                       (N2331)? mem[2016] : 1'b0;
  assign rdata_o[95] = (N2300)? mem[31] : 
                       (N2302)? mem[95] : 
                       (N2304)? mem[159] : 
                       (N2306)? mem[223] : 
                       (N2308)? mem[287] : 
                       (N2310)? mem[351] : 
                       (N2312)? mem[415] : 
                       (N2314)? mem[479] : 
                       (N2316)? mem[543] : 
                       (N2318)? mem[607] : 
                       (N2320)? mem[671] : 
                       (N2322)? mem[735] : 
                       (N2324)? mem[799] : 
                       (N2326)? mem[863] : 
                       (N2328)? mem[927] : 
                       (N2330)? mem[991] : 
                       (N2301)? mem[1055] : 
                       (N2303)? mem[1119] : 
                       (N2305)? mem[1183] : 
                       (N2307)? mem[1247] : 
                       (N2309)? mem[1311] : 
                       (N2311)? mem[1375] : 
                       (N2313)? mem[1439] : 
                       (N2315)? mem[1503] : 
                       (N2317)? mem[1567] : 
                       (N2319)? mem[1631] : 
                       (N2321)? mem[1695] : 
                       (N2323)? mem[1759] : 
                       (N2325)? mem[1823] : 
                       (N2327)? mem[1887] : 
                       (N2329)? mem[1951] : 
                       (N2331)? mem[2015] : 1'b0;
  assign rdata_o[94] = (N2300)? mem[30] : 
                       (N2302)? mem[94] : 
                       (N2304)? mem[158] : 
                       (N2306)? mem[222] : 
                       (N2308)? mem[286] : 
                       (N2310)? mem[350] : 
                       (N2312)? mem[414] : 
                       (N2314)? mem[478] : 
                       (N2316)? mem[542] : 
                       (N2318)? mem[606] : 
                       (N2320)? mem[670] : 
                       (N2322)? mem[734] : 
                       (N2324)? mem[798] : 
                       (N2326)? mem[862] : 
                       (N2328)? mem[926] : 
                       (N2330)? mem[990] : 
                       (N2301)? mem[1054] : 
                       (N2303)? mem[1118] : 
                       (N2305)? mem[1182] : 
                       (N2307)? mem[1246] : 
                       (N2309)? mem[1310] : 
                       (N2311)? mem[1374] : 
                       (N2313)? mem[1438] : 
                       (N2315)? mem[1502] : 
                       (N2317)? mem[1566] : 
                       (N2319)? mem[1630] : 
                       (N2321)? mem[1694] : 
                       (N2323)? mem[1758] : 
                       (N2325)? mem[1822] : 
                       (N2327)? mem[1886] : 
                       (N2329)? mem[1950] : 
                       (N2331)? mem[2014] : 1'b0;
  assign rdata_o[93] = (N2300)? mem[29] : 
                       (N2302)? mem[93] : 
                       (N2304)? mem[157] : 
                       (N2306)? mem[221] : 
                       (N2308)? mem[285] : 
                       (N2310)? mem[349] : 
                       (N2312)? mem[413] : 
                       (N2314)? mem[477] : 
                       (N2316)? mem[541] : 
                       (N2318)? mem[605] : 
                       (N2320)? mem[669] : 
                       (N2322)? mem[733] : 
                       (N2324)? mem[797] : 
                       (N2326)? mem[861] : 
                       (N2328)? mem[925] : 
                       (N2330)? mem[989] : 
                       (N2301)? mem[1053] : 
                       (N2303)? mem[1117] : 
                       (N2305)? mem[1181] : 
                       (N2307)? mem[1245] : 
                       (N2309)? mem[1309] : 
                       (N2311)? mem[1373] : 
                       (N2313)? mem[1437] : 
                       (N2315)? mem[1501] : 
                       (N2317)? mem[1565] : 
                       (N2319)? mem[1629] : 
                       (N2321)? mem[1693] : 
                       (N2323)? mem[1757] : 
                       (N2325)? mem[1821] : 
                       (N2327)? mem[1885] : 
                       (N2329)? mem[1949] : 
                       (N2331)? mem[2013] : 1'b0;
  assign rdata_o[92] = (N2300)? mem[28] : 
                       (N2302)? mem[92] : 
                       (N2304)? mem[156] : 
                       (N2306)? mem[220] : 
                       (N2308)? mem[284] : 
                       (N2310)? mem[348] : 
                       (N2312)? mem[412] : 
                       (N2314)? mem[476] : 
                       (N2316)? mem[540] : 
                       (N2318)? mem[604] : 
                       (N2320)? mem[668] : 
                       (N2322)? mem[732] : 
                       (N2324)? mem[796] : 
                       (N2326)? mem[860] : 
                       (N2328)? mem[924] : 
                       (N2330)? mem[988] : 
                       (N2301)? mem[1052] : 
                       (N2303)? mem[1116] : 
                       (N2305)? mem[1180] : 
                       (N2307)? mem[1244] : 
                       (N2309)? mem[1308] : 
                       (N2311)? mem[1372] : 
                       (N2313)? mem[1436] : 
                       (N2315)? mem[1500] : 
                       (N2317)? mem[1564] : 
                       (N2319)? mem[1628] : 
                       (N2321)? mem[1692] : 
                       (N2323)? mem[1756] : 
                       (N2325)? mem[1820] : 
                       (N2327)? mem[1884] : 
                       (N2329)? mem[1948] : 
                       (N2331)? mem[2012] : 1'b0;
  assign rdata_o[91] = (N2300)? mem[27] : 
                       (N2302)? mem[91] : 
                       (N2304)? mem[155] : 
                       (N2306)? mem[219] : 
                       (N2308)? mem[283] : 
                       (N2310)? mem[347] : 
                       (N2312)? mem[411] : 
                       (N2314)? mem[475] : 
                       (N2316)? mem[539] : 
                       (N2318)? mem[603] : 
                       (N2320)? mem[667] : 
                       (N2322)? mem[731] : 
                       (N2324)? mem[795] : 
                       (N2326)? mem[859] : 
                       (N2328)? mem[923] : 
                       (N2330)? mem[987] : 
                       (N2301)? mem[1051] : 
                       (N2303)? mem[1115] : 
                       (N2305)? mem[1179] : 
                       (N2307)? mem[1243] : 
                       (N2309)? mem[1307] : 
                       (N2311)? mem[1371] : 
                       (N2313)? mem[1435] : 
                       (N2315)? mem[1499] : 
                       (N2317)? mem[1563] : 
                       (N2319)? mem[1627] : 
                       (N2321)? mem[1691] : 
                       (N2323)? mem[1755] : 
                       (N2325)? mem[1819] : 
                       (N2327)? mem[1883] : 
                       (N2329)? mem[1947] : 
                       (N2331)? mem[2011] : 1'b0;
  assign rdata_o[90] = (N2300)? mem[26] : 
                       (N2302)? mem[90] : 
                       (N2304)? mem[154] : 
                       (N2306)? mem[218] : 
                       (N2308)? mem[282] : 
                       (N2310)? mem[346] : 
                       (N2312)? mem[410] : 
                       (N2314)? mem[474] : 
                       (N2316)? mem[538] : 
                       (N2318)? mem[602] : 
                       (N2320)? mem[666] : 
                       (N2322)? mem[730] : 
                       (N2324)? mem[794] : 
                       (N2326)? mem[858] : 
                       (N2328)? mem[922] : 
                       (N2330)? mem[986] : 
                       (N2301)? mem[1050] : 
                       (N2303)? mem[1114] : 
                       (N2305)? mem[1178] : 
                       (N2307)? mem[1242] : 
                       (N2309)? mem[1306] : 
                       (N2311)? mem[1370] : 
                       (N2313)? mem[1434] : 
                       (N2315)? mem[1498] : 
                       (N2317)? mem[1562] : 
                       (N2319)? mem[1626] : 
                       (N2321)? mem[1690] : 
                       (N2323)? mem[1754] : 
                       (N2325)? mem[1818] : 
                       (N2327)? mem[1882] : 
                       (N2329)? mem[1946] : 
                       (N2331)? mem[2010] : 1'b0;
  assign rdata_o[89] = (N2300)? mem[25] : 
                       (N2302)? mem[89] : 
                       (N2304)? mem[153] : 
                       (N2306)? mem[217] : 
                       (N2308)? mem[281] : 
                       (N2310)? mem[345] : 
                       (N2312)? mem[409] : 
                       (N2314)? mem[473] : 
                       (N2316)? mem[537] : 
                       (N2318)? mem[601] : 
                       (N2320)? mem[665] : 
                       (N2322)? mem[729] : 
                       (N2324)? mem[793] : 
                       (N2326)? mem[857] : 
                       (N2328)? mem[921] : 
                       (N2330)? mem[985] : 
                       (N2301)? mem[1049] : 
                       (N2303)? mem[1113] : 
                       (N2305)? mem[1177] : 
                       (N2307)? mem[1241] : 
                       (N2309)? mem[1305] : 
                       (N2311)? mem[1369] : 
                       (N2313)? mem[1433] : 
                       (N2315)? mem[1497] : 
                       (N2317)? mem[1561] : 
                       (N2319)? mem[1625] : 
                       (N2321)? mem[1689] : 
                       (N2323)? mem[1753] : 
                       (N2325)? mem[1817] : 
                       (N2327)? mem[1881] : 
                       (N2329)? mem[1945] : 
                       (N2331)? mem[2009] : 1'b0;
  assign rdata_o[88] = (N2300)? mem[24] : 
                       (N2302)? mem[88] : 
                       (N2304)? mem[152] : 
                       (N2306)? mem[216] : 
                       (N2308)? mem[280] : 
                       (N2310)? mem[344] : 
                       (N2312)? mem[408] : 
                       (N2314)? mem[472] : 
                       (N2316)? mem[536] : 
                       (N2318)? mem[600] : 
                       (N2320)? mem[664] : 
                       (N2322)? mem[728] : 
                       (N2324)? mem[792] : 
                       (N2326)? mem[856] : 
                       (N2328)? mem[920] : 
                       (N2330)? mem[984] : 
                       (N2301)? mem[1048] : 
                       (N2303)? mem[1112] : 
                       (N2305)? mem[1176] : 
                       (N2307)? mem[1240] : 
                       (N2309)? mem[1304] : 
                       (N2311)? mem[1368] : 
                       (N2313)? mem[1432] : 
                       (N2315)? mem[1496] : 
                       (N2317)? mem[1560] : 
                       (N2319)? mem[1624] : 
                       (N2321)? mem[1688] : 
                       (N2323)? mem[1752] : 
                       (N2325)? mem[1816] : 
                       (N2327)? mem[1880] : 
                       (N2329)? mem[1944] : 
                       (N2331)? mem[2008] : 1'b0;
  assign rdata_o[87] = (N2300)? mem[23] : 
                       (N2302)? mem[87] : 
                       (N2304)? mem[151] : 
                       (N2306)? mem[215] : 
                       (N2308)? mem[279] : 
                       (N2310)? mem[343] : 
                       (N2312)? mem[407] : 
                       (N2314)? mem[471] : 
                       (N2316)? mem[535] : 
                       (N2318)? mem[599] : 
                       (N2320)? mem[663] : 
                       (N2322)? mem[727] : 
                       (N2324)? mem[791] : 
                       (N2326)? mem[855] : 
                       (N2328)? mem[919] : 
                       (N2330)? mem[983] : 
                       (N2301)? mem[1047] : 
                       (N2303)? mem[1111] : 
                       (N2305)? mem[1175] : 
                       (N2307)? mem[1239] : 
                       (N2309)? mem[1303] : 
                       (N2311)? mem[1367] : 
                       (N2313)? mem[1431] : 
                       (N2315)? mem[1495] : 
                       (N2317)? mem[1559] : 
                       (N2319)? mem[1623] : 
                       (N2321)? mem[1687] : 
                       (N2323)? mem[1751] : 
                       (N2325)? mem[1815] : 
                       (N2327)? mem[1879] : 
                       (N2329)? mem[1943] : 
                       (N2331)? mem[2007] : 1'b0;
  assign rdata_o[86] = (N2300)? mem[22] : 
                       (N2302)? mem[86] : 
                       (N2304)? mem[150] : 
                       (N2306)? mem[214] : 
                       (N2308)? mem[278] : 
                       (N2310)? mem[342] : 
                       (N2312)? mem[406] : 
                       (N2314)? mem[470] : 
                       (N2316)? mem[534] : 
                       (N2318)? mem[598] : 
                       (N2320)? mem[662] : 
                       (N2322)? mem[726] : 
                       (N2324)? mem[790] : 
                       (N2326)? mem[854] : 
                       (N2328)? mem[918] : 
                       (N2330)? mem[982] : 
                       (N2301)? mem[1046] : 
                       (N2303)? mem[1110] : 
                       (N2305)? mem[1174] : 
                       (N2307)? mem[1238] : 
                       (N2309)? mem[1302] : 
                       (N2311)? mem[1366] : 
                       (N2313)? mem[1430] : 
                       (N2315)? mem[1494] : 
                       (N2317)? mem[1558] : 
                       (N2319)? mem[1622] : 
                       (N2321)? mem[1686] : 
                       (N2323)? mem[1750] : 
                       (N2325)? mem[1814] : 
                       (N2327)? mem[1878] : 
                       (N2329)? mem[1942] : 
                       (N2331)? mem[2006] : 1'b0;
  assign rdata_o[85] = (N2300)? mem[21] : 
                       (N2302)? mem[85] : 
                       (N2304)? mem[149] : 
                       (N2306)? mem[213] : 
                       (N2308)? mem[277] : 
                       (N2310)? mem[341] : 
                       (N2312)? mem[405] : 
                       (N2314)? mem[469] : 
                       (N2316)? mem[533] : 
                       (N2318)? mem[597] : 
                       (N2320)? mem[661] : 
                       (N2322)? mem[725] : 
                       (N2324)? mem[789] : 
                       (N2326)? mem[853] : 
                       (N2328)? mem[917] : 
                       (N2330)? mem[981] : 
                       (N2301)? mem[1045] : 
                       (N2303)? mem[1109] : 
                       (N2305)? mem[1173] : 
                       (N2307)? mem[1237] : 
                       (N2309)? mem[1301] : 
                       (N2311)? mem[1365] : 
                       (N2313)? mem[1429] : 
                       (N2315)? mem[1493] : 
                       (N2317)? mem[1557] : 
                       (N2319)? mem[1621] : 
                       (N2321)? mem[1685] : 
                       (N2323)? mem[1749] : 
                       (N2325)? mem[1813] : 
                       (N2327)? mem[1877] : 
                       (N2329)? mem[1941] : 
                       (N2331)? mem[2005] : 1'b0;
  assign rdata_o[84] = (N2300)? mem[20] : 
                       (N2302)? mem[84] : 
                       (N2304)? mem[148] : 
                       (N2306)? mem[212] : 
                       (N2308)? mem[276] : 
                       (N2310)? mem[340] : 
                       (N2312)? mem[404] : 
                       (N2314)? mem[468] : 
                       (N2316)? mem[532] : 
                       (N2318)? mem[596] : 
                       (N2320)? mem[660] : 
                       (N2322)? mem[724] : 
                       (N2324)? mem[788] : 
                       (N2326)? mem[852] : 
                       (N2328)? mem[916] : 
                       (N2330)? mem[980] : 
                       (N2301)? mem[1044] : 
                       (N2303)? mem[1108] : 
                       (N2305)? mem[1172] : 
                       (N2307)? mem[1236] : 
                       (N2309)? mem[1300] : 
                       (N2311)? mem[1364] : 
                       (N2313)? mem[1428] : 
                       (N2315)? mem[1492] : 
                       (N2317)? mem[1556] : 
                       (N2319)? mem[1620] : 
                       (N2321)? mem[1684] : 
                       (N2323)? mem[1748] : 
                       (N2325)? mem[1812] : 
                       (N2327)? mem[1876] : 
                       (N2329)? mem[1940] : 
                       (N2331)? mem[2004] : 1'b0;
  assign rdata_o[83] = (N2300)? mem[19] : 
                       (N2302)? mem[83] : 
                       (N2304)? mem[147] : 
                       (N2306)? mem[211] : 
                       (N2308)? mem[275] : 
                       (N2310)? mem[339] : 
                       (N2312)? mem[403] : 
                       (N2314)? mem[467] : 
                       (N2316)? mem[531] : 
                       (N2318)? mem[595] : 
                       (N2320)? mem[659] : 
                       (N2322)? mem[723] : 
                       (N2324)? mem[787] : 
                       (N2326)? mem[851] : 
                       (N2328)? mem[915] : 
                       (N2330)? mem[979] : 
                       (N2301)? mem[1043] : 
                       (N2303)? mem[1107] : 
                       (N2305)? mem[1171] : 
                       (N2307)? mem[1235] : 
                       (N2309)? mem[1299] : 
                       (N2311)? mem[1363] : 
                       (N2313)? mem[1427] : 
                       (N2315)? mem[1491] : 
                       (N2317)? mem[1555] : 
                       (N2319)? mem[1619] : 
                       (N2321)? mem[1683] : 
                       (N2323)? mem[1747] : 
                       (N2325)? mem[1811] : 
                       (N2327)? mem[1875] : 
                       (N2329)? mem[1939] : 
                       (N2331)? mem[2003] : 1'b0;
  assign rdata_o[82] = (N2300)? mem[18] : 
                       (N2302)? mem[82] : 
                       (N2304)? mem[146] : 
                       (N2306)? mem[210] : 
                       (N2308)? mem[274] : 
                       (N2310)? mem[338] : 
                       (N2312)? mem[402] : 
                       (N2314)? mem[466] : 
                       (N2316)? mem[530] : 
                       (N2318)? mem[594] : 
                       (N2320)? mem[658] : 
                       (N2322)? mem[722] : 
                       (N2324)? mem[786] : 
                       (N2326)? mem[850] : 
                       (N2328)? mem[914] : 
                       (N2330)? mem[978] : 
                       (N2301)? mem[1042] : 
                       (N2303)? mem[1106] : 
                       (N2305)? mem[1170] : 
                       (N2307)? mem[1234] : 
                       (N2309)? mem[1298] : 
                       (N2311)? mem[1362] : 
                       (N2313)? mem[1426] : 
                       (N2315)? mem[1490] : 
                       (N2317)? mem[1554] : 
                       (N2319)? mem[1618] : 
                       (N2321)? mem[1682] : 
                       (N2323)? mem[1746] : 
                       (N2325)? mem[1810] : 
                       (N2327)? mem[1874] : 
                       (N2329)? mem[1938] : 
                       (N2331)? mem[2002] : 1'b0;
  assign rdata_o[81] = (N2300)? mem[17] : 
                       (N2302)? mem[81] : 
                       (N2304)? mem[145] : 
                       (N2306)? mem[209] : 
                       (N2308)? mem[273] : 
                       (N2310)? mem[337] : 
                       (N2312)? mem[401] : 
                       (N2314)? mem[465] : 
                       (N2316)? mem[529] : 
                       (N2318)? mem[593] : 
                       (N2320)? mem[657] : 
                       (N2322)? mem[721] : 
                       (N2324)? mem[785] : 
                       (N2326)? mem[849] : 
                       (N2328)? mem[913] : 
                       (N2330)? mem[977] : 
                       (N2301)? mem[1041] : 
                       (N2303)? mem[1105] : 
                       (N2305)? mem[1169] : 
                       (N2307)? mem[1233] : 
                       (N2309)? mem[1297] : 
                       (N2311)? mem[1361] : 
                       (N2313)? mem[1425] : 
                       (N2315)? mem[1489] : 
                       (N2317)? mem[1553] : 
                       (N2319)? mem[1617] : 
                       (N2321)? mem[1681] : 
                       (N2323)? mem[1745] : 
                       (N2325)? mem[1809] : 
                       (N2327)? mem[1873] : 
                       (N2329)? mem[1937] : 
                       (N2331)? mem[2001] : 1'b0;
  assign rdata_o[80] = (N2300)? mem[16] : 
                       (N2302)? mem[80] : 
                       (N2304)? mem[144] : 
                       (N2306)? mem[208] : 
                       (N2308)? mem[272] : 
                       (N2310)? mem[336] : 
                       (N2312)? mem[400] : 
                       (N2314)? mem[464] : 
                       (N2316)? mem[528] : 
                       (N2318)? mem[592] : 
                       (N2320)? mem[656] : 
                       (N2322)? mem[720] : 
                       (N2324)? mem[784] : 
                       (N2326)? mem[848] : 
                       (N2328)? mem[912] : 
                       (N2330)? mem[976] : 
                       (N2301)? mem[1040] : 
                       (N2303)? mem[1104] : 
                       (N2305)? mem[1168] : 
                       (N2307)? mem[1232] : 
                       (N2309)? mem[1296] : 
                       (N2311)? mem[1360] : 
                       (N2313)? mem[1424] : 
                       (N2315)? mem[1488] : 
                       (N2317)? mem[1552] : 
                       (N2319)? mem[1616] : 
                       (N2321)? mem[1680] : 
                       (N2323)? mem[1744] : 
                       (N2325)? mem[1808] : 
                       (N2327)? mem[1872] : 
                       (N2329)? mem[1936] : 
                       (N2331)? mem[2000] : 1'b0;
  assign rdata_o[79] = (N2300)? mem[15] : 
                       (N2302)? mem[79] : 
                       (N2304)? mem[143] : 
                       (N2306)? mem[207] : 
                       (N2308)? mem[271] : 
                       (N2310)? mem[335] : 
                       (N2312)? mem[399] : 
                       (N2314)? mem[463] : 
                       (N2316)? mem[527] : 
                       (N2318)? mem[591] : 
                       (N2320)? mem[655] : 
                       (N2322)? mem[719] : 
                       (N2324)? mem[783] : 
                       (N2326)? mem[847] : 
                       (N2328)? mem[911] : 
                       (N2330)? mem[975] : 
                       (N2301)? mem[1039] : 
                       (N2303)? mem[1103] : 
                       (N2305)? mem[1167] : 
                       (N2307)? mem[1231] : 
                       (N2309)? mem[1295] : 
                       (N2311)? mem[1359] : 
                       (N2313)? mem[1423] : 
                       (N2315)? mem[1487] : 
                       (N2317)? mem[1551] : 
                       (N2319)? mem[1615] : 
                       (N2321)? mem[1679] : 
                       (N2323)? mem[1743] : 
                       (N2325)? mem[1807] : 
                       (N2327)? mem[1871] : 
                       (N2329)? mem[1935] : 
                       (N2331)? mem[1999] : 1'b0;
  assign rdata_o[78] = (N2300)? mem[14] : 
                       (N2302)? mem[78] : 
                       (N2304)? mem[142] : 
                       (N2306)? mem[206] : 
                       (N2308)? mem[270] : 
                       (N2310)? mem[334] : 
                       (N2312)? mem[398] : 
                       (N2314)? mem[462] : 
                       (N2316)? mem[526] : 
                       (N2318)? mem[590] : 
                       (N2320)? mem[654] : 
                       (N2322)? mem[718] : 
                       (N2324)? mem[782] : 
                       (N2326)? mem[846] : 
                       (N2328)? mem[910] : 
                       (N2330)? mem[974] : 
                       (N2301)? mem[1038] : 
                       (N2303)? mem[1102] : 
                       (N2305)? mem[1166] : 
                       (N2307)? mem[1230] : 
                       (N2309)? mem[1294] : 
                       (N2311)? mem[1358] : 
                       (N2313)? mem[1422] : 
                       (N2315)? mem[1486] : 
                       (N2317)? mem[1550] : 
                       (N2319)? mem[1614] : 
                       (N2321)? mem[1678] : 
                       (N2323)? mem[1742] : 
                       (N2325)? mem[1806] : 
                       (N2327)? mem[1870] : 
                       (N2329)? mem[1934] : 
                       (N2331)? mem[1998] : 1'b0;
  assign rdata_o[77] = (N2300)? mem[13] : 
                       (N2302)? mem[77] : 
                       (N2304)? mem[141] : 
                       (N2306)? mem[205] : 
                       (N2308)? mem[269] : 
                       (N2310)? mem[333] : 
                       (N2312)? mem[397] : 
                       (N2314)? mem[461] : 
                       (N2316)? mem[525] : 
                       (N2318)? mem[589] : 
                       (N2320)? mem[653] : 
                       (N2322)? mem[717] : 
                       (N2324)? mem[781] : 
                       (N2326)? mem[845] : 
                       (N2328)? mem[909] : 
                       (N2330)? mem[973] : 
                       (N2301)? mem[1037] : 
                       (N2303)? mem[1101] : 
                       (N2305)? mem[1165] : 
                       (N2307)? mem[1229] : 
                       (N2309)? mem[1293] : 
                       (N2311)? mem[1357] : 
                       (N2313)? mem[1421] : 
                       (N2315)? mem[1485] : 
                       (N2317)? mem[1549] : 
                       (N2319)? mem[1613] : 
                       (N2321)? mem[1677] : 
                       (N2323)? mem[1741] : 
                       (N2325)? mem[1805] : 
                       (N2327)? mem[1869] : 
                       (N2329)? mem[1933] : 
                       (N2331)? mem[1997] : 1'b0;
  assign rdata_o[76] = (N2300)? mem[12] : 
                       (N2302)? mem[76] : 
                       (N2304)? mem[140] : 
                       (N2306)? mem[204] : 
                       (N2308)? mem[268] : 
                       (N2310)? mem[332] : 
                       (N2312)? mem[396] : 
                       (N2314)? mem[460] : 
                       (N2316)? mem[524] : 
                       (N2318)? mem[588] : 
                       (N2320)? mem[652] : 
                       (N2322)? mem[716] : 
                       (N2324)? mem[780] : 
                       (N2326)? mem[844] : 
                       (N2328)? mem[908] : 
                       (N2330)? mem[972] : 
                       (N2301)? mem[1036] : 
                       (N2303)? mem[1100] : 
                       (N2305)? mem[1164] : 
                       (N2307)? mem[1228] : 
                       (N2309)? mem[1292] : 
                       (N2311)? mem[1356] : 
                       (N2313)? mem[1420] : 
                       (N2315)? mem[1484] : 
                       (N2317)? mem[1548] : 
                       (N2319)? mem[1612] : 
                       (N2321)? mem[1676] : 
                       (N2323)? mem[1740] : 
                       (N2325)? mem[1804] : 
                       (N2327)? mem[1868] : 
                       (N2329)? mem[1932] : 
                       (N2331)? mem[1996] : 1'b0;
  assign rdata_o[75] = (N2300)? mem[11] : 
                       (N2302)? mem[75] : 
                       (N2304)? mem[139] : 
                       (N2306)? mem[203] : 
                       (N2308)? mem[267] : 
                       (N2310)? mem[331] : 
                       (N2312)? mem[395] : 
                       (N2314)? mem[459] : 
                       (N2316)? mem[523] : 
                       (N2318)? mem[587] : 
                       (N2320)? mem[651] : 
                       (N2322)? mem[715] : 
                       (N2324)? mem[779] : 
                       (N2326)? mem[843] : 
                       (N2328)? mem[907] : 
                       (N2330)? mem[971] : 
                       (N2301)? mem[1035] : 
                       (N2303)? mem[1099] : 
                       (N2305)? mem[1163] : 
                       (N2307)? mem[1227] : 
                       (N2309)? mem[1291] : 
                       (N2311)? mem[1355] : 
                       (N2313)? mem[1419] : 
                       (N2315)? mem[1483] : 
                       (N2317)? mem[1547] : 
                       (N2319)? mem[1611] : 
                       (N2321)? mem[1675] : 
                       (N2323)? mem[1739] : 
                       (N2325)? mem[1803] : 
                       (N2327)? mem[1867] : 
                       (N2329)? mem[1931] : 
                       (N2331)? mem[1995] : 1'b0;
  assign rdata_o[74] = (N2300)? mem[10] : 
                       (N2302)? mem[74] : 
                       (N2304)? mem[138] : 
                       (N2306)? mem[202] : 
                       (N2308)? mem[266] : 
                       (N2310)? mem[330] : 
                       (N2312)? mem[394] : 
                       (N2314)? mem[458] : 
                       (N2316)? mem[522] : 
                       (N2318)? mem[586] : 
                       (N2320)? mem[650] : 
                       (N2322)? mem[714] : 
                       (N2324)? mem[778] : 
                       (N2326)? mem[842] : 
                       (N2328)? mem[906] : 
                       (N2330)? mem[970] : 
                       (N2301)? mem[1034] : 
                       (N2303)? mem[1098] : 
                       (N2305)? mem[1162] : 
                       (N2307)? mem[1226] : 
                       (N2309)? mem[1290] : 
                       (N2311)? mem[1354] : 
                       (N2313)? mem[1418] : 
                       (N2315)? mem[1482] : 
                       (N2317)? mem[1546] : 
                       (N2319)? mem[1610] : 
                       (N2321)? mem[1674] : 
                       (N2323)? mem[1738] : 
                       (N2325)? mem[1802] : 
                       (N2327)? mem[1866] : 
                       (N2329)? mem[1930] : 
                       (N2331)? mem[1994] : 1'b0;
  assign rdata_o[73] = (N2300)? mem[9] : 
                       (N2302)? mem[73] : 
                       (N2304)? mem[137] : 
                       (N2306)? mem[201] : 
                       (N2308)? mem[265] : 
                       (N2310)? mem[329] : 
                       (N2312)? mem[393] : 
                       (N2314)? mem[457] : 
                       (N2316)? mem[521] : 
                       (N2318)? mem[585] : 
                       (N2320)? mem[649] : 
                       (N2322)? mem[713] : 
                       (N2324)? mem[777] : 
                       (N2326)? mem[841] : 
                       (N2328)? mem[905] : 
                       (N2330)? mem[969] : 
                       (N2301)? mem[1033] : 
                       (N2303)? mem[1097] : 
                       (N2305)? mem[1161] : 
                       (N2307)? mem[1225] : 
                       (N2309)? mem[1289] : 
                       (N2311)? mem[1353] : 
                       (N2313)? mem[1417] : 
                       (N2315)? mem[1481] : 
                       (N2317)? mem[1545] : 
                       (N2319)? mem[1609] : 
                       (N2321)? mem[1673] : 
                       (N2323)? mem[1737] : 
                       (N2325)? mem[1801] : 
                       (N2327)? mem[1865] : 
                       (N2329)? mem[1929] : 
                       (N2331)? mem[1993] : 1'b0;
  assign rdata_o[72] = (N2300)? mem[8] : 
                       (N2302)? mem[72] : 
                       (N2304)? mem[136] : 
                       (N2306)? mem[200] : 
                       (N2308)? mem[264] : 
                       (N2310)? mem[328] : 
                       (N2312)? mem[392] : 
                       (N2314)? mem[456] : 
                       (N2316)? mem[520] : 
                       (N2318)? mem[584] : 
                       (N2320)? mem[648] : 
                       (N2322)? mem[712] : 
                       (N2324)? mem[776] : 
                       (N2326)? mem[840] : 
                       (N2328)? mem[904] : 
                       (N2330)? mem[968] : 
                       (N2301)? mem[1032] : 
                       (N2303)? mem[1096] : 
                       (N2305)? mem[1160] : 
                       (N2307)? mem[1224] : 
                       (N2309)? mem[1288] : 
                       (N2311)? mem[1352] : 
                       (N2313)? mem[1416] : 
                       (N2315)? mem[1480] : 
                       (N2317)? mem[1544] : 
                       (N2319)? mem[1608] : 
                       (N2321)? mem[1672] : 
                       (N2323)? mem[1736] : 
                       (N2325)? mem[1800] : 
                       (N2327)? mem[1864] : 
                       (N2329)? mem[1928] : 
                       (N2331)? mem[1992] : 1'b0;
  assign rdata_o[71] = (N2300)? mem[7] : 
                       (N2302)? mem[71] : 
                       (N2304)? mem[135] : 
                       (N2306)? mem[199] : 
                       (N2308)? mem[263] : 
                       (N2310)? mem[327] : 
                       (N2312)? mem[391] : 
                       (N2314)? mem[455] : 
                       (N2316)? mem[519] : 
                       (N2318)? mem[583] : 
                       (N2320)? mem[647] : 
                       (N2322)? mem[711] : 
                       (N2324)? mem[775] : 
                       (N2326)? mem[839] : 
                       (N2328)? mem[903] : 
                       (N2330)? mem[967] : 
                       (N2301)? mem[1031] : 
                       (N2303)? mem[1095] : 
                       (N2305)? mem[1159] : 
                       (N2307)? mem[1223] : 
                       (N2309)? mem[1287] : 
                       (N2311)? mem[1351] : 
                       (N2313)? mem[1415] : 
                       (N2315)? mem[1479] : 
                       (N2317)? mem[1543] : 
                       (N2319)? mem[1607] : 
                       (N2321)? mem[1671] : 
                       (N2323)? mem[1735] : 
                       (N2325)? mem[1799] : 
                       (N2327)? mem[1863] : 
                       (N2329)? mem[1927] : 
                       (N2331)? mem[1991] : 1'b0;
  assign rdata_o[70] = (N2300)? mem[6] : 
                       (N2302)? mem[70] : 
                       (N2304)? mem[134] : 
                       (N2306)? mem[198] : 
                       (N2308)? mem[262] : 
                       (N2310)? mem[326] : 
                       (N2312)? mem[390] : 
                       (N2314)? mem[454] : 
                       (N2316)? mem[518] : 
                       (N2318)? mem[582] : 
                       (N2320)? mem[646] : 
                       (N2322)? mem[710] : 
                       (N2324)? mem[774] : 
                       (N2326)? mem[838] : 
                       (N2328)? mem[902] : 
                       (N2330)? mem[966] : 
                       (N2301)? mem[1030] : 
                       (N2303)? mem[1094] : 
                       (N2305)? mem[1158] : 
                       (N2307)? mem[1222] : 
                       (N2309)? mem[1286] : 
                       (N2311)? mem[1350] : 
                       (N2313)? mem[1414] : 
                       (N2315)? mem[1478] : 
                       (N2317)? mem[1542] : 
                       (N2319)? mem[1606] : 
                       (N2321)? mem[1670] : 
                       (N2323)? mem[1734] : 
                       (N2325)? mem[1798] : 
                       (N2327)? mem[1862] : 
                       (N2329)? mem[1926] : 
                       (N2331)? mem[1990] : 1'b0;
  assign rdata_o[69] = (N2300)? mem[5] : 
                       (N2302)? mem[69] : 
                       (N2304)? mem[133] : 
                       (N2306)? mem[197] : 
                       (N2308)? mem[261] : 
                       (N2310)? mem[325] : 
                       (N2312)? mem[389] : 
                       (N2314)? mem[453] : 
                       (N2316)? mem[517] : 
                       (N2318)? mem[581] : 
                       (N2320)? mem[645] : 
                       (N2322)? mem[709] : 
                       (N2324)? mem[773] : 
                       (N2326)? mem[837] : 
                       (N2328)? mem[901] : 
                       (N2330)? mem[965] : 
                       (N2301)? mem[1029] : 
                       (N2303)? mem[1093] : 
                       (N2305)? mem[1157] : 
                       (N2307)? mem[1221] : 
                       (N2309)? mem[1285] : 
                       (N2311)? mem[1349] : 
                       (N2313)? mem[1413] : 
                       (N2315)? mem[1477] : 
                       (N2317)? mem[1541] : 
                       (N2319)? mem[1605] : 
                       (N2321)? mem[1669] : 
                       (N2323)? mem[1733] : 
                       (N2325)? mem[1797] : 
                       (N2327)? mem[1861] : 
                       (N2329)? mem[1925] : 
                       (N2331)? mem[1989] : 1'b0;
  assign rdata_o[68] = (N2300)? mem[4] : 
                       (N2302)? mem[68] : 
                       (N2304)? mem[132] : 
                       (N2306)? mem[196] : 
                       (N2308)? mem[260] : 
                       (N2310)? mem[324] : 
                       (N2312)? mem[388] : 
                       (N2314)? mem[452] : 
                       (N2316)? mem[516] : 
                       (N2318)? mem[580] : 
                       (N2320)? mem[644] : 
                       (N2322)? mem[708] : 
                       (N2324)? mem[772] : 
                       (N2326)? mem[836] : 
                       (N2328)? mem[900] : 
                       (N2330)? mem[964] : 
                       (N2301)? mem[1028] : 
                       (N2303)? mem[1092] : 
                       (N2305)? mem[1156] : 
                       (N2307)? mem[1220] : 
                       (N2309)? mem[1284] : 
                       (N2311)? mem[1348] : 
                       (N2313)? mem[1412] : 
                       (N2315)? mem[1476] : 
                       (N2317)? mem[1540] : 
                       (N2319)? mem[1604] : 
                       (N2321)? mem[1668] : 
                       (N2323)? mem[1732] : 
                       (N2325)? mem[1796] : 
                       (N2327)? mem[1860] : 
                       (N2329)? mem[1924] : 
                       (N2331)? mem[1988] : 1'b0;
  assign rdata_o[67] = (N2300)? mem[3] : 
                       (N2302)? mem[67] : 
                       (N2304)? mem[131] : 
                       (N2306)? mem[195] : 
                       (N2308)? mem[259] : 
                       (N2310)? mem[323] : 
                       (N2312)? mem[387] : 
                       (N2314)? mem[451] : 
                       (N2316)? mem[515] : 
                       (N2318)? mem[579] : 
                       (N2320)? mem[643] : 
                       (N2322)? mem[707] : 
                       (N2324)? mem[771] : 
                       (N2326)? mem[835] : 
                       (N2328)? mem[899] : 
                       (N2330)? mem[963] : 
                       (N2301)? mem[1027] : 
                       (N2303)? mem[1091] : 
                       (N2305)? mem[1155] : 
                       (N2307)? mem[1219] : 
                       (N2309)? mem[1283] : 
                       (N2311)? mem[1347] : 
                       (N2313)? mem[1411] : 
                       (N2315)? mem[1475] : 
                       (N2317)? mem[1539] : 
                       (N2319)? mem[1603] : 
                       (N2321)? mem[1667] : 
                       (N2323)? mem[1731] : 
                       (N2325)? mem[1795] : 
                       (N2327)? mem[1859] : 
                       (N2329)? mem[1923] : 
                       (N2331)? mem[1987] : 1'b0;
  assign rdata_o[66] = (N2300)? mem[2] : 
                       (N2302)? mem[66] : 
                       (N2304)? mem[130] : 
                       (N2306)? mem[194] : 
                       (N2308)? mem[258] : 
                       (N2310)? mem[322] : 
                       (N2312)? mem[386] : 
                       (N2314)? mem[450] : 
                       (N2316)? mem[514] : 
                       (N2318)? mem[578] : 
                       (N2320)? mem[642] : 
                       (N2322)? mem[706] : 
                       (N2324)? mem[770] : 
                       (N2326)? mem[834] : 
                       (N2328)? mem[898] : 
                       (N2330)? mem[962] : 
                       (N2301)? mem[1026] : 
                       (N2303)? mem[1090] : 
                       (N2305)? mem[1154] : 
                       (N2307)? mem[1218] : 
                       (N2309)? mem[1282] : 
                       (N2311)? mem[1346] : 
                       (N2313)? mem[1410] : 
                       (N2315)? mem[1474] : 
                       (N2317)? mem[1538] : 
                       (N2319)? mem[1602] : 
                       (N2321)? mem[1666] : 
                       (N2323)? mem[1730] : 
                       (N2325)? mem[1794] : 
                       (N2327)? mem[1858] : 
                       (N2329)? mem[1922] : 
                       (N2331)? mem[1986] : 1'b0;
  assign rdata_o[65] = (N2300)? mem[1] : 
                       (N2302)? mem[65] : 
                       (N2304)? mem[129] : 
                       (N2306)? mem[193] : 
                       (N2308)? mem[257] : 
                       (N2310)? mem[321] : 
                       (N2312)? mem[385] : 
                       (N2314)? mem[449] : 
                       (N2316)? mem[513] : 
                       (N2318)? mem[577] : 
                       (N2320)? mem[641] : 
                       (N2322)? mem[705] : 
                       (N2324)? mem[769] : 
                       (N2326)? mem[833] : 
                       (N2328)? mem[897] : 
                       (N2330)? mem[961] : 
                       (N2301)? mem[1025] : 
                       (N2303)? mem[1089] : 
                       (N2305)? mem[1153] : 
                       (N2307)? mem[1217] : 
                       (N2309)? mem[1281] : 
                       (N2311)? mem[1345] : 
                       (N2313)? mem[1409] : 
                       (N2315)? mem[1473] : 
                       (N2317)? mem[1537] : 
                       (N2319)? mem[1601] : 
                       (N2321)? mem[1665] : 
                       (N2323)? mem[1729] : 
                       (N2325)? mem[1793] : 
                       (N2327)? mem[1857] : 
                       (N2329)? mem[1921] : 
                       (N2331)? mem[1985] : 1'b0;
  assign rdata_o[64] = (N2300)? mem[0] : 
                       (N2302)? mem[64] : 
                       (N2304)? mem[128] : 
                       (N2306)? mem[192] : 
                       (N2308)? mem[256] : 
                       (N2310)? mem[320] : 
                       (N2312)? mem[384] : 
                       (N2314)? mem[448] : 
                       (N2316)? mem[512] : 
                       (N2318)? mem[576] : 
                       (N2320)? mem[640] : 
                       (N2322)? mem[704] : 
                       (N2324)? mem[768] : 
                       (N2326)? mem[832] : 
                       (N2328)? mem[896] : 
                       (N2330)? mem[960] : 
                       (N2301)? mem[1024] : 
                       (N2303)? mem[1088] : 
                       (N2305)? mem[1152] : 
                       (N2307)? mem[1216] : 
                       (N2309)? mem[1280] : 
                       (N2311)? mem[1344] : 
                       (N2313)? mem[1408] : 
                       (N2315)? mem[1472] : 
                       (N2317)? mem[1536] : 
                       (N2319)? mem[1600] : 
                       (N2321)? mem[1664] : 
                       (N2323)? mem[1728] : 
                       (N2325)? mem[1792] : 
                       (N2327)? mem[1856] : 
                       (N2329)? mem[1920] : 
                       (N2331)? mem[1984] : 1'b0;
  assign N2332 = waddr_i[8] & waddr_i[9];
  assign N2333 = waddr_i[7] & N2332;
  assign N2334 = waddr_i[6] & N2333;
  assign N2335 = waddr_i[5] & N2334;
  assign N2336 = ~waddr_i[9];
  assign N2337 = ~waddr_i[8];
  assign N2338 = ~waddr_i[7];
  assign N2339 = ~waddr_i[6];
  assign N2340 = N2337 | N2336;
  assign N2341 = N2338 | N2340;
  assign N2342 = N2339 | N2341;
  assign N2343 = waddr_i[5] | N2342;
  assign N2344 = ~N2343;
  assign N2345 = ~waddr_i[5];
  assign N2346 = waddr_i[6] | N2341;
  assign N2347 = N2345 | N2346;
  assign N2348 = ~N2347;
  assign N2349 = waddr_i[5] | N2346;
  assign N2350 = ~N2349;
  assign N2351 = waddr_i[7] | N2340;
  assign N2352 = N2339 | N2351;
  assign N2353 = N2345 | N2352;
  assign N2354 = ~N2353;
  assign N2355 = waddr_i[5] | N2352;
  assign N2356 = ~N2355;
  assign N2357 = waddr_i[6] | N2351;
  assign N2358 = N2345 | N2357;
  assign N2359 = ~N2358;
  assign N2360 = waddr_i[5] | N2357;
  assign N2361 = ~N2360;
  assign N2362 = waddr_i[8] | N2336;
  assign N2363 = N2338 | N2362;
  assign N2364 = N2339 | N2363;
  assign N2365 = N2345 | N2364;
  assign N2366 = ~N2365;
  assign N2367 = waddr_i[5] | N2364;
  assign N2368 = ~N2367;
  assign N2369 = waddr_i[6] | N2363;
  assign N2370 = N2345 | N2369;
  assign N2371 = ~N2370;
  assign N2372 = waddr_i[5] | N2369;
  assign N2373 = ~N2372;
  assign N2374 = waddr_i[7] | N2362;
  assign N2375 = N2339 | N2374;
  assign N2376 = N2345 | N2375;
  assign N2377 = ~N2376;
  assign N2378 = waddr_i[5] | N2375;
  assign N2379 = ~N2378;
  assign N2380 = waddr_i[6] | N2374;
  assign N2381 = N2345 | N2380;
  assign N2382 = ~N2381;
  assign N2383 = waddr_i[5] | N2380;
  assign N2384 = ~N2383;
  assign N2385 = N2337 | waddr_i[9];
  assign N2386 = N2338 | N2385;
  assign N2387 = N2339 | N2386;
  assign N2388 = N2345 | N2387;
  assign N2389 = ~N2388;
  assign N2390 = waddr_i[5] | N2387;
  assign N2391 = ~N2390;
  assign N2392 = waddr_i[6] | N2386;
  assign N2393 = N2345 | N2392;
  assign N2394 = ~N2393;
  assign N2395 = waddr_i[5] | N2392;
  assign N2396 = ~N2395;
  assign N2397 = waddr_i[7] | N2385;
  assign N2398 = N2339 | N2397;
  assign N2399 = N2345 | N2398;
  assign N2400 = ~N2399;
  assign N2401 = waddr_i[5] | N2398;
  assign N2402 = ~N2401;
  assign N2403 = waddr_i[6] | N2397;
  assign N2404 = N2345 | N2403;
  assign N2405 = ~N2404;
  assign N2406 = waddr_i[5] | N2403;
  assign N2407 = ~N2406;
  assign N2408 = waddr_i[8] | waddr_i[9];
  assign N2409 = N2338 | N2408;
  assign N2410 = N2339 | N2409;
  assign N2411 = N2345 | N2410;
  assign N2412 = ~N2411;
  assign N2413 = waddr_i[5] | N2410;
  assign N2414 = ~N2413;
  assign N2415 = waddr_i[6] | N2409;
  assign N2416 = N2345 | N2415;
  assign N2417 = ~N2416;
  assign N2418 = waddr_i[5] | N2415;
  assign N2419 = ~N2418;
  assign N2420 = waddr_i[7] | N2408;
  assign N2421 = N2339 | N2420;
  assign N2422 = N2345 | N2421;
  assign N2423 = ~N2422;
  assign N2424 = waddr_i[5] | N2421;
  assign N2425 = ~N2424;
  assign N2426 = waddr_i[6] | N2420;
  assign N2427 = N2345 | N2426;
  assign N2428 = ~N2427;
  assign N2429 = waddr_i[3] & waddr_i[4];
  assign N2430 = waddr_i[2] & N2429;
  assign N2431 = waddr_i[1] & N2430;
  assign N2432 = waddr_i[0] & N2431;
  assign N2433 = ~waddr_i[4];
  assign N2434 = ~waddr_i[3];
  assign N2435 = ~waddr_i[2];
  assign N2436 = ~waddr_i[1];
  assign N2437 = N2434 | N2433;
  assign N2438 = N2435 | N2437;
  assign N2439 = N2436 | N2438;
  assign N2440 = waddr_i[0] | N2439;
  assign N2441 = ~N2440;
  assign N2442 = ~waddr_i[0];
  assign N2443 = waddr_i[1] | N2438;
  assign N2444 = N2442 | N2443;
  assign N2445 = ~N2444;
  assign N2446 = waddr_i[0] | N2443;
  assign N2447 = ~N2446;
  assign N2448 = waddr_i[2] | N2437;
  assign N2449 = N2436 | N2448;
  assign N2450 = N2442 | N2449;
  assign N2451 = ~N2450;
  assign N2452 = waddr_i[0] | N2449;
  assign N2453 = ~N2452;
  assign N2454 = waddr_i[1] | N2448;
  assign N2455 = N2442 | N2454;
  assign N2456 = ~N2455;
  assign N2457 = waddr_i[0] | N2454;
  assign N2458 = ~N2457;
  assign N2459 = waddr_i[3] | N2433;
  assign N2460 = N2435 | N2459;
  assign N2461 = N2436 | N2460;
  assign N2462 = N2442 | N2461;
  assign N2463 = ~N2462;
  assign N2464 = waddr_i[0] | N2461;
  assign N2465 = ~N2464;
  assign N2466 = waddr_i[1] | N2460;
  assign N2467 = N2442 | N2466;
  assign N2468 = ~N2467;
  assign N2469 = waddr_i[0] | N2466;
  assign N2470 = ~N2469;
  assign N2471 = waddr_i[2] | N2459;
  assign N2472 = N2436 | N2471;
  assign N2473 = N2442 | N2472;
  assign N2474 = ~N2473;
  assign N2475 = waddr_i[0] | N2472;
  assign N2476 = ~N2475;
  assign N2477 = waddr_i[1] | N2471;
  assign N2478 = N2442 | N2477;
  assign N2479 = ~N2478;
  assign N2480 = waddr_i[0] | N2477;
  assign N2481 = ~N2480;
  assign N2482 = N2434 | waddr_i[4];
  assign N2483 = N2435 | N2482;
  assign N2484 = N2436 | N2483;
  assign N2485 = N2442 | N2484;
  assign N2486 = ~N2485;
  assign N2487 = waddr_i[0] | N2484;
  assign N2488 = ~N2487;
  assign N2489 = waddr_i[1] | N2483;
  assign N2490 = N2442 | N2489;
  assign N2491 = ~N2490;
  assign N2492 = waddr_i[0] | N2489;
  assign N2493 = ~N2492;
  assign N2494 = waddr_i[2] | N2482;
  assign N2495 = N2436 | N2494;
  assign N2496 = N2442 | N2495;
  assign N2497 = ~N2496;
  assign N2498 = waddr_i[0] | N2495;
  assign N2499 = ~N2498;
  assign N2500 = waddr_i[1] | N2494;
  assign N2501 = N2442 | N2500;
  assign N2502 = ~N2501;
  assign N2503 = waddr_i[0] | N2500;
  assign N2504 = ~N2503;
  assign N2505 = waddr_i[3] | waddr_i[4];
  assign N2506 = N2435 | N2505;
  assign N2507 = N2436 | N2506;
  assign N2508 = N2442 | N2507;
  assign N2509 = ~N2508;
  assign N2510 = waddr_i[0] | N2507;
  assign N2511 = ~N2510;
  assign N2512 = waddr_i[1] | N2506;
  assign N2513 = N2442 | N2512;
  assign N2514 = ~N2513;
  assign N2515 = waddr_i[0] | N2512;
  assign N2516 = ~N2515;
  assign N2517 = waddr_i[2] | N2505;
  assign N2518 = N2436 | N2517;
  assign N2519 = N2442 | N2518;
  assign N2520 = ~N2519;
  assign N2521 = waddr_i[0] | N2518;
  assign N2522 = ~N2521;
  assign N2523 = waddr_i[1] | N2517;
  assign N2524 = N2442 | N2523;
  assign N2525 = ~N2524;
  assign we_dec_0__1_ = (N0)? we_i[0] : 
                        (N1)? 1'b0 : 1'b0;
  assign N0 = N2525;
  assign N1 = N2524;
  assign we_dec_0__2_ = (N2)? we_i[0] : 
                        (N3)? 1'b0 : 1'b0;
  assign N2 = N2522;
  assign N3 = N2521;
  assign we_dec_0__3_ = (N4)? we_i[0] : 
                        (N5)? 1'b0 : 1'b0;
  assign N4 = N2520;
  assign N5 = N2519;
  assign we_dec_0__4_ = (N6)? we_i[0] : 
                        (N7)? 1'b0 : 1'b0;
  assign N6 = N2516;
  assign N7 = N2515;
  assign we_dec_0__5_ = (N8)? we_i[0] : 
                        (N9)? 1'b0 : 1'b0;
  assign N8 = N2514;
  assign N9 = N2513;
  assign we_dec_0__6_ = (N10)? we_i[0] : 
                        (N11)? 1'b0 : 1'b0;
  assign N10 = N2511;
  assign N11 = N2510;
  assign we_dec_0__7_ = (N12)? we_i[0] : 
                        (N13)? 1'b0 : 1'b0;
  assign N12 = N2509;
  assign N13 = N2508;
  assign we_dec_0__8_ = (N14)? we_i[0] : 
                        (N15)? 1'b0 : 1'b0;
  assign N14 = N2504;
  assign N15 = N2503;
  assign we_dec_0__9_ = (N16)? we_i[0] : 
                        (N17)? 1'b0 : 1'b0;
  assign N16 = N2502;
  assign N17 = N2501;
  assign we_dec_0__10_ = (N18)? we_i[0] : 
                         (N19)? 1'b0 : 1'b0;
  assign N18 = N2499;
  assign N19 = N2498;
  assign we_dec_0__11_ = (N20)? we_i[0] : 
                         (N21)? 1'b0 : 1'b0;
  assign N20 = N2497;
  assign N21 = N2496;
  assign we_dec_0__12_ = (N22)? we_i[0] : 
                         (N23)? 1'b0 : 1'b0;
  assign N22 = N2493;
  assign N23 = N2492;
  assign we_dec_0__13_ = (N24)? we_i[0] : 
                         (N25)? 1'b0 : 1'b0;
  assign N24 = N2491;
  assign N25 = N2490;
  assign we_dec_0__14_ = (N26)? we_i[0] : 
                         (N27)? 1'b0 : 1'b0;
  assign N26 = N2488;
  assign N27 = N2487;
  assign we_dec_0__15_ = (N28)? we_i[0] : 
                         (N29)? 1'b0 : 1'b0;
  assign N28 = N2486;
  assign N29 = N2485;
  assign we_dec_0__16_ = (N30)? we_i[0] : 
                         (N31)? 1'b0 : 1'b0;
  assign N30 = N2481;
  assign N31 = N2480;
  assign we_dec_0__17_ = (N32)? we_i[0] : 
                         (N33)? 1'b0 : 1'b0;
  assign N32 = N2479;
  assign N33 = N2478;
  assign we_dec_0__18_ = (N34)? we_i[0] : 
                         (N35)? 1'b0 : 1'b0;
  assign N34 = N2476;
  assign N35 = N2475;
  assign we_dec_0__19_ = (N36)? we_i[0] : 
                         (N37)? 1'b0 : 1'b0;
  assign N36 = N2474;
  assign N37 = N2473;
  assign we_dec_0__20_ = (N38)? we_i[0] : 
                         (N39)? 1'b0 : 1'b0;
  assign N38 = N2470;
  assign N39 = N2469;
  assign we_dec_0__21_ = (N40)? we_i[0] : 
                         (N41)? 1'b0 : 1'b0;
  assign N40 = N2468;
  assign N41 = N2467;
  assign we_dec_0__22_ = (N42)? we_i[0] : 
                         (N43)? 1'b0 : 1'b0;
  assign N42 = N2465;
  assign N43 = N2464;
  assign we_dec_0__23_ = (N44)? we_i[0] : 
                         (N45)? 1'b0 : 1'b0;
  assign N44 = N2463;
  assign N45 = N2462;
  assign we_dec_0__24_ = (N46)? we_i[0] : 
                         (N47)? 1'b0 : 1'b0;
  assign N46 = N2458;
  assign N47 = N2457;
  assign we_dec_0__25_ = (N48)? we_i[0] : 
                         (N49)? 1'b0 : 1'b0;
  assign N48 = N2456;
  assign N49 = N2455;
  assign we_dec_0__26_ = (N50)? we_i[0] : 
                         (N51)? 1'b0 : 1'b0;
  assign N50 = N2453;
  assign N51 = N2452;
  assign we_dec_0__27_ = (N52)? we_i[0] : 
                         (N53)? 1'b0 : 1'b0;
  assign N52 = N2451;
  assign N53 = N2450;
  assign we_dec_0__28_ = (N54)? we_i[0] : 
                         (N55)? 1'b0 : 1'b0;
  assign N54 = N2447;
  assign N55 = N2446;
  assign we_dec_0__29_ = (N56)? we_i[0] : 
                         (N57)? 1'b0 : 1'b0;
  assign N56 = N2445;
  assign N57 = N2444;
  assign we_dec_0__30_ = (N58)? we_i[0] : 
                         (N59)? 1'b0 : 1'b0;
  assign N58 = N2441;
  assign N59 = N2440;
  assign we_dec_0__31_ = (N60)? we_i[0] : 
                         (N153)? 1'b0 : 1'b0;
  assign N60 = N2432;
  assign we_dec_1__1_ = (N61)? we_i[1] : 
                        (N62)? 1'b0 : 1'b0;
  assign N61 = N2428;
  assign N62 = N2427;
  assign we_dec_1__2_ = (N63)? we_i[1] : 
                        (N64)? 1'b0 : 1'b0;
  assign N63 = N2425;
  assign N64 = N2424;
  assign we_dec_1__3_ = (N65)? we_i[1] : 
                        (N66)? 1'b0 : 1'b0;
  assign N65 = N2423;
  assign N66 = N2422;
  assign we_dec_1__4_ = (N67)? we_i[1] : 
                        (N68)? 1'b0 : 1'b0;
  assign N67 = N2419;
  assign N68 = N2418;
  assign we_dec_1__5_ = (N69)? we_i[1] : 
                        (N70)? 1'b0 : 1'b0;
  assign N69 = N2417;
  assign N70 = N2416;
  assign we_dec_1__6_ = (N71)? we_i[1] : 
                        (N72)? 1'b0 : 1'b0;
  assign N71 = N2414;
  assign N72 = N2413;
  assign we_dec_1__7_ = (N73)? we_i[1] : 
                        (N74)? 1'b0 : 1'b0;
  assign N73 = N2412;
  assign N74 = N2411;
  assign we_dec_1__8_ = (N75)? we_i[1] : 
                        (N76)? 1'b0 : 1'b0;
  assign N75 = N2407;
  assign N76 = N2406;
  assign we_dec_1__9_ = (N77)? we_i[1] : 
                        (N78)? 1'b0 : 1'b0;
  assign N77 = N2405;
  assign N78 = N2404;
  assign we_dec_1__10_ = (N79)? we_i[1] : 
                         (N80)? 1'b0 : 1'b0;
  assign N79 = N2402;
  assign N80 = N2401;
  assign we_dec_1__11_ = (N81)? we_i[1] : 
                         (N82)? 1'b0 : 1'b0;
  assign N81 = N2400;
  assign N82 = N2399;
  assign we_dec_1__12_ = (N83)? we_i[1] : 
                         (N84)? 1'b0 : 1'b0;
  assign N83 = N2396;
  assign N84 = N2395;
  assign we_dec_1__13_ = (N85)? we_i[1] : 
                         (N86)? 1'b0 : 1'b0;
  assign N85 = N2394;
  assign N86 = N2393;
  assign we_dec_1__14_ = (N87)? we_i[1] : 
                         (N88)? 1'b0 : 1'b0;
  assign N87 = N2391;
  assign N88 = N2390;
  assign we_dec_1__15_ = (N89)? we_i[1] : 
                         (N90)? 1'b0 : 1'b0;
  assign N89 = N2389;
  assign N90 = N2388;
  assign we_dec_1__16_ = (N91)? we_i[1] : 
                         (N92)? 1'b0 : 1'b0;
  assign N91 = N2384;
  assign N92 = N2383;
  assign we_dec_1__17_ = (N93)? we_i[1] : 
                         (N94)? 1'b0 : 1'b0;
  assign N93 = N2382;
  assign N94 = N2381;
  assign we_dec_1__18_ = (N95)? we_i[1] : 
                         (N96)? 1'b0 : 1'b0;
  assign N95 = N2379;
  assign N96 = N2378;
  assign we_dec_1__19_ = (N97)? we_i[1] : 
                         (N98)? 1'b0 : 1'b0;
  assign N97 = N2377;
  assign N98 = N2376;
  assign we_dec_1__20_ = (N99)? we_i[1] : 
                         (N100)? 1'b0 : 1'b0;
  assign N99 = N2373;
  assign N100 = N2372;
  assign we_dec_1__21_ = (N101)? we_i[1] : 
                         (N102)? 1'b0 : 1'b0;
  assign N101 = N2371;
  assign N102 = N2370;
  assign we_dec_1__22_ = (N103)? we_i[1] : 
                         (N104)? 1'b0 : 1'b0;
  assign N103 = N2368;
  assign N104 = N2367;
  assign we_dec_1__23_ = (N105)? we_i[1] : 
                         (N106)? 1'b0 : 1'b0;
  assign N105 = N2366;
  assign N106 = N2365;
  assign we_dec_1__24_ = (N107)? we_i[1] : 
                         (N108)? 1'b0 : 1'b0;
  assign N107 = N2361;
  assign N108 = N2360;
  assign we_dec_1__25_ = (N109)? we_i[1] : 
                         (N110)? 1'b0 : 1'b0;
  assign N109 = N2359;
  assign N110 = N2358;
  assign we_dec_1__26_ = (N111)? we_i[1] : 
                         (N112)? 1'b0 : 1'b0;
  assign N111 = N2356;
  assign N112 = N2355;
  assign we_dec_1__27_ = (N113)? we_i[1] : 
                         (N114)? 1'b0 : 1'b0;
  assign N113 = N2354;
  assign N114 = N2353;
  assign we_dec_1__28_ = (N115)? we_i[1] : 
                         (N116)? 1'b0 : 1'b0;
  assign N115 = N2350;
  assign N116 = N2349;
  assign we_dec_1__29_ = (N117)? we_i[1] : 
                         (N118)? 1'b0 : 1'b0;
  assign N117 = N2348;
  assign N118 = N2347;
  assign we_dec_1__30_ = (N119)? we_i[1] : 
                         (N120)? 1'b0 : 1'b0;
  assign N119 = N2344;
  assign N120 = N2343;
  assign we_dec_1__31_ = (N121)? we_i[1] : 
                         (N154)? 1'b0 : 1'b0;
  assign N121 = N2335;
  assign N157 = (N122)? 1'b1 : 
                (N156)? we_dec_0__1_ : 1'b0;
  assign N122 = we_dec_1__1_;
  assign { N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158 } = (N122)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N156)? wdata_i[63:0] : 1'b0;
  assign N223 = (N123)? 1'b1 : 
                (N222)? we_dec_0__2_ : 1'b0;
  assign N123 = we_dec_1__2_;
  assign { N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224 } = (N123)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N222)? wdata_i[63:0] : 1'b0;
  assign N289 = (N124)? 1'b1 : 
                (N288)? we_dec_0__3_ : 1'b0;
  assign N124 = we_dec_1__3_;
  assign { N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290 } = (N124)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N288)? wdata_i[63:0] : 1'b0;
  assign N355 = (N125)? 1'b1 : 
                (N354)? we_dec_0__4_ : 1'b0;
  assign N125 = we_dec_1__4_;
  assign { N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356 } = (N125)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N354)? wdata_i[63:0] : 1'b0;
  assign N421 = (N126)? 1'b1 : 
                (N420)? we_dec_0__5_ : 1'b0;
  assign N126 = we_dec_1__5_;
  assign { N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422 } = (N126)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N420)? wdata_i[63:0] : 1'b0;
  assign N487 = (N127)? 1'b1 : 
                (N486)? we_dec_0__6_ : 1'b0;
  assign N127 = we_dec_1__6_;
  assign { N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488 } = (N127)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N486)? wdata_i[63:0] : 1'b0;
  assign N553 = (N128)? 1'b1 : 
                (N552)? we_dec_0__7_ : 1'b0;
  assign N128 = we_dec_1__7_;
  assign { N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554 } = (N128)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N552)? wdata_i[63:0] : 1'b0;
  assign N619 = (N129)? 1'b1 : 
                (N618)? we_dec_0__8_ : 1'b0;
  assign N129 = we_dec_1__8_;
  assign { N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620 } = (N129)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N618)? wdata_i[63:0] : 1'b0;
  assign N685 = (N130)? 1'b1 : 
                (N684)? we_dec_0__9_ : 1'b0;
  assign N130 = we_dec_1__9_;
  assign { N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686 } = (N130)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N684)? wdata_i[63:0] : 1'b0;
  assign N751 = (N131)? 1'b1 : 
                (N750)? we_dec_0__10_ : 1'b0;
  assign N131 = we_dec_1__10_;
  assign { N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752 } = (N131)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N750)? wdata_i[63:0] : 1'b0;
  assign N817 = (N132)? 1'b1 : 
                (N816)? we_dec_0__11_ : 1'b0;
  assign N132 = we_dec_1__11_;
  assign { N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818 } = (N132)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N816)? wdata_i[63:0] : 1'b0;
  assign N883 = (N133)? 1'b1 : 
                (N882)? we_dec_0__12_ : 1'b0;
  assign N133 = we_dec_1__12_;
  assign { N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884 } = (N133)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N882)? wdata_i[63:0] : 1'b0;
  assign N949 = (N134)? 1'b1 : 
                (N948)? we_dec_0__13_ : 1'b0;
  assign N134 = we_dec_1__13_;
  assign { N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950 } = (N134)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                            (N948)? wdata_i[63:0] : 1'b0;
  assign N1015 = (N135)? 1'b1 : 
                 (N1014)? we_dec_0__14_ : 1'b0;
  assign N135 = we_dec_1__14_;
  assign { N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016 } = (N135)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1014)? wdata_i[63:0] : 1'b0;
  assign N1081 = (N136)? 1'b1 : 
                 (N1080)? we_dec_0__15_ : 1'b0;
  assign N136 = we_dec_1__15_;
  assign { N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082 } = (N136)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1080)? wdata_i[63:0] : 1'b0;
  assign N1147 = (N137)? 1'b1 : 
                 (N1146)? we_dec_0__16_ : 1'b0;
  assign N137 = we_dec_1__16_;
  assign { N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148 } = (N137)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1146)? wdata_i[63:0] : 1'b0;
  assign N1213 = (N138)? 1'b1 : 
                 (N1212)? we_dec_0__17_ : 1'b0;
  assign N138 = we_dec_1__17_;
  assign { N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214 } = (N138)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1212)? wdata_i[63:0] : 1'b0;
  assign N1279 = (N139)? 1'b1 : 
                 (N1278)? we_dec_0__18_ : 1'b0;
  assign N139 = we_dec_1__18_;
  assign { N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280 } = (N139)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1278)? wdata_i[63:0] : 1'b0;
  assign N1345 = (N140)? 1'b1 : 
                 (N1344)? we_dec_0__19_ : 1'b0;
  assign N140 = we_dec_1__19_;
  assign { N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346 } = (N140)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1344)? wdata_i[63:0] : 1'b0;
  assign N1411 = (N141)? 1'b1 : 
                 (N1410)? we_dec_0__20_ : 1'b0;
  assign N141 = we_dec_1__20_;
  assign { N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412 } = (N141)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1410)? wdata_i[63:0] : 1'b0;
  assign N1477 = (N142)? 1'b1 : 
                 (N1476)? we_dec_0__21_ : 1'b0;
  assign N142 = we_dec_1__21_;
  assign { N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478 } = (N142)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1476)? wdata_i[63:0] : 1'b0;
  assign N1543 = (N143)? 1'b1 : 
                 (N1542)? we_dec_0__22_ : 1'b0;
  assign N143 = we_dec_1__22_;
  assign { N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544 } = (N143)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1542)? wdata_i[63:0] : 1'b0;
  assign N1609 = (N144)? 1'b1 : 
                 (N1608)? we_dec_0__23_ : 1'b0;
  assign N144 = we_dec_1__23_;
  assign { N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610 } = (N144)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1608)? wdata_i[63:0] : 1'b0;
  assign N1675 = (N145)? 1'b1 : 
                 (N1674)? we_dec_0__24_ : 1'b0;
  assign N145 = we_dec_1__24_;
  assign { N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676 } = (N145)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1674)? wdata_i[63:0] : 1'b0;
  assign N1741 = (N146)? 1'b1 : 
                 (N1740)? we_dec_0__25_ : 1'b0;
  assign N146 = we_dec_1__25_;
  assign { N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742 } = (N146)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1740)? wdata_i[63:0] : 1'b0;
  assign N1807 = (N147)? 1'b1 : 
                 (N1806)? we_dec_0__26_ : 1'b0;
  assign N147 = we_dec_1__26_;
  assign { N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808 } = (N147)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1806)? wdata_i[63:0] : 1'b0;
  assign N1873 = (N148)? 1'b1 : 
                 (N1872)? we_dec_0__27_ : 1'b0;
  assign N148 = we_dec_1__27_;
  assign { N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874 } = (N148)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1872)? wdata_i[63:0] : 1'b0;
  assign N1939 = (N149)? 1'b1 : 
                 (N1938)? we_dec_0__28_ : 1'b0;
  assign N149 = we_dec_1__28_;
  assign { N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940 } = (N149)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1938)? wdata_i[63:0] : 1'b0;
  assign N2005 = (N150)? 1'b1 : 
                 (N2004)? we_dec_0__29_ : 1'b0;
  assign N150 = we_dec_1__29_;
  assign { N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006 } = (N150)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2004)? wdata_i[63:0] : 1'b0;
  assign N2071 = (N151)? 1'b1 : 
                 (N2070)? we_dec_0__30_ : 1'b0;
  assign N151 = we_dec_1__30_;
  assign { N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072 } = (N151)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2070)? wdata_i[63:0] : 1'b0;
  assign N2137 = (N152)? 1'b1 : 
                 (N2136)? we_dec_0__31_ : 1'b0;
  assign N152 = we_dec_1__31_;
  assign { N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138 } = (N152)? wdata_i[127:64] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N2136)? wdata_i[63:0] : 1'b0;
  assign N153 = ~N2432;
  assign N154 = ~N2335;
  assign N155 = ~rst_ni;
  assign N156 = ~we_dec_1__1_;
  assign N222 = ~we_dec_1__2_;
  assign N288 = ~we_dec_1__3_;
  assign N354 = ~we_dec_1__4_;
  assign N420 = ~we_dec_1__5_;
  assign N486 = ~we_dec_1__6_;
  assign N552 = ~we_dec_1__7_;
  assign N618 = ~we_dec_1__8_;
  assign N684 = ~we_dec_1__9_;
  assign N750 = ~we_dec_1__10_;
  assign N816 = ~we_dec_1__11_;
  assign N882 = ~we_dec_1__12_;
  assign N948 = ~we_dec_1__13_;
  assign N1014 = ~we_dec_1__14_;
  assign N1080 = ~we_dec_1__15_;
  assign N1146 = ~we_dec_1__16_;
  assign N1212 = ~we_dec_1__17_;
  assign N1278 = ~we_dec_1__18_;
  assign N1344 = ~we_dec_1__19_;
  assign N1410 = ~we_dec_1__20_;
  assign N1476 = ~we_dec_1__21_;
  assign N1542 = ~we_dec_1__22_;
  assign N1608 = ~we_dec_1__23_;
  assign N1674 = ~we_dec_1__24_;
  assign N1740 = ~we_dec_1__25_;
  assign N1806 = ~we_dec_1__26_;
  assign N1872 = ~we_dec_1__27_;
  assign N1938 = ~we_dec_1__28_;
  assign N2004 = ~we_dec_1__29_;
  assign N2070 = ~we_dec_1__30_;
  assign N2136 = ~we_dec_1__31_;
  assign N2202 = ~raddr_i[0];
  assign N2203 = ~raddr_i[1];
  assign N2204 = N2202 & N2203;
  assign N2205 = N2202 & raddr_i[1];
  assign N2206 = raddr_i[0] & N2203;
  assign N2207 = raddr_i[0] & raddr_i[1];
  assign N2208 = ~raddr_i[2];
  assign N2209 = N2204 & N2208;
  assign N2210 = N2204 & raddr_i[2];
  assign N2211 = N2206 & N2208;
  assign N2212 = N2206 & raddr_i[2];
  assign N2213 = N2205 & N2208;
  assign N2214 = N2205 & raddr_i[2];
  assign N2215 = N2207 & N2208;
  assign N2216 = N2207 & raddr_i[2];
  assign N2217 = ~raddr_i[3];
  assign N2218 = N2209 & N2217;
  assign N2219 = N2209 & raddr_i[3];
  assign N2220 = N2211 & N2217;
  assign N2221 = N2211 & raddr_i[3];
  assign N2222 = N2213 & N2217;
  assign N2223 = N2213 & raddr_i[3];
  assign N2224 = N2215 & N2217;
  assign N2225 = N2215 & raddr_i[3];
  assign N2226 = N2210 & N2217;
  assign N2227 = N2210 & raddr_i[3];
  assign N2228 = N2212 & N2217;
  assign N2229 = N2212 & raddr_i[3];
  assign N2230 = N2214 & N2217;
  assign N2231 = N2214 & raddr_i[3];
  assign N2232 = N2216 & N2217;
  assign N2233 = N2216 & raddr_i[3];
  assign N2234 = ~raddr_i[4];
  assign N2235 = N2218 & N2234;
  assign N2236 = N2218 & raddr_i[4];
  assign N2237 = N2220 & N2234;
  assign N2238 = N2220 & raddr_i[4];
  assign N2239 = N2222 & N2234;
  assign N2240 = N2222 & raddr_i[4];
  assign N2241 = N2224 & N2234;
  assign N2242 = N2224 & raddr_i[4];
  assign N2243 = N2226 & N2234;
  assign N2244 = N2226 & raddr_i[4];
  assign N2245 = N2228 & N2234;
  assign N2246 = N2228 & raddr_i[4];
  assign N2247 = N2230 & N2234;
  assign N2248 = N2230 & raddr_i[4];
  assign N2249 = N2232 & N2234;
  assign N2250 = N2232 & raddr_i[4];
  assign N2251 = N2219 & N2234;
  assign N2252 = N2219 & raddr_i[4];
  assign N2253 = N2221 & N2234;
  assign N2254 = N2221 & raddr_i[4];
  assign N2255 = N2223 & N2234;
  assign N2256 = N2223 & raddr_i[4];
  assign N2257 = N2225 & N2234;
  assign N2258 = N2225 & raddr_i[4];
  assign N2259 = N2227 & N2234;
  assign N2260 = N2227 & raddr_i[4];
  assign N2261 = N2229 & N2234;
  assign N2262 = N2229 & raddr_i[4];
  assign N2263 = N2231 & N2234;
  assign N2264 = N2231 & raddr_i[4];
  assign N2265 = N2233 & N2234;
  assign N2266 = N2233 & raddr_i[4];
  assign N2267 = ~raddr_i[5];
  assign N2268 = ~raddr_i[6];
  assign N2269 = N2267 & N2268;
  assign N2270 = N2267 & raddr_i[6];
  assign N2271 = raddr_i[5] & N2268;
  assign N2272 = raddr_i[5] & raddr_i[6];
  assign N2273 = ~raddr_i[7];
  assign N2274 = N2269 & N2273;
  assign N2275 = N2269 & raddr_i[7];
  assign N2276 = N2271 & N2273;
  assign N2277 = N2271 & raddr_i[7];
  assign N2278 = N2270 & N2273;
  assign N2279 = N2270 & raddr_i[7];
  assign N2280 = N2272 & N2273;
  assign N2281 = N2272 & raddr_i[7];
  assign N2282 = ~raddr_i[8];
  assign N2283 = N2274 & N2282;
  assign N2284 = N2274 & raddr_i[8];
  assign N2285 = N2276 & N2282;
  assign N2286 = N2276 & raddr_i[8];
  assign N2287 = N2278 & N2282;
  assign N2288 = N2278 & raddr_i[8];
  assign N2289 = N2280 & N2282;
  assign N2290 = N2280 & raddr_i[8];
  assign N2291 = N2275 & N2282;
  assign N2292 = N2275 & raddr_i[8];
  assign N2293 = N2277 & N2282;
  assign N2294 = N2277 & raddr_i[8];
  assign N2295 = N2279 & N2282;
  assign N2296 = N2279 & raddr_i[8];
  assign N2297 = N2281 & N2282;
  assign N2298 = N2281 & raddr_i[8];
  assign N2299 = ~raddr_i[9];
  assign N2300 = N2283 & N2299;
  assign N2301 = N2283 & raddr_i[9];
  assign N2302 = N2285 & N2299;
  assign N2303 = N2285 & raddr_i[9];
  assign N2304 = N2287 & N2299;
  assign N2305 = N2287 & raddr_i[9];
  assign N2306 = N2289 & N2299;
  assign N2307 = N2289 & raddr_i[9];
  assign N2308 = N2291 & N2299;
  assign N2309 = N2291 & raddr_i[9];
  assign N2310 = N2293 & N2299;
  assign N2311 = N2293 & raddr_i[9];
  assign N2312 = N2295 & N2299;
  assign N2313 = N2295 & raddr_i[9];
  assign N2314 = N2297 & N2299;
  assign N2315 = N2297 & raddr_i[9];
  assign N2316 = N2284 & N2299;
  assign N2317 = N2284 & raddr_i[9];
  assign N2318 = N2286 & N2299;
  assign N2319 = N2286 & raddr_i[9];
  assign N2320 = N2288 & N2299;
  assign N2321 = N2288 & raddr_i[9];
  assign N2322 = N2290 & N2299;
  assign N2323 = N2290 & raddr_i[9];
  assign N2324 = N2292 & N2299;
  assign N2325 = N2292 & raddr_i[9];
  assign N2326 = N2294 & N2299;
  assign N2327 = N2294 & raddr_i[9];
  assign N2328 = N2296 & N2299;
  assign N2329 = N2296 & raddr_i[9];
  assign N2330 = N2298 & N2299;
  assign N2331 = N2298 & raddr_i[9];

endmodule