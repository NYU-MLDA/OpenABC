module bsg_mem_2r1w_sync_synth_width_p64_els_p32_read_write_same_addr_p1_harden_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r0_v_i,
  r0_addr_i,
  r0_data_o,
  r1_v_i,
  r1_addr_i,
  r1_data_o
);

  input [4:0] w_addr_i;
  input [63:0] w_data_i;
  input [4:0] r0_addr_i;
  output [63:0] r0_data_o;
  input [4:0] r1_addr_i;
  output [63:0] r1_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r0_v_i;
  input r1_v_i;
  wire [63:0] r0_data_o,r1_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221;
  reg [4:0] r0_addr_r,r1_addr_r;
  reg [2047:0] mem;
  assign r0_data_o[63] = (N43)? mem[63] : 
                         (N45)? mem[127] : 
                         (N47)? mem[191] : 
                         (N49)? mem[255] : 
                         (N51)? mem[319] : 
                         (N53)? mem[383] : 
                         (N55)? mem[447] : 
                         (N57)? mem[511] : 
                         (N59)? mem[575] : 
                         (N61)? mem[639] : 
                         (N63)? mem[703] : 
                         (N65)? mem[767] : 
                         (N67)? mem[831] : 
                         (N69)? mem[895] : 
                         (N71)? mem[959] : 
                         (N73)? mem[1023] : 
                         (N44)? mem[1087] : 
                         (N46)? mem[1151] : 
                         (N48)? mem[1215] : 
                         (N50)? mem[1279] : 
                         (N52)? mem[1343] : 
                         (N54)? mem[1407] : 
                         (N56)? mem[1471] : 
                         (N58)? mem[1535] : 
                         (N60)? mem[1599] : 
                         (N62)? mem[1663] : 
                         (N64)? mem[1727] : 
                         (N66)? mem[1791] : 
                         (N68)? mem[1855] : 
                         (N70)? mem[1919] : 
                         (N72)? mem[1983] : 
                         (N74)? mem[2047] : 1'b0;
  assign r0_data_o[62] = (N43)? mem[62] : 
                         (N45)? mem[126] : 
                         (N47)? mem[190] : 
                         (N49)? mem[254] : 
                         (N51)? mem[318] : 
                         (N53)? mem[382] : 
                         (N55)? mem[446] : 
                         (N57)? mem[510] : 
                         (N59)? mem[574] : 
                         (N61)? mem[638] : 
                         (N63)? mem[702] : 
                         (N65)? mem[766] : 
                         (N67)? mem[830] : 
                         (N69)? mem[894] : 
                         (N71)? mem[958] : 
                         (N73)? mem[1022] : 
                         (N44)? mem[1086] : 
                         (N46)? mem[1150] : 
                         (N48)? mem[1214] : 
                         (N50)? mem[1278] : 
                         (N52)? mem[1342] : 
                         (N54)? mem[1406] : 
                         (N56)? mem[1470] : 
                         (N58)? mem[1534] : 
                         (N60)? mem[1598] : 
                         (N62)? mem[1662] : 
                         (N64)? mem[1726] : 
                         (N66)? mem[1790] : 
                         (N68)? mem[1854] : 
                         (N70)? mem[1918] : 
                         (N72)? mem[1982] : 
                         (N74)? mem[2046] : 1'b0;
  assign r0_data_o[61] = (N43)? mem[61] : 
                         (N45)? mem[125] : 
                         (N47)? mem[189] : 
                         (N49)? mem[253] : 
                         (N51)? mem[317] : 
                         (N53)? mem[381] : 
                         (N55)? mem[445] : 
                         (N57)? mem[509] : 
                         (N59)? mem[573] : 
                         (N61)? mem[637] : 
                         (N63)? mem[701] : 
                         (N65)? mem[765] : 
                         (N67)? mem[829] : 
                         (N69)? mem[893] : 
                         (N71)? mem[957] : 
                         (N73)? mem[1021] : 
                         (N44)? mem[1085] : 
                         (N46)? mem[1149] : 
                         (N48)? mem[1213] : 
                         (N50)? mem[1277] : 
                         (N52)? mem[1341] : 
                         (N54)? mem[1405] : 
                         (N56)? mem[1469] : 
                         (N58)? mem[1533] : 
                         (N60)? mem[1597] : 
                         (N62)? mem[1661] : 
                         (N64)? mem[1725] : 
                         (N66)? mem[1789] : 
                         (N68)? mem[1853] : 
                         (N70)? mem[1917] : 
                         (N72)? mem[1981] : 
                         (N74)? mem[2045] : 1'b0;
  assign r0_data_o[60] = (N43)? mem[60] : 
                         (N45)? mem[124] : 
                         (N47)? mem[188] : 
                         (N49)? mem[252] : 
                         (N51)? mem[316] : 
                         (N53)? mem[380] : 
                         (N55)? mem[444] : 
                         (N57)? mem[508] : 
                         (N59)? mem[572] : 
                         (N61)? mem[636] : 
                         (N63)? mem[700] : 
                         (N65)? mem[764] : 
                         (N67)? mem[828] : 
                         (N69)? mem[892] : 
                         (N71)? mem[956] : 
                         (N73)? mem[1020] : 
                         (N44)? mem[1084] : 
                         (N46)? mem[1148] : 
                         (N48)? mem[1212] : 
                         (N50)? mem[1276] : 
                         (N52)? mem[1340] : 
                         (N54)? mem[1404] : 
                         (N56)? mem[1468] : 
                         (N58)? mem[1532] : 
                         (N60)? mem[1596] : 
                         (N62)? mem[1660] : 
                         (N64)? mem[1724] : 
                         (N66)? mem[1788] : 
                         (N68)? mem[1852] : 
                         (N70)? mem[1916] : 
                         (N72)? mem[1980] : 
                         (N74)? mem[2044] : 1'b0;
  assign r0_data_o[59] = (N43)? mem[59] : 
                         (N45)? mem[123] : 
                         (N47)? mem[187] : 
                         (N49)? mem[251] : 
                         (N51)? mem[315] : 
                         (N53)? mem[379] : 
                         (N55)? mem[443] : 
                         (N57)? mem[507] : 
                         (N59)? mem[571] : 
                         (N61)? mem[635] : 
                         (N63)? mem[699] : 
                         (N65)? mem[763] : 
                         (N67)? mem[827] : 
                         (N69)? mem[891] : 
                         (N71)? mem[955] : 
                         (N73)? mem[1019] : 
                         (N44)? mem[1083] : 
                         (N46)? mem[1147] : 
                         (N48)? mem[1211] : 
                         (N50)? mem[1275] : 
                         (N52)? mem[1339] : 
                         (N54)? mem[1403] : 
                         (N56)? mem[1467] : 
                         (N58)? mem[1531] : 
                         (N60)? mem[1595] : 
                         (N62)? mem[1659] : 
                         (N64)? mem[1723] : 
                         (N66)? mem[1787] : 
                         (N68)? mem[1851] : 
                         (N70)? mem[1915] : 
                         (N72)? mem[1979] : 
                         (N74)? mem[2043] : 1'b0;
  assign r0_data_o[58] = (N43)? mem[58] : 
                         (N45)? mem[122] : 
                         (N47)? mem[186] : 
                         (N49)? mem[250] : 
                         (N51)? mem[314] : 
                         (N53)? mem[378] : 
                         (N55)? mem[442] : 
                         (N57)? mem[506] : 
                         (N59)? mem[570] : 
                         (N61)? mem[634] : 
                         (N63)? mem[698] : 
                         (N65)? mem[762] : 
                         (N67)? mem[826] : 
                         (N69)? mem[890] : 
                         (N71)? mem[954] : 
                         (N73)? mem[1018] : 
                         (N44)? mem[1082] : 
                         (N46)? mem[1146] : 
                         (N48)? mem[1210] : 
                         (N50)? mem[1274] : 
                         (N52)? mem[1338] : 
                         (N54)? mem[1402] : 
                         (N56)? mem[1466] : 
                         (N58)? mem[1530] : 
                         (N60)? mem[1594] : 
                         (N62)? mem[1658] : 
                         (N64)? mem[1722] : 
                         (N66)? mem[1786] : 
                         (N68)? mem[1850] : 
                         (N70)? mem[1914] : 
                         (N72)? mem[1978] : 
                         (N74)? mem[2042] : 1'b0;
  assign r0_data_o[57] = (N43)? mem[57] : 
                         (N45)? mem[121] : 
                         (N47)? mem[185] : 
                         (N49)? mem[249] : 
                         (N51)? mem[313] : 
                         (N53)? mem[377] : 
                         (N55)? mem[441] : 
                         (N57)? mem[505] : 
                         (N59)? mem[569] : 
                         (N61)? mem[633] : 
                         (N63)? mem[697] : 
                         (N65)? mem[761] : 
                         (N67)? mem[825] : 
                         (N69)? mem[889] : 
                         (N71)? mem[953] : 
                         (N73)? mem[1017] : 
                         (N44)? mem[1081] : 
                         (N46)? mem[1145] : 
                         (N48)? mem[1209] : 
                         (N50)? mem[1273] : 
                         (N52)? mem[1337] : 
                         (N54)? mem[1401] : 
                         (N56)? mem[1465] : 
                         (N58)? mem[1529] : 
                         (N60)? mem[1593] : 
                         (N62)? mem[1657] : 
                         (N64)? mem[1721] : 
                         (N66)? mem[1785] : 
                         (N68)? mem[1849] : 
                         (N70)? mem[1913] : 
                         (N72)? mem[1977] : 
                         (N74)? mem[2041] : 1'b0;
  assign r0_data_o[56] = (N43)? mem[56] : 
                         (N45)? mem[120] : 
                         (N47)? mem[184] : 
                         (N49)? mem[248] : 
                         (N51)? mem[312] : 
                         (N53)? mem[376] : 
                         (N55)? mem[440] : 
                         (N57)? mem[504] : 
                         (N59)? mem[568] : 
                         (N61)? mem[632] : 
                         (N63)? mem[696] : 
                         (N65)? mem[760] : 
                         (N67)? mem[824] : 
                         (N69)? mem[888] : 
                         (N71)? mem[952] : 
                         (N73)? mem[1016] : 
                         (N44)? mem[1080] : 
                         (N46)? mem[1144] : 
                         (N48)? mem[1208] : 
                         (N50)? mem[1272] : 
                         (N52)? mem[1336] : 
                         (N54)? mem[1400] : 
                         (N56)? mem[1464] : 
                         (N58)? mem[1528] : 
                         (N60)? mem[1592] : 
                         (N62)? mem[1656] : 
                         (N64)? mem[1720] : 
                         (N66)? mem[1784] : 
                         (N68)? mem[1848] : 
                         (N70)? mem[1912] : 
                         (N72)? mem[1976] : 
                         (N74)? mem[2040] : 1'b0;
  assign r0_data_o[55] = (N43)? mem[55] : 
                         (N45)? mem[119] : 
                         (N47)? mem[183] : 
                         (N49)? mem[247] : 
                         (N51)? mem[311] : 
                         (N53)? mem[375] : 
                         (N55)? mem[439] : 
                         (N57)? mem[503] : 
                         (N59)? mem[567] : 
                         (N61)? mem[631] : 
                         (N63)? mem[695] : 
                         (N65)? mem[759] : 
                         (N67)? mem[823] : 
                         (N69)? mem[887] : 
                         (N71)? mem[951] : 
                         (N73)? mem[1015] : 
                         (N44)? mem[1079] : 
                         (N46)? mem[1143] : 
                         (N48)? mem[1207] : 
                         (N50)? mem[1271] : 
                         (N52)? mem[1335] : 
                         (N54)? mem[1399] : 
                         (N56)? mem[1463] : 
                         (N58)? mem[1527] : 
                         (N60)? mem[1591] : 
                         (N62)? mem[1655] : 
                         (N64)? mem[1719] : 
                         (N66)? mem[1783] : 
                         (N68)? mem[1847] : 
                         (N70)? mem[1911] : 
                         (N72)? mem[1975] : 
                         (N74)? mem[2039] : 1'b0;
  assign r0_data_o[54] = (N43)? mem[54] : 
                         (N45)? mem[118] : 
                         (N47)? mem[182] : 
                         (N49)? mem[246] : 
                         (N51)? mem[310] : 
                         (N53)? mem[374] : 
                         (N55)? mem[438] : 
                         (N57)? mem[502] : 
                         (N59)? mem[566] : 
                         (N61)? mem[630] : 
                         (N63)? mem[694] : 
                         (N65)? mem[758] : 
                         (N67)? mem[822] : 
                         (N69)? mem[886] : 
                         (N71)? mem[950] : 
                         (N73)? mem[1014] : 
                         (N44)? mem[1078] : 
                         (N46)? mem[1142] : 
                         (N48)? mem[1206] : 
                         (N50)? mem[1270] : 
                         (N52)? mem[1334] : 
                         (N54)? mem[1398] : 
                         (N56)? mem[1462] : 
                         (N58)? mem[1526] : 
                         (N60)? mem[1590] : 
                         (N62)? mem[1654] : 
                         (N64)? mem[1718] : 
                         (N66)? mem[1782] : 
                         (N68)? mem[1846] : 
                         (N70)? mem[1910] : 
                         (N72)? mem[1974] : 
                         (N74)? mem[2038] : 1'b0;
  assign r0_data_o[53] = (N43)? mem[53] : 
                         (N45)? mem[117] : 
                         (N47)? mem[181] : 
                         (N49)? mem[245] : 
                         (N51)? mem[309] : 
                         (N53)? mem[373] : 
                         (N55)? mem[437] : 
                         (N57)? mem[501] : 
                         (N59)? mem[565] : 
                         (N61)? mem[629] : 
                         (N63)? mem[693] : 
                         (N65)? mem[757] : 
                         (N67)? mem[821] : 
                         (N69)? mem[885] : 
                         (N71)? mem[949] : 
                         (N73)? mem[1013] : 
                         (N44)? mem[1077] : 
                         (N46)? mem[1141] : 
                         (N48)? mem[1205] : 
                         (N50)? mem[1269] : 
                         (N52)? mem[1333] : 
                         (N54)? mem[1397] : 
                         (N56)? mem[1461] : 
                         (N58)? mem[1525] : 
                         (N60)? mem[1589] : 
                         (N62)? mem[1653] : 
                         (N64)? mem[1717] : 
                         (N66)? mem[1781] : 
                         (N68)? mem[1845] : 
                         (N70)? mem[1909] : 
                         (N72)? mem[1973] : 
                         (N74)? mem[2037] : 1'b0;
  assign r0_data_o[52] = (N43)? mem[52] : 
                         (N45)? mem[116] : 
                         (N47)? mem[180] : 
                         (N49)? mem[244] : 
                         (N51)? mem[308] : 
                         (N53)? mem[372] : 
                         (N55)? mem[436] : 
                         (N57)? mem[500] : 
                         (N59)? mem[564] : 
                         (N61)? mem[628] : 
                         (N63)? mem[692] : 
                         (N65)? mem[756] : 
                         (N67)? mem[820] : 
                         (N69)? mem[884] : 
                         (N71)? mem[948] : 
                         (N73)? mem[1012] : 
                         (N44)? mem[1076] : 
                         (N46)? mem[1140] : 
                         (N48)? mem[1204] : 
                         (N50)? mem[1268] : 
                         (N52)? mem[1332] : 
                         (N54)? mem[1396] : 
                         (N56)? mem[1460] : 
                         (N58)? mem[1524] : 
                         (N60)? mem[1588] : 
                         (N62)? mem[1652] : 
                         (N64)? mem[1716] : 
                         (N66)? mem[1780] : 
                         (N68)? mem[1844] : 
                         (N70)? mem[1908] : 
                         (N72)? mem[1972] : 
                         (N74)? mem[2036] : 1'b0;
  assign r0_data_o[51] = (N43)? mem[51] : 
                         (N45)? mem[115] : 
                         (N47)? mem[179] : 
                         (N49)? mem[243] : 
                         (N51)? mem[307] : 
                         (N53)? mem[371] : 
                         (N55)? mem[435] : 
                         (N57)? mem[499] : 
                         (N59)? mem[563] : 
                         (N61)? mem[627] : 
                         (N63)? mem[691] : 
                         (N65)? mem[755] : 
                         (N67)? mem[819] : 
                         (N69)? mem[883] : 
                         (N71)? mem[947] : 
                         (N73)? mem[1011] : 
                         (N44)? mem[1075] : 
                         (N46)? mem[1139] : 
                         (N48)? mem[1203] : 
                         (N50)? mem[1267] : 
                         (N52)? mem[1331] : 
                         (N54)? mem[1395] : 
                         (N56)? mem[1459] : 
                         (N58)? mem[1523] : 
                         (N60)? mem[1587] : 
                         (N62)? mem[1651] : 
                         (N64)? mem[1715] : 
                         (N66)? mem[1779] : 
                         (N68)? mem[1843] : 
                         (N70)? mem[1907] : 
                         (N72)? mem[1971] : 
                         (N74)? mem[2035] : 1'b0;
  assign r0_data_o[50] = (N43)? mem[50] : 
                         (N45)? mem[114] : 
                         (N47)? mem[178] : 
                         (N49)? mem[242] : 
                         (N51)? mem[306] : 
                         (N53)? mem[370] : 
                         (N55)? mem[434] : 
                         (N57)? mem[498] : 
                         (N59)? mem[562] : 
                         (N61)? mem[626] : 
                         (N63)? mem[690] : 
                         (N65)? mem[754] : 
                         (N67)? mem[818] : 
                         (N69)? mem[882] : 
                         (N71)? mem[946] : 
                         (N73)? mem[1010] : 
                         (N44)? mem[1074] : 
                         (N46)? mem[1138] : 
                         (N48)? mem[1202] : 
                         (N50)? mem[1266] : 
                         (N52)? mem[1330] : 
                         (N54)? mem[1394] : 
                         (N56)? mem[1458] : 
                         (N58)? mem[1522] : 
                         (N60)? mem[1586] : 
                         (N62)? mem[1650] : 
                         (N64)? mem[1714] : 
                         (N66)? mem[1778] : 
                         (N68)? mem[1842] : 
                         (N70)? mem[1906] : 
                         (N72)? mem[1970] : 
                         (N74)? mem[2034] : 1'b0;
  assign r0_data_o[49] = (N43)? mem[49] : 
                         (N45)? mem[113] : 
                         (N47)? mem[177] : 
                         (N49)? mem[241] : 
                         (N51)? mem[305] : 
                         (N53)? mem[369] : 
                         (N55)? mem[433] : 
                         (N57)? mem[497] : 
                         (N59)? mem[561] : 
                         (N61)? mem[625] : 
                         (N63)? mem[689] : 
                         (N65)? mem[753] : 
                         (N67)? mem[817] : 
                         (N69)? mem[881] : 
                         (N71)? mem[945] : 
                         (N73)? mem[1009] : 
                         (N44)? mem[1073] : 
                         (N46)? mem[1137] : 
                         (N48)? mem[1201] : 
                         (N50)? mem[1265] : 
                         (N52)? mem[1329] : 
                         (N54)? mem[1393] : 
                         (N56)? mem[1457] : 
                         (N58)? mem[1521] : 
                         (N60)? mem[1585] : 
                         (N62)? mem[1649] : 
                         (N64)? mem[1713] : 
                         (N66)? mem[1777] : 
                         (N68)? mem[1841] : 
                         (N70)? mem[1905] : 
                         (N72)? mem[1969] : 
                         (N74)? mem[2033] : 1'b0;
  assign r0_data_o[48] = (N43)? mem[48] : 
                         (N45)? mem[112] : 
                         (N47)? mem[176] : 
                         (N49)? mem[240] : 
                         (N51)? mem[304] : 
                         (N53)? mem[368] : 
                         (N55)? mem[432] : 
                         (N57)? mem[496] : 
                         (N59)? mem[560] : 
                         (N61)? mem[624] : 
                         (N63)? mem[688] : 
                         (N65)? mem[752] : 
                         (N67)? mem[816] : 
                         (N69)? mem[880] : 
                         (N71)? mem[944] : 
                         (N73)? mem[1008] : 
                         (N44)? mem[1072] : 
                         (N46)? mem[1136] : 
                         (N48)? mem[1200] : 
                         (N50)? mem[1264] : 
                         (N52)? mem[1328] : 
                         (N54)? mem[1392] : 
                         (N56)? mem[1456] : 
                         (N58)? mem[1520] : 
                         (N60)? mem[1584] : 
                         (N62)? mem[1648] : 
                         (N64)? mem[1712] : 
                         (N66)? mem[1776] : 
                         (N68)? mem[1840] : 
                         (N70)? mem[1904] : 
                         (N72)? mem[1968] : 
                         (N74)? mem[2032] : 1'b0;
  assign r0_data_o[47] = (N43)? mem[47] : 
                         (N45)? mem[111] : 
                         (N47)? mem[175] : 
                         (N49)? mem[239] : 
                         (N51)? mem[303] : 
                         (N53)? mem[367] : 
                         (N55)? mem[431] : 
                         (N57)? mem[495] : 
                         (N59)? mem[559] : 
                         (N61)? mem[623] : 
                         (N63)? mem[687] : 
                         (N65)? mem[751] : 
                         (N67)? mem[815] : 
                         (N69)? mem[879] : 
                         (N71)? mem[943] : 
                         (N73)? mem[1007] : 
                         (N44)? mem[1071] : 
                         (N46)? mem[1135] : 
                         (N48)? mem[1199] : 
                         (N50)? mem[1263] : 
                         (N52)? mem[1327] : 
                         (N54)? mem[1391] : 
                         (N56)? mem[1455] : 
                         (N58)? mem[1519] : 
                         (N60)? mem[1583] : 
                         (N62)? mem[1647] : 
                         (N64)? mem[1711] : 
                         (N66)? mem[1775] : 
                         (N68)? mem[1839] : 
                         (N70)? mem[1903] : 
                         (N72)? mem[1967] : 
                         (N74)? mem[2031] : 1'b0;
  assign r0_data_o[46] = (N43)? mem[46] : 
                         (N45)? mem[110] : 
                         (N47)? mem[174] : 
                         (N49)? mem[238] : 
                         (N51)? mem[302] : 
                         (N53)? mem[366] : 
                         (N55)? mem[430] : 
                         (N57)? mem[494] : 
                         (N59)? mem[558] : 
                         (N61)? mem[622] : 
                         (N63)? mem[686] : 
                         (N65)? mem[750] : 
                         (N67)? mem[814] : 
                         (N69)? mem[878] : 
                         (N71)? mem[942] : 
                         (N73)? mem[1006] : 
                         (N44)? mem[1070] : 
                         (N46)? mem[1134] : 
                         (N48)? mem[1198] : 
                         (N50)? mem[1262] : 
                         (N52)? mem[1326] : 
                         (N54)? mem[1390] : 
                         (N56)? mem[1454] : 
                         (N58)? mem[1518] : 
                         (N60)? mem[1582] : 
                         (N62)? mem[1646] : 
                         (N64)? mem[1710] : 
                         (N66)? mem[1774] : 
                         (N68)? mem[1838] : 
                         (N70)? mem[1902] : 
                         (N72)? mem[1966] : 
                         (N74)? mem[2030] : 1'b0;
  assign r0_data_o[45] = (N43)? mem[45] : 
                         (N45)? mem[109] : 
                         (N47)? mem[173] : 
                         (N49)? mem[237] : 
                         (N51)? mem[301] : 
                         (N53)? mem[365] : 
                         (N55)? mem[429] : 
                         (N57)? mem[493] : 
                         (N59)? mem[557] : 
                         (N61)? mem[621] : 
                         (N63)? mem[685] : 
                         (N65)? mem[749] : 
                         (N67)? mem[813] : 
                         (N69)? mem[877] : 
                         (N71)? mem[941] : 
                         (N73)? mem[1005] : 
                         (N44)? mem[1069] : 
                         (N46)? mem[1133] : 
                         (N48)? mem[1197] : 
                         (N50)? mem[1261] : 
                         (N52)? mem[1325] : 
                         (N54)? mem[1389] : 
                         (N56)? mem[1453] : 
                         (N58)? mem[1517] : 
                         (N60)? mem[1581] : 
                         (N62)? mem[1645] : 
                         (N64)? mem[1709] : 
                         (N66)? mem[1773] : 
                         (N68)? mem[1837] : 
                         (N70)? mem[1901] : 
                         (N72)? mem[1965] : 
                         (N74)? mem[2029] : 1'b0;
  assign r0_data_o[44] = (N43)? mem[44] : 
                         (N45)? mem[108] : 
                         (N47)? mem[172] : 
                         (N49)? mem[236] : 
                         (N51)? mem[300] : 
                         (N53)? mem[364] : 
                         (N55)? mem[428] : 
                         (N57)? mem[492] : 
                         (N59)? mem[556] : 
                         (N61)? mem[620] : 
                         (N63)? mem[684] : 
                         (N65)? mem[748] : 
                         (N67)? mem[812] : 
                         (N69)? mem[876] : 
                         (N71)? mem[940] : 
                         (N73)? mem[1004] : 
                         (N44)? mem[1068] : 
                         (N46)? mem[1132] : 
                         (N48)? mem[1196] : 
                         (N50)? mem[1260] : 
                         (N52)? mem[1324] : 
                         (N54)? mem[1388] : 
                         (N56)? mem[1452] : 
                         (N58)? mem[1516] : 
                         (N60)? mem[1580] : 
                         (N62)? mem[1644] : 
                         (N64)? mem[1708] : 
                         (N66)? mem[1772] : 
                         (N68)? mem[1836] : 
                         (N70)? mem[1900] : 
                         (N72)? mem[1964] : 
                         (N74)? mem[2028] : 1'b0;
  assign r0_data_o[43] = (N43)? mem[43] : 
                         (N45)? mem[107] : 
                         (N47)? mem[171] : 
                         (N49)? mem[235] : 
                         (N51)? mem[299] : 
                         (N53)? mem[363] : 
                         (N55)? mem[427] : 
                         (N57)? mem[491] : 
                         (N59)? mem[555] : 
                         (N61)? mem[619] : 
                         (N63)? mem[683] : 
                         (N65)? mem[747] : 
                         (N67)? mem[811] : 
                         (N69)? mem[875] : 
                         (N71)? mem[939] : 
                         (N73)? mem[1003] : 
                         (N44)? mem[1067] : 
                         (N46)? mem[1131] : 
                         (N48)? mem[1195] : 
                         (N50)? mem[1259] : 
                         (N52)? mem[1323] : 
                         (N54)? mem[1387] : 
                         (N56)? mem[1451] : 
                         (N58)? mem[1515] : 
                         (N60)? mem[1579] : 
                         (N62)? mem[1643] : 
                         (N64)? mem[1707] : 
                         (N66)? mem[1771] : 
                         (N68)? mem[1835] : 
                         (N70)? mem[1899] : 
                         (N72)? mem[1963] : 
                         (N74)? mem[2027] : 1'b0;
  assign r0_data_o[42] = (N43)? mem[42] : 
                         (N45)? mem[106] : 
                         (N47)? mem[170] : 
                         (N49)? mem[234] : 
                         (N51)? mem[298] : 
                         (N53)? mem[362] : 
                         (N55)? mem[426] : 
                         (N57)? mem[490] : 
                         (N59)? mem[554] : 
                         (N61)? mem[618] : 
                         (N63)? mem[682] : 
                         (N65)? mem[746] : 
                         (N67)? mem[810] : 
                         (N69)? mem[874] : 
                         (N71)? mem[938] : 
                         (N73)? mem[1002] : 
                         (N44)? mem[1066] : 
                         (N46)? mem[1130] : 
                         (N48)? mem[1194] : 
                         (N50)? mem[1258] : 
                         (N52)? mem[1322] : 
                         (N54)? mem[1386] : 
                         (N56)? mem[1450] : 
                         (N58)? mem[1514] : 
                         (N60)? mem[1578] : 
                         (N62)? mem[1642] : 
                         (N64)? mem[1706] : 
                         (N66)? mem[1770] : 
                         (N68)? mem[1834] : 
                         (N70)? mem[1898] : 
                         (N72)? mem[1962] : 
                         (N74)? mem[2026] : 1'b0;
  assign r0_data_o[41] = (N43)? mem[41] : 
                         (N45)? mem[105] : 
                         (N47)? mem[169] : 
                         (N49)? mem[233] : 
                         (N51)? mem[297] : 
                         (N53)? mem[361] : 
                         (N55)? mem[425] : 
                         (N57)? mem[489] : 
                         (N59)? mem[553] : 
                         (N61)? mem[617] : 
                         (N63)? mem[681] : 
                         (N65)? mem[745] : 
                         (N67)? mem[809] : 
                         (N69)? mem[873] : 
                         (N71)? mem[937] : 
                         (N73)? mem[1001] : 
                         (N44)? mem[1065] : 
                         (N46)? mem[1129] : 
                         (N48)? mem[1193] : 
                         (N50)? mem[1257] : 
                         (N52)? mem[1321] : 
                         (N54)? mem[1385] : 
                         (N56)? mem[1449] : 
                         (N58)? mem[1513] : 
                         (N60)? mem[1577] : 
                         (N62)? mem[1641] : 
                         (N64)? mem[1705] : 
                         (N66)? mem[1769] : 
                         (N68)? mem[1833] : 
                         (N70)? mem[1897] : 
                         (N72)? mem[1961] : 
                         (N74)? mem[2025] : 1'b0;
  assign r0_data_o[40] = (N43)? mem[40] : 
                         (N45)? mem[104] : 
                         (N47)? mem[168] : 
                         (N49)? mem[232] : 
                         (N51)? mem[296] : 
                         (N53)? mem[360] : 
                         (N55)? mem[424] : 
                         (N57)? mem[488] : 
                         (N59)? mem[552] : 
                         (N61)? mem[616] : 
                         (N63)? mem[680] : 
                         (N65)? mem[744] : 
                         (N67)? mem[808] : 
                         (N69)? mem[872] : 
                         (N71)? mem[936] : 
                         (N73)? mem[1000] : 
                         (N44)? mem[1064] : 
                         (N46)? mem[1128] : 
                         (N48)? mem[1192] : 
                         (N50)? mem[1256] : 
                         (N52)? mem[1320] : 
                         (N54)? mem[1384] : 
                         (N56)? mem[1448] : 
                         (N58)? mem[1512] : 
                         (N60)? mem[1576] : 
                         (N62)? mem[1640] : 
                         (N64)? mem[1704] : 
                         (N66)? mem[1768] : 
                         (N68)? mem[1832] : 
                         (N70)? mem[1896] : 
                         (N72)? mem[1960] : 
                         (N74)? mem[2024] : 1'b0;
  assign r0_data_o[39] = (N43)? mem[39] : 
                         (N45)? mem[103] : 
                         (N47)? mem[167] : 
                         (N49)? mem[231] : 
                         (N51)? mem[295] : 
                         (N53)? mem[359] : 
                         (N55)? mem[423] : 
                         (N57)? mem[487] : 
                         (N59)? mem[551] : 
                         (N61)? mem[615] : 
                         (N63)? mem[679] : 
                         (N65)? mem[743] : 
                         (N67)? mem[807] : 
                         (N69)? mem[871] : 
                         (N71)? mem[935] : 
                         (N73)? mem[999] : 
                         (N44)? mem[1063] : 
                         (N46)? mem[1127] : 
                         (N48)? mem[1191] : 
                         (N50)? mem[1255] : 
                         (N52)? mem[1319] : 
                         (N54)? mem[1383] : 
                         (N56)? mem[1447] : 
                         (N58)? mem[1511] : 
                         (N60)? mem[1575] : 
                         (N62)? mem[1639] : 
                         (N64)? mem[1703] : 
                         (N66)? mem[1767] : 
                         (N68)? mem[1831] : 
                         (N70)? mem[1895] : 
                         (N72)? mem[1959] : 
                         (N74)? mem[2023] : 1'b0;
  assign r0_data_o[38] = (N43)? mem[38] : 
                         (N45)? mem[102] : 
                         (N47)? mem[166] : 
                         (N49)? mem[230] : 
                         (N51)? mem[294] : 
                         (N53)? mem[358] : 
                         (N55)? mem[422] : 
                         (N57)? mem[486] : 
                         (N59)? mem[550] : 
                         (N61)? mem[614] : 
                         (N63)? mem[678] : 
                         (N65)? mem[742] : 
                         (N67)? mem[806] : 
                         (N69)? mem[870] : 
                         (N71)? mem[934] : 
                         (N73)? mem[998] : 
                         (N44)? mem[1062] : 
                         (N46)? mem[1126] : 
                         (N48)? mem[1190] : 
                         (N50)? mem[1254] : 
                         (N52)? mem[1318] : 
                         (N54)? mem[1382] : 
                         (N56)? mem[1446] : 
                         (N58)? mem[1510] : 
                         (N60)? mem[1574] : 
                         (N62)? mem[1638] : 
                         (N64)? mem[1702] : 
                         (N66)? mem[1766] : 
                         (N68)? mem[1830] : 
                         (N70)? mem[1894] : 
                         (N72)? mem[1958] : 
                         (N74)? mem[2022] : 1'b0;
  assign r0_data_o[37] = (N43)? mem[37] : 
                         (N45)? mem[101] : 
                         (N47)? mem[165] : 
                         (N49)? mem[229] : 
                         (N51)? mem[293] : 
                         (N53)? mem[357] : 
                         (N55)? mem[421] : 
                         (N57)? mem[485] : 
                         (N59)? mem[549] : 
                         (N61)? mem[613] : 
                         (N63)? mem[677] : 
                         (N65)? mem[741] : 
                         (N67)? mem[805] : 
                         (N69)? mem[869] : 
                         (N71)? mem[933] : 
                         (N73)? mem[997] : 
                         (N44)? mem[1061] : 
                         (N46)? mem[1125] : 
                         (N48)? mem[1189] : 
                         (N50)? mem[1253] : 
                         (N52)? mem[1317] : 
                         (N54)? mem[1381] : 
                         (N56)? mem[1445] : 
                         (N58)? mem[1509] : 
                         (N60)? mem[1573] : 
                         (N62)? mem[1637] : 
                         (N64)? mem[1701] : 
                         (N66)? mem[1765] : 
                         (N68)? mem[1829] : 
                         (N70)? mem[1893] : 
                         (N72)? mem[1957] : 
                         (N74)? mem[2021] : 1'b0;
  assign r0_data_o[36] = (N43)? mem[36] : 
                         (N45)? mem[100] : 
                         (N47)? mem[164] : 
                         (N49)? mem[228] : 
                         (N51)? mem[292] : 
                         (N53)? mem[356] : 
                         (N55)? mem[420] : 
                         (N57)? mem[484] : 
                         (N59)? mem[548] : 
                         (N61)? mem[612] : 
                         (N63)? mem[676] : 
                         (N65)? mem[740] : 
                         (N67)? mem[804] : 
                         (N69)? mem[868] : 
                         (N71)? mem[932] : 
                         (N73)? mem[996] : 
                         (N44)? mem[1060] : 
                         (N46)? mem[1124] : 
                         (N48)? mem[1188] : 
                         (N50)? mem[1252] : 
                         (N52)? mem[1316] : 
                         (N54)? mem[1380] : 
                         (N56)? mem[1444] : 
                         (N58)? mem[1508] : 
                         (N60)? mem[1572] : 
                         (N62)? mem[1636] : 
                         (N64)? mem[1700] : 
                         (N66)? mem[1764] : 
                         (N68)? mem[1828] : 
                         (N70)? mem[1892] : 
                         (N72)? mem[1956] : 
                         (N74)? mem[2020] : 1'b0;
  assign r0_data_o[35] = (N43)? mem[35] : 
                         (N45)? mem[99] : 
                         (N47)? mem[163] : 
                         (N49)? mem[227] : 
                         (N51)? mem[291] : 
                         (N53)? mem[355] : 
                         (N55)? mem[419] : 
                         (N57)? mem[483] : 
                         (N59)? mem[547] : 
                         (N61)? mem[611] : 
                         (N63)? mem[675] : 
                         (N65)? mem[739] : 
                         (N67)? mem[803] : 
                         (N69)? mem[867] : 
                         (N71)? mem[931] : 
                         (N73)? mem[995] : 
                         (N44)? mem[1059] : 
                         (N46)? mem[1123] : 
                         (N48)? mem[1187] : 
                         (N50)? mem[1251] : 
                         (N52)? mem[1315] : 
                         (N54)? mem[1379] : 
                         (N56)? mem[1443] : 
                         (N58)? mem[1507] : 
                         (N60)? mem[1571] : 
                         (N62)? mem[1635] : 
                         (N64)? mem[1699] : 
                         (N66)? mem[1763] : 
                         (N68)? mem[1827] : 
                         (N70)? mem[1891] : 
                         (N72)? mem[1955] : 
                         (N74)? mem[2019] : 1'b0;
  assign r0_data_o[34] = (N43)? mem[34] : 
                         (N45)? mem[98] : 
                         (N47)? mem[162] : 
                         (N49)? mem[226] : 
                         (N51)? mem[290] : 
                         (N53)? mem[354] : 
                         (N55)? mem[418] : 
                         (N57)? mem[482] : 
                         (N59)? mem[546] : 
                         (N61)? mem[610] : 
                         (N63)? mem[674] : 
                         (N65)? mem[738] : 
                         (N67)? mem[802] : 
                         (N69)? mem[866] : 
                         (N71)? mem[930] : 
                         (N73)? mem[994] : 
                         (N44)? mem[1058] : 
                         (N46)? mem[1122] : 
                         (N48)? mem[1186] : 
                         (N50)? mem[1250] : 
                         (N52)? mem[1314] : 
                         (N54)? mem[1378] : 
                         (N56)? mem[1442] : 
                         (N58)? mem[1506] : 
                         (N60)? mem[1570] : 
                         (N62)? mem[1634] : 
                         (N64)? mem[1698] : 
                         (N66)? mem[1762] : 
                         (N68)? mem[1826] : 
                         (N70)? mem[1890] : 
                         (N72)? mem[1954] : 
                         (N74)? mem[2018] : 1'b0;
  assign r0_data_o[33] = (N43)? mem[33] : 
                         (N45)? mem[97] : 
                         (N47)? mem[161] : 
                         (N49)? mem[225] : 
                         (N51)? mem[289] : 
                         (N53)? mem[353] : 
                         (N55)? mem[417] : 
                         (N57)? mem[481] : 
                         (N59)? mem[545] : 
                         (N61)? mem[609] : 
                         (N63)? mem[673] : 
                         (N65)? mem[737] : 
                         (N67)? mem[801] : 
                         (N69)? mem[865] : 
                         (N71)? mem[929] : 
                         (N73)? mem[993] : 
                         (N44)? mem[1057] : 
                         (N46)? mem[1121] : 
                         (N48)? mem[1185] : 
                         (N50)? mem[1249] : 
                         (N52)? mem[1313] : 
                         (N54)? mem[1377] : 
                         (N56)? mem[1441] : 
                         (N58)? mem[1505] : 
                         (N60)? mem[1569] : 
                         (N62)? mem[1633] : 
                         (N64)? mem[1697] : 
                         (N66)? mem[1761] : 
                         (N68)? mem[1825] : 
                         (N70)? mem[1889] : 
                         (N72)? mem[1953] : 
                         (N74)? mem[2017] : 1'b0;
  assign r0_data_o[32] = (N43)? mem[32] : 
                         (N45)? mem[96] : 
                         (N47)? mem[160] : 
                         (N49)? mem[224] : 
                         (N51)? mem[288] : 
                         (N53)? mem[352] : 
                         (N55)? mem[416] : 
                         (N57)? mem[480] : 
                         (N59)? mem[544] : 
                         (N61)? mem[608] : 
                         (N63)? mem[672] : 
                         (N65)? mem[736] : 
                         (N67)? mem[800] : 
                         (N69)? mem[864] : 
                         (N71)? mem[928] : 
                         (N73)? mem[992] : 
                         (N44)? mem[1056] : 
                         (N46)? mem[1120] : 
                         (N48)? mem[1184] : 
                         (N50)? mem[1248] : 
                         (N52)? mem[1312] : 
                         (N54)? mem[1376] : 
                         (N56)? mem[1440] : 
                         (N58)? mem[1504] : 
                         (N60)? mem[1568] : 
                         (N62)? mem[1632] : 
                         (N64)? mem[1696] : 
                         (N66)? mem[1760] : 
                         (N68)? mem[1824] : 
                         (N70)? mem[1888] : 
                         (N72)? mem[1952] : 
                         (N74)? mem[2016] : 1'b0;
  assign r0_data_o[31] = (N43)? mem[31] : 
                         (N45)? mem[95] : 
                         (N47)? mem[159] : 
                         (N49)? mem[223] : 
                         (N51)? mem[287] : 
                         (N53)? mem[351] : 
                         (N55)? mem[415] : 
                         (N57)? mem[479] : 
                         (N59)? mem[543] : 
                         (N61)? mem[607] : 
                         (N63)? mem[671] : 
                         (N65)? mem[735] : 
                         (N67)? mem[799] : 
                         (N69)? mem[863] : 
                         (N71)? mem[927] : 
                         (N73)? mem[991] : 
                         (N44)? mem[1055] : 
                         (N46)? mem[1119] : 
                         (N48)? mem[1183] : 
                         (N50)? mem[1247] : 
                         (N52)? mem[1311] : 
                         (N54)? mem[1375] : 
                         (N56)? mem[1439] : 
                         (N58)? mem[1503] : 
                         (N60)? mem[1567] : 
                         (N62)? mem[1631] : 
                         (N64)? mem[1695] : 
                         (N66)? mem[1759] : 
                         (N68)? mem[1823] : 
                         (N70)? mem[1887] : 
                         (N72)? mem[1951] : 
                         (N74)? mem[2015] : 1'b0;
  assign r0_data_o[30] = (N43)? mem[30] : 
                         (N45)? mem[94] : 
                         (N47)? mem[158] : 
                         (N49)? mem[222] : 
                         (N51)? mem[286] : 
                         (N53)? mem[350] : 
                         (N55)? mem[414] : 
                         (N57)? mem[478] : 
                         (N59)? mem[542] : 
                         (N61)? mem[606] : 
                         (N63)? mem[670] : 
                         (N65)? mem[734] : 
                         (N67)? mem[798] : 
                         (N69)? mem[862] : 
                         (N71)? mem[926] : 
                         (N73)? mem[990] : 
                         (N44)? mem[1054] : 
                         (N46)? mem[1118] : 
                         (N48)? mem[1182] : 
                         (N50)? mem[1246] : 
                         (N52)? mem[1310] : 
                         (N54)? mem[1374] : 
                         (N56)? mem[1438] : 
                         (N58)? mem[1502] : 
                         (N60)? mem[1566] : 
                         (N62)? mem[1630] : 
                         (N64)? mem[1694] : 
                         (N66)? mem[1758] : 
                         (N68)? mem[1822] : 
                         (N70)? mem[1886] : 
                         (N72)? mem[1950] : 
                         (N74)? mem[2014] : 1'b0;
  assign r0_data_o[29] = (N43)? mem[29] : 
                         (N45)? mem[93] : 
                         (N47)? mem[157] : 
                         (N49)? mem[221] : 
                         (N51)? mem[285] : 
                         (N53)? mem[349] : 
                         (N55)? mem[413] : 
                         (N57)? mem[477] : 
                         (N59)? mem[541] : 
                         (N61)? mem[605] : 
                         (N63)? mem[669] : 
                         (N65)? mem[733] : 
                         (N67)? mem[797] : 
                         (N69)? mem[861] : 
                         (N71)? mem[925] : 
                         (N73)? mem[989] : 
                         (N44)? mem[1053] : 
                         (N46)? mem[1117] : 
                         (N48)? mem[1181] : 
                         (N50)? mem[1245] : 
                         (N52)? mem[1309] : 
                         (N54)? mem[1373] : 
                         (N56)? mem[1437] : 
                         (N58)? mem[1501] : 
                         (N60)? mem[1565] : 
                         (N62)? mem[1629] : 
                         (N64)? mem[1693] : 
                         (N66)? mem[1757] : 
                         (N68)? mem[1821] : 
                         (N70)? mem[1885] : 
                         (N72)? mem[1949] : 
                         (N74)? mem[2013] : 1'b0;
  assign r0_data_o[28] = (N43)? mem[28] : 
                         (N45)? mem[92] : 
                         (N47)? mem[156] : 
                         (N49)? mem[220] : 
                         (N51)? mem[284] : 
                         (N53)? mem[348] : 
                         (N55)? mem[412] : 
                         (N57)? mem[476] : 
                         (N59)? mem[540] : 
                         (N61)? mem[604] : 
                         (N63)? mem[668] : 
                         (N65)? mem[732] : 
                         (N67)? mem[796] : 
                         (N69)? mem[860] : 
                         (N71)? mem[924] : 
                         (N73)? mem[988] : 
                         (N44)? mem[1052] : 
                         (N46)? mem[1116] : 
                         (N48)? mem[1180] : 
                         (N50)? mem[1244] : 
                         (N52)? mem[1308] : 
                         (N54)? mem[1372] : 
                         (N56)? mem[1436] : 
                         (N58)? mem[1500] : 
                         (N60)? mem[1564] : 
                         (N62)? mem[1628] : 
                         (N64)? mem[1692] : 
                         (N66)? mem[1756] : 
                         (N68)? mem[1820] : 
                         (N70)? mem[1884] : 
                         (N72)? mem[1948] : 
                         (N74)? mem[2012] : 1'b0;
  assign r0_data_o[27] = (N43)? mem[27] : 
                         (N45)? mem[91] : 
                         (N47)? mem[155] : 
                         (N49)? mem[219] : 
                         (N51)? mem[283] : 
                         (N53)? mem[347] : 
                         (N55)? mem[411] : 
                         (N57)? mem[475] : 
                         (N59)? mem[539] : 
                         (N61)? mem[603] : 
                         (N63)? mem[667] : 
                         (N65)? mem[731] : 
                         (N67)? mem[795] : 
                         (N69)? mem[859] : 
                         (N71)? mem[923] : 
                         (N73)? mem[987] : 
                         (N44)? mem[1051] : 
                         (N46)? mem[1115] : 
                         (N48)? mem[1179] : 
                         (N50)? mem[1243] : 
                         (N52)? mem[1307] : 
                         (N54)? mem[1371] : 
                         (N56)? mem[1435] : 
                         (N58)? mem[1499] : 
                         (N60)? mem[1563] : 
                         (N62)? mem[1627] : 
                         (N64)? mem[1691] : 
                         (N66)? mem[1755] : 
                         (N68)? mem[1819] : 
                         (N70)? mem[1883] : 
                         (N72)? mem[1947] : 
                         (N74)? mem[2011] : 1'b0;
  assign r0_data_o[26] = (N43)? mem[26] : 
                         (N45)? mem[90] : 
                         (N47)? mem[154] : 
                         (N49)? mem[218] : 
                         (N51)? mem[282] : 
                         (N53)? mem[346] : 
                         (N55)? mem[410] : 
                         (N57)? mem[474] : 
                         (N59)? mem[538] : 
                         (N61)? mem[602] : 
                         (N63)? mem[666] : 
                         (N65)? mem[730] : 
                         (N67)? mem[794] : 
                         (N69)? mem[858] : 
                         (N71)? mem[922] : 
                         (N73)? mem[986] : 
                         (N44)? mem[1050] : 
                         (N46)? mem[1114] : 
                         (N48)? mem[1178] : 
                         (N50)? mem[1242] : 
                         (N52)? mem[1306] : 
                         (N54)? mem[1370] : 
                         (N56)? mem[1434] : 
                         (N58)? mem[1498] : 
                         (N60)? mem[1562] : 
                         (N62)? mem[1626] : 
                         (N64)? mem[1690] : 
                         (N66)? mem[1754] : 
                         (N68)? mem[1818] : 
                         (N70)? mem[1882] : 
                         (N72)? mem[1946] : 
                         (N74)? mem[2010] : 1'b0;
  assign r0_data_o[25] = (N43)? mem[25] : 
                         (N45)? mem[89] : 
                         (N47)? mem[153] : 
                         (N49)? mem[217] : 
                         (N51)? mem[281] : 
                         (N53)? mem[345] : 
                         (N55)? mem[409] : 
                         (N57)? mem[473] : 
                         (N59)? mem[537] : 
                         (N61)? mem[601] : 
                         (N63)? mem[665] : 
                         (N65)? mem[729] : 
                         (N67)? mem[793] : 
                         (N69)? mem[857] : 
                         (N71)? mem[921] : 
                         (N73)? mem[985] : 
                         (N44)? mem[1049] : 
                         (N46)? mem[1113] : 
                         (N48)? mem[1177] : 
                         (N50)? mem[1241] : 
                         (N52)? mem[1305] : 
                         (N54)? mem[1369] : 
                         (N56)? mem[1433] : 
                         (N58)? mem[1497] : 
                         (N60)? mem[1561] : 
                         (N62)? mem[1625] : 
                         (N64)? mem[1689] : 
                         (N66)? mem[1753] : 
                         (N68)? mem[1817] : 
                         (N70)? mem[1881] : 
                         (N72)? mem[1945] : 
                         (N74)? mem[2009] : 1'b0;
  assign r0_data_o[24] = (N43)? mem[24] : 
                         (N45)? mem[88] : 
                         (N47)? mem[152] : 
                         (N49)? mem[216] : 
                         (N51)? mem[280] : 
                         (N53)? mem[344] : 
                         (N55)? mem[408] : 
                         (N57)? mem[472] : 
                         (N59)? mem[536] : 
                         (N61)? mem[600] : 
                         (N63)? mem[664] : 
                         (N65)? mem[728] : 
                         (N67)? mem[792] : 
                         (N69)? mem[856] : 
                         (N71)? mem[920] : 
                         (N73)? mem[984] : 
                         (N44)? mem[1048] : 
                         (N46)? mem[1112] : 
                         (N48)? mem[1176] : 
                         (N50)? mem[1240] : 
                         (N52)? mem[1304] : 
                         (N54)? mem[1368] : 
                         (N56)? mem[1432] : 
                         (N58)? mem[1496] : 
                         (N60)? mem[1560] : 
                         (N62)? mem[1624] : 
                         (N64)? mem[1688] : 
                         (N66)? mem[1752] : 
                         (N68)? mem[1816] : 
                         (N70)? mem[1880] : 
                         (N72)? mem[1944] : 
                         (N74)? mem[2008] : 1'b0;
  assign r0_data_o[23] = (N43)? mem[23] : 
                         (N45)? mem[87] : 
                         (N47)? mem[151] : 
                         (N49)? mem[215] : 
                         (N51)? mem[279] : 
                         (N53)? mem[343] : 
                         (N55)? mem[407] : 
                         (N57)? mem[471] : 
                         (N59)? mem[535] : 
                         (N61)? mem[599] : 
                         (N63)? mem[663] : 
                         (N65)? mem[727] : 
                         (N67)? mem[791] : 
                         (N69)? mem[855] : 
                         (N71)? mem[919] : 
                         (N73)? mem[983] : 
                         (N44)? mem[1047] : 
                         (N46)? mem[1111] : 
                         (N48)? mem[1175] : 
                         (N50)? mem[1239] : 
                         (N52)? mem[1303] : 
                         (N54)? mem[1367] : 
                         (N56)? mem[1431] : 
                         (N58)? mem[1495] : 
                         (N60)? mem[1559] : 
                         (N62)? mem[1623] : 
                         (N64)? mem[1687] : 
                         (N66)? mem[1751] : 
                         (N68)? mem[1815] : 
                         (N70)? mem[1879] : 
                         (N72)? mem[1943] : 
                         (N74)? mem[2007] : 1'b0;
  assign r0_data_o[22] = (N43)? mem[22] : 
                         (N45)? mem[86] : 
                         (N47)? mem[150] : 
                         (N49)? mem[214] : 
                         (N51)? mem[278] : 
                         (N53)? mem[342] : 
                         (N55)? mem[406] : 
                         (N57)? mem[470] : 
                         (N59)? mem[534] : 
                         (N61)? mem[598] : 
                         (N63)? mem[662] : 
                         (N65)? mem[726] : 
                         (N67)? mem[790] : 
                         (N69)? mem[854] : 
                         (N71)? mem[918] : 
                         (N73)? mem[982] : 
                         (N44)? mem[1046] : 
                         (N46)? mem[1110] : 
                         (N48)? mem[1174] : 
                         (N50)? mem[1238] : 
                         (N52)? mem[1302] : 
                         (N54)? mem[1366] : 
                         (N56)? mem[1430] : 
                         (N58)? mem[1494] : 
                         (N60)? mem[1558] : 
                         (N62)? mem[1622] : 
                         (N64)? mem[1686] : 
                         (N66)? mem[1750] : 
                         (N68)? mem[1814] : 
                         (N70)? mem[1878] : 
                         (N72)? mem[1942] : 
                         (N74)? mem[2006] : 1'b0;
  assign r0_data_o[21] = (N43)? mem[21] : 
                         (N45)? mem[85] : 
                         (N47)? mem[149] : 
                         (N49)? mem[213] : 
                         (N51)? mem[277] : 
                         (N53)? mem[341] : 
                         (N55)? mem[405] : 
                         (N57)? mem[469] : 
                         (N59)? mem[533] : 
                         (N61)? mem[597] : 
                         (N63)? mem[661] : 
                         (N65)? mem[725] : 
                         (N67)? mem[789] : 
                         (N69)? mem[853] : 
                         (N71)? mem[917] : 
                         (N73)? mem[981] : 
                         (N44)? mem[1045] : 
                         (N46)? mem[1109] : 
                         (N48)? mem[1173] : 
                         (N50)? mem[1237] : 
                         (N52)? mem[1301] : 
                         (N54)? mem[1365] : 
                         (N56)? mem[1429] : 
                         (N58)? mem[1493] : 
                         (N60)? mem[1557] : 
                         (N62)? mem[1621] : 
                         (N64)? mem[1685] : 
                         (N66)? mem[1749] : 
                         (N68)? mem[1813] : 
                         (N70)? mem[1877] : 
                         (N72)? mem[1941] : 
                         (N74)? mem[2005] : 1'b0;
  assign r0_data_o[20] = (N43)? mem[20] : 
                         (N45)? mem[84] : 
                         (N47)? mem[148] : 
                         (N49)? mem[212] : 
                         (N51)? mem[276] : 
                         (N53)? mem[340] : 
                         (N55)? mem[404] : 
                         (N57)? mem[468] : 
                         (N59)? mem[532] : 
                         (N61)? mem[596] : 
                         (N63)? mem[660] : 
                         (N65)? mem[724] : 
                         (N67)? mem[788] : 
                         (N69)? mem[852] : 
                         (N71)? mem[916] : 
                         (N73)? mem[980] : 
                         (N44)? mem[1044] : 
                         (N46)? mem[1108] : 
                         (N48)? mem[1172] : 
                         (N50)? mem[1236] : 
                         (N52)? mem[1300] : 
                         (N54)? mem[1364] : 
                         (N56)? mem[1428] : 
                         (N58)? mem[1492] : 
                         (N60)? mem[1556] : 
                         (N62)? mem[1620] : 
                         (N64)? mem[1684] : 
                         (N66)? mem[1748] : 
                         (N68)? mem[1812] : 
                         (N70)? mem[1876] : 
                         (N72)? mem[1940] : 
                         (N74)? mem[2004] : 1'b0;
  assign r0_data_o[19] = (N43)? mem[19] : 
                         (N45)? mem[83] : 
                         (N47)? mem[147] : 
                         (N49)? mem[211] : 
                         (N51)? mem[275] : 
                         (N53)? mem[339] : 
                         (N55)? mem[403] : 
                         (N57)? mem[467] : 
                         (N59)? mem[531] : 
                         (N61)? mem[595] : 
                         (N63)? mem[659] : 
                         (N65)? mem[723] : 
                         (N67)? mem[787] : 
                         (N69)? mem[851] : 
                         (N71)? mem[915] : 
                         (N73)? mem[979] : 
                         (N44)? mem[1043] : 
                         (N46)? mem[1107] : 
                         (N48)? mem[1171] : 
                         (N50)? mem[1235] : 
                         (N52)? mem[1299] : 
                         (N54)? mem[1363] : 
                         (N56)? mem[1427] : 
                         (N58)? mem[1491] : 
                         (N60)? mem[1555] : 
                         (N62)? mem[1619] : 
                         (N64)? mem[1683] : 
                         (N66)? mem[1747] : 
                         (N68)? mem[1811] : 
                         (N70)? mem[1875] : 
                         (N72)? mem[1939] : 
                         (N74)? mem[2003] : 1'b0;
  assign r0_data_o[18] = (N43)? mem[18] : 
                         (N45)? mem[82] : 
                         (N47)? mem[146] : 
                         (N49)? mem[210] : 
                         (N51)? mem[274] : 
                         (N53)? mem[338] : 
                         (N55)? mem[402] : 
                         (N57)? mem[466] : 
                         (N59)? mem[530] : 
                         (N61)? mem[594] : 
                         (N63)? mem[658] : 
                         (N65)? mem[722] : 
                         (N67)? mem[786] : 
                         (N69)? mem[850] : 
                         (N71)? mem[914] : 
                         (N73)? mem[978] : 
                         (N44)? mem[1042] : 
                         (N46)? mem[1106] : 
                         (N48)? mem[1170] : 
                         (N50)? mem[1234] : 
                         (N52)? mem[1298] : 
                         (N54)? mem[1362] : 
                         (N56)? mem[1426] : 
                         (N58)? mem[1490] : 
                         (N60)? mem[1554] : 
                         (N62)? mem[1618] : 
                         (N64)? mem[1682] : 
                         (N66)? mem[1746] : 
                         (N68)? mem[1810] : 
                         (N70)? mem[1874] : 
                         (N72)? mem[1938] : 
                         (N74)? mem[2002] : 1'b0;
  assign r0_data_o[17] = (N43)? mem[17] : 
                         (N45)? mem[81] : 
                         (N47)? mem[145] : 
                         (N49)? mem[209] : 
                         (N51)? mem[273] : 
                         (N53)? mem[337] : 
                         (N55)? mem[401] : 
                         (N57)? mem[465] : 
                         (N59)? mem[529] : 
                         (N61)? mem[593] : 
                         (N63)? mem[657] : 
                         (N65)? mem[721] : 
                         (N67)? mem[785] : 
                         (N69)? mem[849] : 
                         (N71)? mem[913] : 
                         (N73)? mem[977] : 
                         (N44)? mem[1041] : 
                         (N46)? mem[1105] : 
                         (N48)? mem[1169] : 
                         (N50)? mem[1233] : 
                         (N52)? mem[1297] : 
                         (N54)? mem[1361] : 
                         (N56)? mem[1425] : 
                         (N58)? mem[1489] : 
                         (N60)? mem[1553] : 
                         (N62)? mem[1617] : 
                         (N64)? mem[1681] : 
                         (N66)? mem[1745] : 
                         (N68)? mem[1809] : 
                         (N70)? mem[1873] : 
                         (N72)? mem[1937] : 
                         (N74)? mem[2001] : 1'b0;
  assign r0_data_o[16] = (N43)? mem[16] : 
                         (N45)? mem[80] : 
                         (N47)? mem[144] : 
                         (N49)? mem[208] : 
                         (N51)? mem[272] : 
                         (N53)? mem[336] : 
                         (N55)? mem[400] : 
                         (N57)? mem[464] : 
                         (N59)? mem[528] : 
                         (N61)? mem[592] : 
                         (N63)? mem[656] : 
                         (N65)? mem[720] : 
                         (N67)? mem[784] : 
                         (N69)? mem[848] : 
                         (N71)? mem[912] : 
                         (N73)? mem[976] : 
                         (N44)? mem[1040] : 
                         (N46)? mem[1104] : 
                         (N48)? mem[1168] : 
                         (N50)? mem[1232] : 
                         (N52)? mem[1296] : 
                         (N54)? mem[1360] : 
                         (N56)? mem[1424] : 
                         (N58)? mem[1488] : 
                         (N60)? mem[1552] : 
                         (N62)? mem[1616] : 
                         (N64)? mem[1680] : 
                         (N66)? mem[1744] : 
                         (N68)? mem[1808] : 
                         (N70)? mem[1872] : 
                         (N72)? mem[1936] : 
                         (N74)? mem[2000] : 1'b0;
  assign r0_data_o[15] = (N43)? mem[15] : 
                         (N45)? mem[79] : 
                         (N47)? mem[143] : 
                         (N49)? mem[207] : 
                         (N51)? mem[271] : 
                         (N53)? mem[335] : 
                         (N55)? mem[399] : 
                         (N57)? mem[463] : 
                         (N59)? mem[527] : 
                         (N61)? mem[591] : 
                         (N63)? mem[655] : 
                         (N65)? mem[719] : 
                         (N67)? mem[783] : 
                         (N69)? mem[847] : 
                         (N71)? mem[911] : 
                         (N73)? mem[975] : 
                         (N44)? mem[1039] : 
                         (N46)? mem[1103] : 
                         (N48)? mem[1167] : 
                         (N50)? mem[1231] : 
                         (N52)? mem[1295] : 
                         (N54)? mem[1359] : 
                         (N56)? mem[1423] : 
                         (N58)? mem[1487] : 
                         (N60)? mem[1551] : 
                         (N62)? mem[1615] : 
                         (N64)? mem[1679] : 
                         (N66)? mem[1743] : 
                         (N68)? mem[1807] : 
                         (N70)? mem[1871] : 
                         (N72)? mem[1935] : 
                         (N74)? mem[1999] : 1'b0;
  assign r0_data_o[14] = (N43)? mem[14] : 
                         (N45)? mem[78] : 
                         (N47)? mem[142] : 
                         (N49)? mem[206] : 
                         (N51)? mem[270] : 
                         (N53)? mem[334] : 
                         (N55)? mem[398] : 
                         (N57)? mem[462] : 
                         (N59)? mem[526] : 
                         (N61)? mem[590] : 
                         (N63)? mem[654] : 
                         (N65)? mem[718] : 
                         (N67)? mem[782] : 
                         (N69)? mem[846] : 
                         (N71)? mem[910] : 
                         (N73)? mem[974] : 
                         (N44)? mem[1038] : 
                         (N46)? mem[1102] : 
                         (N48)? mem[1166] : 
                         (N50)? mem[1230] : 
                         (N52)? mem[1294] : 
                         (N54)? mem[1358] : 
                         (N56)? mem[1422] : 
                         (N58)? mem[1486] : 
                         (N60)? mem[1550] : 
                         (N62)? mem[1614] : 
                         (N64)? mem[1678] : 
                         (N66)? mem[1742] : 
                         (N68)? mem[1806] : 
                         (N70)? mem[1870] : 
                         (N72)? mem[1934] : 
                         (N74)? mem[1998] : 1'b0;
  assign r0_data_o[13] = (N43)? mem[13] : 
                         (N45)? mem[77] : 
                         (N47)? mem[141] : 
                         (N49)? mem[205] : 
                         (N51)? mem[269] : 
                         (N53)? mem[333] : 
                         (N55)? mem[397] : 
                         (N57)? mem[461] : 
                         (N59)? mem[525] : 
                         (N61)? mem[589] : 
                         (N63)? mem[653] : 
                         (N65)? mem[717] : 
                         (N67)? mem[781] : 
                         (N69)? mem[845] : 
                         (N71)? mem[909] : 
                         (N73)? mem[973] : 
                         (N44)? mem[1037] : 
                         (N46)? mem[1101] : 
                         (N48)? mem[1165] : 
                         (N50)? mem[1229] : 
                         (N52)? mem[1293] : 
                         (N54)? mem[1357] : 
                         (N56)? mem[1421] : 
                         (N58)? mem[1485] : 
                         (N60)? mem[1549] : 
                         (N62)? mem[1613] : 
                         (N64)? mem[1677] : 
                         (N66)? mem[1741] : 
                         (N68)? mem[1805] : 
                         (N70)? mem[1869] : 
                         (N72)? mem[1933] : 
                         (N74)? mem[1997] : 1'b0;
  assign r0_data_o[12] = (N43)? mem[12] : 
                         (N45)? mem[76] : 
                         (N47)? mem[140] : 
                         (N49)? mem[204] : 
                         (N51)? mem[268] : 
                         (N53)? mem[332] : 
                         (N55)? mem[396] : 
                         (N57)? mem[460] : 
                         (N59)? mem[524] : 
                         (N61)? mem[588] : 
                         (N63)? mem[652] : 
                         (N65)? mem[716] : 
                         (N67)? mem[780] : 
                         (N69)? mem[844] : 
                         (N71)? mem[908] : 
                         (N73)? mem[972] : 
                         (N44)? mem[1036] : 
                         (N46)? mem[1100] : 
                         (N48)? mem[1164] : 
                         (N50)? mem[1228] : 
                         (N52)? mem[1292] : 
                         (N54)? mem[1356] : 
                         (N56)? mem[1420] : 
                         (N58)? mem[1484] : 
                         (N60)? mem[1548] : 
                         (N62)? mem[1612] : 
                         (N64)? mem[1676] : 
                         (N66)? mem[1740] : 
                         (N68)? mem[1804] : 
                         (N70)? mem[1868] : 
                         (N72)? mem[1932] : 
                         (N74)? mem[1996] : 1'b0;
  assign r0_data_o[11] = (N43)? mem[11] : 
                         (N45)? mem[75] : 
                         (N47)? mem[139] : 
                         (N49)? mem[203] : 
                         (N51)? mem[267] : 
                         (N53)? mem[331] : 
                         (N55)? mem[395] : 
                         (N57)? mem[459] : 
                         (N59)? mem[523] : 
                         (N61)? mem[587] : 
                         (N63)? mem[651] : 
                         (N65)? mem[715] : 
                         (N67)? mem[779] : 
                         (N69)? mem[843] : 
                         (N71)? mem[907] : 
                         (N73)? mem[971] : 
                         (N44)? mem[1035] : 
                         (N46)? mem[1099] : 
                         (N48)? mem[1163] : 
                         (N50)? mem[1227] : 
                         (N52)? mem[1291] : 
                         (N54)? mem[1355] : 
                         (N56)? mem[1419] : 
                         (N58)? mem[1483] : 
                         (N60)? mem[1547] : 
                         (N62)? mem[1611] : 
                         (N64)? mem[1675] : 
                         (N66)? mem[1739] : 
                         (N68)? mem[1803] : 
                         (N70)? mem[1867] : 
                         (N72)? mem[1931] : 
                         (N74)? mem[1995] : 1'b0;
  assign r0_data_o[10] = (N43)? mem[10] : 
                         (N45)? mem[74] : 
                         (N47)? mem[138] : 
                         (N49)? mem[202] : 
                         (N51)? mem[266] : 
                         (N53)? mem[330] : 
                         (N55)? mem[394] : 
                         (N57)? mem[458] : 
                         (N59)? mem[522] : 
                         (N61)? mem[586] : 
                         (N63)? mem[650] : 
                         (N65)? mem[714] : 
                         (N67)? mem[778] : 
                         (N69)? mem[842] : 
                         (N71)? mem[906] : 
                         (N73)? mem[970] : 
                         (N44)? mem[1034] : 
                         (N46)? mem[1098] : 
                         (N48)? mem[1162] : 
                         (N50)? mem[1226] : 
                         (N52)? mem[1290] : 
                         (N54)? mem[1354] : 
                         (N56)? mem[1418] : 
                         (N58)? mem[1482] : 
                         (N60)? mem[1546] : 
                         (N62)? mem[1610] : 
                         (N64)? mem[1674] : 
                         (N66)? mem[1738] : 
                         (N68)? mem[1802] : 
                         (N70)? mem[1866] : 
                         (N72)? mem[1930] : 
                         (N74)? mem[1994] : 1'b0;
  assign r0_data_o[9] = (N43)? mem[9] : 
                        (N45)? mem[73] : 
                        (N47)? mem[137] : 
                        (N49)? mem[201] : 
                        (N51)? mem[265] : 
                        (N53)? mem[329] : 
                        (N55)? mem[393] : 
                        (N57)? mem[457] : 
                        (N59)? mem[521] : 
                        (N61)? mem[585] : 
                        (N63)? mem[649] : 
                        (N65)? mem[713] : 
                        (N67)? mem[777] : 
                        (N69)? mem[841] : 
                        (N71)? mem[905] : 
                        (N73)? mem[969] : 
                        (N44)? mem[1033] : 
                        (N46)? mem[1097] : 
                        (N48)? mem[1161] : 
                        (N50)? mem[1225] : 
                        (N52)? mem[1289] : 
                        (N54)? mem[1353] : 
                        (N56)? mem[1417] : 
                        (N58)? mem[1481] : 
                        (N60)? mem[1545] : 
                        (N62)? mem[1609] : 
                        (N64)? mem[1673] : 
                        (N66)? mem[1737] : 
                        (N68)? mem[1801] : 
                        (N70)? mem[1865] : 
                        (N72)? mem[1929] : 
                        (N74)? mem[1993] : 1'b0;
  assign r0_data_o[8] = (N43)? mem[8] : 
                        (N45)? mem[72] : 
                        (N47)? mem[136] : 
                        (N49)? mem[200] : 
                        (N51)? mem[264] : 
                        (N53)? mem[328] : 
                        (N55)? mem[392] : 
                        (N57)? mem[456] : 
                        (N59)? mem[520] : 
                        (N61)? mem[584] : 
                        (N63)? mem[648] : 
                        (N65)? mem[712] : 
                        (N67)? mem[776] : 
                        (N69)? mem[840] : 
                        (N71)? mem[904] : 
                        (N73)? mem[968] : 
                        (N44)? mem[1032] : 
                        (N46)? mem[1096] : 
                        (N48)? mem[1160] : 
                        (N50)? mem[1224] : 
                        (N52)? mem[1288] : 
                        (N54)? mem[1352] : 
                        (N56)? mem[1416] : 
                        (N58)? mem[1480] : 
                        (N60)? mem[1544] : 
                        (N62)? mem[1608] : 
                        (N64)? mem[1672] : 
                        (N66)? mem[1736] : 
                        (N68)? mem[1800] : 
                        (N70)? mem[1864] : 
                        (N72)? mem[1928] : 
                        (N74)? mem[1992] : 1'b0;
  assign r0_data_o[7] = (N43)? mem[7] : 
                        (N45)? mem[71] : 
                        (N47)? mem[135] : 
                        (N49)? mem[199] : 
                        (N51)? mem[263] : 
                        (N53)? mem[327] : 
                        (N55)? mem[391] : 
                        (N57)? mem[455] : 
                        (N59)? mem[519] : 
                        (N61)? mem[583] : 
                        (N63)? mem[647] : 
                        (N65)? mem[711] : 
                        (N67)? mem[775] : 
                        (N69)? mem[839] : 
                        (N71)? mem[903] : 
                        (N73)? mem[967] : 
                        (N44)? mem[1031] : 
                        (N46)? mem[1095] : 
                        (N48)? mem[1159] : 
                        (N50)? mem[1223] : 
                        (N52)? mem[1287] : 
                        (N54)? mem[1351] : 
                        (N56)? mem[1415] : 
                        (N58)? mem[1479] : 
                        (N60)? mem[1543] : 
                        (N62)? mem[1607] : 
                        (N64)? mem[1671] : 
                        (N66)? mem[1735] : 
                        (N68)? mem[1799] : 
                        (N70)? mem[1863] : 
                        (N72)? mem[1927] : 
                        (N74)? mem[1991] : 1'b0;
  assign r0_data_o[6] = (N43)? mem[6] : 
                        (N45)? mem[70] : 
                        (N47)? mem[134] : 
                        (N49)? mem[198] : 
                        (N51)? mem[262] : 
                        (N53)? mem[326] : 
                        (N55)? mem[390] : 
                        (N57)? mem[454] : 
                        (N59)? mem[518] : 
                        (N61)? mem[582] : 
                        (N63)? mem[646] : 
                        (N65)? mem[710] : 
                        (N67)? mem[774] : 
                        (N69)? mem[838] : 
                        (N71)? mem[902] : 
                        (N73)? mem[966] : 
                        (N44)? mem[1030] : 
                        (N46)? mem[1094] : 
                        (N48)? mem[1158] : 
                        (N50)? mem[1222] : 
                        (N52)? mem[1286] : 
                        (N54)? mem[1350] : 
                        (N56)? mem[1414] : 
                        (N58)? mem[1478] : 
                        (N60)? mem[1542] : 
                        (N62)? mem[1606] : 
                        (N64)? mem[1670] : 
                        (N66)? mem[1734] : 
                        (N68)? mem[1798] : 
                        (N70)? mem[1862] : 
                        (N72)? mem[1926] : 
                        (N74)? mem[1990] : 1'b0;
  assign r0_data_o[5] = (N43)? mem[5] : 
                        (N45)? mem[69] : 
                        (N47)? mem[133] : 
                        (N49)? mem[197] : 
                        (N51)? mem[261] : 
                        (N53)? mem[325] : 
                        (N55)? mem[389] : 
                        (N57)? mem[453] : 
                        (N59)? mem[517] : 
                        (N61)? mem[581] : 
                        (N63)? mem[645] : 
                        (N65)? mem[709] : 
                        (N67)? mem[773] : 
                        (N69)? mem[837] : 
                        (N71)? mem[901] : 
                        (N73)? mem[965] : 
                        (N44)? mem[1029] : 
                        (N46)? mem[1093] : 
                        (N48)? mem[1157] : 
                        (N50)? mem[1221] : 
                        (N52)? mem[1285] : 
                        (N54)? mem[1349] : 
                        (N56)? mem[1413] : 
                        (N58)? mem[1477] : 
                        (N60)? mem[1541] : 
                        (N62)? mem[1605] : 
                        (N64)? mem[1669] : 
                        (N66)? mem[1733] : 
                        (N68)? mem[1797] : 
                        (N70)? mem[1861] : 
                        (N72)? mem[1925] : 
                        (N74)? mem[1989] : 1'b0;
  assign r0_data_o[4] = (N43)? mem[4] : 
                        (N45)? mem[68] : 
                        (N47)? mem[132] : 
                        (N49)? mem[196] : 
                        (N51)? mem[260] : 
                        (N53)? mem[324] : 
                        (N55)? mem[388] : 
                        (N57)? mem[452] : 
                        (N59)? mem[516] : 
                        (N61)? mem[580] : 
                        (N63)? mem[644] : 
                        (N65)? mem[708] : 
                        (N67)? mem[772] : 
                        (N69)? mem[836] : 
                        (N71)? mem[900] : 
                        (N73)? mem[964] : 
                        (N44)? mem[1028] : 
                        (N46)? mem[1092] : 
                        (N48)? mem[1156] : 
                        (N50)? mem[1220] : 
                        (N52)? mem[1284] : 
                        (N54)? mem[1348] : 
                        (N56)? mem[1412] : 
                        (N58)? mem[1476] : 
                        (N60)? mem[1540] : 
                        (N62)? mem[1604] : 
                        (N64)? mem[1668] : 
                        (N66)? mem[1732] : 
                        (N68)? mem[1796] : 
                        (N70)? mem[1860] : 
                        (N72)? mem[1924] : 
                        (N74)? mem[1988] : 1'b0;
  assign r0_data_o[3] = (N43)? mem[3] : 
                        (N45)? mem[67] : 
                        (N47)? mem[131] : 
                        (N49)? mem[195] : 
                        (N51)? mem[259] : 
                        (N53)? mem[323] : 
                        (N55)? mem[387] : 
                        (N57)? mem[451] : 
                        (N59)? mem[515] : 
                        (N61)? mem[579] : 
                        (N63)? mem[643] : 
                        (N65)? mem[707] : 
                        (N67)? mem[771] : 
                        (N69)? mem[835] : 
                        (N71)? mem[899] : 
                        (N73)? mem[963] : 
                        (N44)? mem[1027] : 
                        (N46)? mem[1091] : 
                        (N48)? mem[1155] : 
                        (N50)? mem[1219] : 
                        (N52)? mem[1283] : 
                        (N54)? mem[1347] : 
                        (N56)? mem[1411] : 
                        (N58)? mem[1475] : 
                        (N60)? mem[1539] : 
                        (N62)? mem[1603] : 
                        (N64)? mem[1667] : 
                        (N66)? mem[1731] : 
                        (N68)? mem[1795] : 
                        (N70)? mem[1859] : 
                        (N72)? mem[1923] : 
                        (N74)? mem[1987] : 1'b0;
  assign r0_data_o[2] = (N43)? mem[2] : 
                        (N45)? mem[66] : 
                        (N47)? mem[130] : 
                        (N49)? mem[194] : 
                        (N51)? mem[258] : 
                        (N53)? mem[322] : 
                        (N55)? mem[386] : 
                        (N57)? mem[450] : 
                        (N59)? mem[514] : 
                        (N61)? mem[578] : 
                        (N63)? mem[642] : 
                        (N65)? mem[706] : 
                        (N67)? mem[770] : 
                        (N69)? mem[834] : 
                        (N71)? mem[898] : 
                        (N73)? mem[962] : 
                        (N44)? mem[1026] : 
                        (N46)? mem[1090] : 
                        (N48)? mem[1154] : 
                        (N50)? mem[1218] : 
                        (N52)? mem[1282] : 
                        (N54)? mem[1346] : 
                        (N56)? mem[1410] : 
                        (N58)? mem[1474] : 
                        (N60)? mem[1538] : 
                        (N62)? mem[1602] : 
                        (N64)? mem[1666] : 
                        (N66)? mem[1730] : 
                        (N68)? mem[1794] : 
                        (N70)? mem[1858] : 
                        (N72)? mem[1922] : 
                        (N74)? mem[1986] : 1'b0;
  assign r0_data_o[1] = (N43)? mem[1] : 
                        (N45)? mem[65] : 
                        (N47)? mem[129] : 
                        (N49)? mem[193] : 
                        (N51)? mem[257] : 
                        (N53)? mem[321] : 
                        (N55)? mem[385] : 
                        (N57)? mem[449] : 
                        (N59)? mem[513] : 
                        (N61)? mem[577] : 
                        (N63)? mem[641] : 
                        (N65)? mem[705] : 
                        (N67)? mem[769] : 
                        (N69)? mem[833] : 
                        (N71)? mem[897] : 
                        (N73)? mem[961] : 
                        (N44)? mem[1025] : 
                        (N46)? mem[1089] : 
                        (N48)? mem[1153] : 
                        (N50)? mem[1217] : 
                        (N52)? mem[1281] : 
                        (N54)? mem[1345] : 
                        (N56)? mem[1409] : 
                        (N58)? mem[1473] : 
                        (N60)? mem[1537] : 
                        (N62)? mem[1601] : 
                        (N64)? mem[1665] : 
                        (N66)? mem[1729] : 
                        (N68)? mem[1793] : 
                        (N70)? mem[1857] : 
                        (N72)? mem[1921] : 
                        (N74)? mem[1985] : 1'b0;
  assign r0_data_o[0] = (N43)? mem[0] : 
                        (N45)? mem[64] : 
                        (N47)? mem[128] : 
                        (N49)? mem[192] : 
                        (N51)? mem[256] : 
                        (N53)? mem[320] : 
                        (N55)? mem[384] : 
                        (N57)? mem[448] : 
                        (N59)? mem[512] : 
                        (N61)? mem[576] : 
                        (N63)? mem[640] : 
                        (N65)? mem[704] : 
                        (N67)? mem[768] : 
                        (N69)? mem[832] : 
                        (N71)? mem[896] : 
                        (N73)? mem[960] : 
                        (N44)? mem[1024] : 
                        (N46)? mem[1088] : 
                        (N48)? mem[1152] : 
                        (N50)? mem[1216] : 
                        (N52)? mem[1280] : 
                        (N54)? mem[1344] : 
                        (N56)? mem[1408] : 
                        (N58)? mem[1472] : 
                        (N60)? mem[1536] : 
                        (N62)? mem[1600] : 
                        (N64)? mem[1664] : 
                        (N66)? mem[1728] : 
                        (N68)? mem[1792] : 
                        (N70)? mem[1856] : 
                        (N72)? mem[1920] : 
                        (N74)? mem[1984] : 1'b0;
  assign r1_data_o[63] = (N108)? mem[63] : 
                         (N110)? mem[127] : 
                         (N112)? mem[191] : 
                         (N114)? mem[255] : 
                         (N116)? mem[319] : 
                         (N118)? mem[383] : 
                         (N120)? mem[447] : 
                         (N122)? mem[511] : 
                         (N124)? mem[575] : 
                         (N126)? mem[639] : 
                         (N128)? mem[703] : 
                         (N130)? mem[767] : 
                         (N132)? mem[831] : 
                         (N134)? mem[895] : 
                         (N136)? mem[959] : 
                         (N138)? mem[1023] : 
                         (N109)? mem[1087] : 
                         (N111)? mem[1151] : 
                         (N113)? mem[1215] : 
                         (N115)? mem[1279] : 
                         (N117)? mem[1343] : 
                         (N119)? mem[1407] : 
                         (N121)? mem[1471] : 
                         (N123)? mem[1535] : 
                         (N125)? mem[1599] : 
                         (N127)? mem[1663] : 
                         (N129)? mem[1727] : 
                         (N131)? mem[1791] : 
                         (N133)? mem[1855] : 
                         (N135)? mem[1919] : 
                         (N137)? mem[1983] : 
                         (N139)? mem[2047] : 1'b0;
  assign r1_data_o[62] = (N108)? mem[62] : 
                         (N110)? mem[126] : 
                         (N112)? mem[190] : 
                         (N114)? mem[254] : 
                         (N116)? mem[318] : 
                         (N118)? mem[382] : 
                         (N120)? mem[446] : 
                         (N122)? mem[510] : 
                         (N124)? mem[574] : 
                         (N126)? mem[638] : 
                         (N128)? mem[702] : 
                         (N130)? mem[766] : 
                         (N132)? mem[830] : 
                         (N134)? mem[894] : 
                         (N136)? mem[958] : 
                         (N138)? mem[1022] : 
                         (N109)? mem[1086] : 
                         (N111)? mem[1150] : 
                         (N113)? mem[1214] : 
                         (N115)? mem[1278] : 
                         (N117)? mem[1342] : 
                         (N119)? mem[1406] : 
                         (N121)? mem[1470] : 
                         (N123)? mem[1534] : 
                         (N125)? mem[1598] : 
                         (N127)? mem[1662] : 
                         (N129)? mem[1726] : 
                         (N131)? mem[1790] : 
                         (N133)? mem[1854] : 
                         (N135)? mem[1918] : 
                         (N137)? mem[1982] : 
                         (N139)? mem[2046] : 1'b0;
  assign r1_data_o[61] = (N108)? mem[61] : 
                         (N110)? mem[125] : 
                         (N112)? mem[189] : 
                         (N114)? mem[253] : 
                         (N116)? mem[317] : 
                         (N118)? mem[381] : 
                         (N120)? mem[445] : 
                         (N122)? mem[509] : 
                         (N124)? mem[573] : 
                         (N126)? mem[637] : 
                         (N128)? mem[701] : 
                         (N130)? mem[765] : 
                         (N132)? mem[829] : 
                         (N134)? mem[893] : 
                         (N136)? mem[957] : 
                         (N138)? mem[1021] : 
                         (N109)? mem[1085] : 
                         (N111)? mem[1149] : 
                         (N113)? mem[1213] : 
                         (N115)? mem[1277] : 
                         (N117)? mem[1341] : 
                         (N119)? mem[1405] : 
                         (N121)? mem[1469] : 
                         (N123)? mem[1533] : 
                         (N125)? mem[1597] : 
                         (N127)? mem[1661] : 
                         (N129)? mem[1725] : 
                         (N131)? mem[1789] : 
                         (N133)? mem[1853] : 
                         (N135)? mem[1917] : 
                         (N137)? mem[1981] : 
                         (N139)? mem[2045] : 1'b0;
  assign r1_data_o[60] = (N108)? mem[60] : 
                         (N110)? mem[124] : 
                         (N112)? mem[188] : 
                         (N114)? mem[252] : 
                         (N116)? mem[316] : 
                         (N118)? mem[380] : 
                         (N120)? mem[444] : 
                         (N122)? mem[508] : 
                         (N124)? mem[572] : 
                         (N126)? mem[636] : 
                         (N128)? mem[700] : 
                         (N130)? mem[764] : 
                         (N132)? mem[828] : 
                         (N134)? mem[892] : 
                         (N136)? mem[956] : 
                         (N138)? mem[1020] : 
                         (N109)? mem[1084] : 
                         (N111)? mem[1148] : 
                         (N113)? mem[1212] : 
                         (N115)? mem[1276] : 
                         (N117)? mem[1340] : 
                         (N119)? mem[1404] : 
                         (N121)? mem[1468] : 
                         (N123)? mem[1532] : 
                         (N125)? mem[1596] : 
                         (N127)? mem[1660] : 
                         (N129)? mem[1724] : 
                         (N131)? mem[1788] : 
                         (N133)? mem[1852] : 
                         (N135)? mem[1916] : 
                         (N137)? mem[1980] : 
                         (N139)? mem[2044] : 1'b0;
  assign r1_data_o[59] = (N108)? mem[59] : 
                         (N110)? mem[123] : 
                         (N112)? mem[187] : 
                         (N114)? mem[251] : 
                         (N116)? mem[315] : 
                         (N118)? mem[379] : 
                         (N120)? mem[443] : 
                         (N122)? mem[507] : 
                         (N124)? mem[571] : 
                         (N126)? mem[635] : 
                         (N128)? mem[699] : 
                         (N130)? mem[763] : 
                         (N132)? mem[827] : 
                         (N134)? mem[891] : 
                         (N136)? mem[955] : 
                         (N138)? mem[1019] : 
                         (N109)? mem[1083] : 
                         (N111)? mem[1147] : 
                         (N113)? mem[1211] : 
                         (N115)? mem[1275] : 
                         (N117)? mem[1339] : 
                         (N119)? mem[1403] : 
                         (N121)? mem[1467] : 
                         (N123)? mem[1531] : 
                         (N125)? mem[1595] : 
                         (N127)? mem[1659] : 
                         (N129)? mem[1723] : 
                         (N131)? mem[1787] : 
                         (N133)? mem[1851] : 
                         (N135)? mem[1915] : 
                         (N137)? mem[1979] : 
                         (N139)? mem[2043] : 1'b0;
  assign r1_data_o[58] = (N108)? mem[58] : 
                         (N110)? mem[122] : 
                         (N112)? mem[186] : 
                         (N114)? mem[250] : 
                         (N116)? mem[314] : 
                         (N118)? mem[378] : 
                         (N120)? mem[442] : 
                         (N122)? mem[506] : 
                         (N124)? mem[570] : 
                         (N126)? mem[634] : 
                         (N128)? mem[698] : 
                         (N130)? mem[762] : 
                         (N132)? mem[826] : 
                         (N134)? mem[890] : 
                         (N136)? mem[954] : 
                         (N138)? mem[1018] : 
                         (N109)? mem[1082] : 
                         (N111)? mem[1146] : 
                         (N113)? mem[1210] : 
                         (N115)? mem[1274] : 
                         (N117)? mem[1338] : 
                         (N119)? mem[1402] : 
                         (N121)? mem[1466] : 
                         (N123)? mem[1530] : 
                         (N125)? mem[1594] : 
                         (N127)? mem[1658] : 
                         (N129)? mem[1722] : 
                         (N131)? mem[1786] : 
                         (N133)? mem[1850] : 
                         (N135)? mem[1914] : 
                         (N137)? mem[1978] : 
                         (N139)? mem[2042] : 1'b0;
  assign r1_data_o[57] = (N108)? mem[57] : 
                         (N110)? mem[121] : 
                         (N112)? mem[185] : 
                         (N114)? mem[249] : 
                         (N116)? mem[313] : 
                         (N118)? mem[377] : 
                         (N120)? mem[441] : 
                         (N122)? mem[505] : 
                         (N124)? mem[569] : 
                         (N126)? mem[633] : 
                         (N128)? mem[697] : 
                         (N130)? mem[761] : 
                         (N132)? mem[825] : 
                         (N134)? mem[889] : 
                         (N136)? mem[953] : 
                         (N138)? mem[1017] : 
                         (N109)? mem[1081] : 
                         (N111)? mem[1145] : 
                         (N113)? mem[1209] : 
                         (N115)? mem[1273] : 
                         (N117)? mem[1337] : 
                         (N119)? mem[1401] : 
                         (N121)? mem[1465] : 
                         (N123)? mem[1529] : 
                         (N125)? mem[1593] : 
                         (N127)? mem[1657] : 
                         (N129)? mem[1721] : 
                         (N131)? mem[1785] : 
                         (N133)? mem[1849] : 
                         (N135)? mem[1913] : 
                         (N137)? mem[1977] : 
                         (N139)? mem[2041] : 1'b0;
  assign r1_data_o[56] = (N108)? mem[56] : 
                         (N110)? mem[120] : 
                         (N112)? mem[184] : 
                         (N114)? mem[248] : 
                         (N116)? mem[312] : 
                         (N118)? mem[376] : 
                         (N120)? mem[440] : 
                         (N122)? mem[504] : 
                         (N124)? mem[568] : 
                         (N126)? mem[632] : 
                         (N128)? mem[696] : 
                         (N130)? mem[760] : 
                         (N132)? mem[824] : 
                         (N134)? mem[888] : 
                         (N136)? mem[952] : 
                         (N138)? mem[1016] : 
                         (N109)? mem[1080] : 
                         (N111)? mem[1144] : 
                         (N113)? mem[1208] : 
                         (N115)? mem[1272] : 
                         (N117)? mem[1336] : 
                         (N119)? mem[1400] : 
                         (N121)? mem[1464] : 
                         (N123)? mem[1528] : 
                         (N125)? mem[1592] : 
                         (N127)? mem[1656] : 
                         (N129)? mem[1720] : 
                         (N131)? mem[1784] : 
                         (N133)? mem[1848] : 
                         (N135)? mem[1912] : 
                         (N137)? mem[1976] : 
                         (N139)? mem[2040] : 1'b0;
  assign r1_data_o[55] = (N108)? mem[55] : 
                         (N110)? mem[119] : 
                         (N112)? mem[183] : 
                         (N114)? mem[247] : 
                         (N116)? mem[311] : 
                         (N118)? mem[375] : 
                         (N120)? mem[439] : 
                         (N122)? mem[503] : 
                         (N124)? mem[567] : 
                         (N126)? mem[631] : 
                         (N128)? mem[695] : 
                         (N130)? mem[759] : 
                         (N132)? mem[823] : 
                         (N134)? mem[887] : 
                         (N136)? mem[951] : 
                         (N138)? mem[1015] : 
                         (N109)? mem[1079] : 
                         (N111)? mem[1143] : 
                         (N113)? mem[1207] : 
                         (N115)? mem[1271] : 
                         (N117)? mem[1335] : 
                         (N119)? mem[1399] : 
                         (N121)? mem[1463] : 
                         (N123)? mem[1527] : 
                         (N125)? mem[1591] : 
                         (N127)? mem[1655] : 
                         (N129)? mem[1719] : 
                         (N131)? mem[1783] : 
                         (N133)? mem[1847] : 
                         (N135)? mem[1911] : 
                         (N137)? mem[1975] : 
                         (N139)? mem[2039] : 1'b0;
  assign r1_data_o[54] = (N108)? mem[54] : 
                         (N110)? mem[118] : 
                         (N112)? mem[182] : 
                         (N114)? mem[246] : 
                         (N116)? mem[310] : 
                         (N118)? mem[374] : 
                         (N120)? mem[438] : 
                         (N122)? mem[502] : 
                         (N124)? mem[566] : 
                         (N126)? mem[630] : 
                         (N128)? mem[694] : 
                         (N130)? mem[758] : 
                         (N132)? mem[822] : 
                         (N134)? mem[886] : 
                         (N136)? mem[950] : 
                         (N138)? mem[1014] : 
                         (N109)? mem[1078] : 
                         (N111)? mem[1142] : 
                         (N113)? mem[1206] : 
                         (N115)? mem[1270] : 
                         (N117)? mem[1334] : 
                         (N119)? mem[1398] : 
                         (N121)? mem[1462] : 
                         (N123)? mem[1526] : 
                         (N125)? mem[1590] : 
                         (N127)? mem[1654] : 
                         (N129)? mem[1718] : 
                         (N131)? mem[1782] : 
                         (N133)? mem[1846] : 
                         (N135)? mem[1910] : 
                         (N137)? mem[1974] : 
                         (N139)? mem[2038] : 1'b0;
  assign r1_data_o[53] = (N108)? mem[53] : 
                         (N110)? mem[117] : 
                         (N112)? mem[181] : 
                         (N114)? mem[245] : 
                         (N116)? mem[309] : 
                         (N118)? mem[373] : 
                         (N120)? mem[437] : 
                         (N122)? mem[501] : 
                         (N124)? mem[565] : 
                         (N126)? mem[629] : 
                         (N128)? mem[693] : 
                         (N130)? mem[757] : 
                         (N132)? mem[821] : 
                         (N134)? mem[885] : 
                         (N136)? mem[949] : 
                         (N138)? mem[1013] : 
                         (N109)? mem[1077] : 
                         (N111)? mem[1141] : 
                         (N113)? mem[1205] : 
                         (N115)? mem[1269] : 
                         (N117)? mem[1333] : 
                         (N119)? mem[1397] : 
                         (N121)? mem[1461] : 
                         (N123)? mem[1525] : 
                         (N125)? mem[1589] : 
                         (N127)? mem[1653] : 
                         (N129)? mem[1717] : 
                         (N131)? mem[1781] : 
                         (N133)? mem[1845] : 
                         (N135)? mem[1909] : 
                         (N137)? mem[1973] : 
                         (N139)? mem[2037] : 1'b0;
  assign r1_data_o[52] = (N108)? mem[52] : 
                         (N110)? mem[116] : 
                         (N112)? mem[180] : 
                         (N114)? mem[244] : 
                         (N116)? mem[308] : 
                         (N118)? mem[372] : 
                         (N120)? mem[436] : 
                         (N122)? mem[500] : 
                         (N124)? mem[564] : 
                         (N126)? mem[628] : 
                         (N128)? mem[692] : 
                         (N130)? mem[756] : 
                         (N132)? mem[820] : 
                         (N134)? mem[884] : 
                         (N136)? mem[948] : 
                         (N138)? mem[1012] : 
                         (N109)? mem[1076] : 
                         (N111)? mem[1140] : 
                         (N113)? mem[1204] : 
                         (N115)? mem[1268] : 
                         (N117)? mem[1332] : 
                         (N119)? mem[1396] : 
                         (N121)? mem[1460] : 
                         (N123)? mem[1524] : 
                         (N125)? mem[1588] : 
                         (N127)? mem[1652] : 
                         (N129)? mem[1716] : 
                         (N131)? mem[1780] : 
                         (N133)? mem[1844] : 
                         (N135)? mem[1908] : 
                         (N137)? mem[1972] : 
                         (N139)? mem[2036] : 1'b0;
  assign r1_data_o[51] = (N108)? mem[51] : 
                         (N110)? mem[115] : 
                         (N112)? mem[179] : 
                         (N114)? mem[243] : 
                         (N116)? mem[307] : 
                         (N118)? mem[371] : 
                         (N120)? mem[435] : 
                         (N122)? mem[499] : 
                         (N124)? mem[563] : 
                         (N126)? mem[627] : 
                         (N128)? mem[691] : 
                         (N130)? mem[755] : 
                         (N132)? mem[819] : 
                         (N134)? mem[883] : 
                         (N136)? mem[947] : 
                         (N138)? mem[1011] : 
                         (N109)? mem[1075] : 
                         (N111)? mem[1139] : 
                         (N113)? mem[1203] : 
                         (N115)? mem[1267] : 
                         (N117)? mem[1331] : 
                         (N119)? mem[1395] : 
                         (N121)? mem[1459] : 
                         (N123)? mem[1523] : 
                         (N125)? mem[1587] : 
                         (N127)? mem[1651] : 
                         (N129)? mem[1715] : 
                         (N131)? mem[1779] : 
                         (N133)? mem[1843] : 
                         (N135)? mem[1907] : 
                         (N137)? mem[1971] : 
                         (N139)? mem[2035] : 1'b0;
  assign r1_data_o[50] = (N108)? mem[50] : 
                         (N110)? mem[114] : 
                         (N112)? mem[178] : 
                         (N114)? mem[242] : 
                         (N116)? mem[306] : 
                         (N118)? mem[370] : 
                         (N120)? mem[434] : 
                         (N122)? mem[498] : 
                         (N124)? mem[562] : 
                         (N126)? mem[626] : 
                         (N128)? mem[690] : 
                         (N130)? mem[754] : 
                         (N132)? mem[818] : 
                         (N134)? mem[882] : 
                         (N136)? mem[946] : 
                         (N138)? mem[1010] : 
                         (N109)? mem[1074] : 
                         (N111)? mem[1138] : 
                         (N113)? mem[1202] : 
                         (N115)? mem[1266] : 
                         (N117)? mem[1330] : 
                         (N119)? mem[1394] : 
                         (N121)? mem[1458] : 
                         (N123)? mem[1522] : 
                         (N125)? mem[1586] : 
                         (N127)? mem[1650] : 
                         (N129)? mem[1714] : 
                         (N131)? mem[1778] : 
                         (N133)? mem[1842] : 
                         (N135)? mem[1906] : 
                         (N137)? mem[1970] : 
                         (N139)? mem[2034] : 1'b0;
  assign r1_data_o[49] = (N108)? mem[49] : 
                         (N110)? mem[113] : 
                         (N112)? mem[177] : 
                         (N114)? mem[241] : 
                         (N116)? mem[305] : 
                         (N118)? mem[369] : 
                         (N120)? mem[433] : 
                         (N122)? mem[497] : 
                         (N124)? mem[561] : 
                         (N126)? mem[625] : 
                         (N128)? mem[689] : 
                         (N130)? mem[753] : 
                         (N132)? mem[817] : 
                         (N134)? mem[881] : 
                         (N136)? mem[945] : 
                         (N138)? mem[1009] : 
                         (N109)? mem[1073] : 
                         (N111)? mem[1137] : 
                         (N113)? mem[1201] : 
                         (N115)? mem[1265] : 
                         (N117)? mem[1329] : 
                         (N119)? mem[1393] : 
                         (N121)? mem[1457] : 
                         (N123)? mem[1521] : 
                         (N125)? mem[1585] : 
                         (N127)? mem[1649] : 
                         (N129)? mem[1713] : 
                         (N131)? mem[1777] : 
                         (N133)? mem[1841] : 
                         (N135)? mem[1905] : 
                         (N137)? mem[1969] : 
                         (N139)? mem[2033] : 1'b0;
  assign r1_data_o[48] = (N108)? mem[48] : 
                         (N110)? mem[112] : 
                         (N112)? mem[176] : 
                         (N114)? mem[240] : 
                         (N116)? mem[304] : 
                         (N118)? mem[368] : 
                         (N120)? mem[432] : 
                         (N122)? mem[496] : 
                         (N124)? mem[560] : 
                         (N126)? mem[624] : 
                         (N128)? mem[688] : 
                         (N130)? mem[752] : 
                         (N132)? mem[816] : 
                         (N134)? mem[880] : 
                         (N136)? mem[944] : 
                         (N138)? mem[1008] : 
                         (N109)? mem[1072] : 
                         (N111)? mem[1136] : 
                         (N113)? mem[1200] : 
                         (N115)? mem[1264] : 
                         (N117)? mem[1328] : 
                         (N119)? mem[1392] : 
                         (N121)? mem[1456] : 
                         (N123)? mem[1520] : 
                         (N125)? mem[1584] : 
                         (N127)? mem[1648] : 
                         (N129)? mem[1712] : 
                         (N131)? mem[1776] : 
                         (N133)? mem[1840] : 
                         (N135)? mem[1904] : 
                         (N137)? mem[1968] : 
                         (N139)? mem[2032] : 1'b0;
  assign r1_data_o[47] = (N108)? mem[47] : 
                         (N110)? mem[111] : 
                         (N112)? mem[175] : 
                         (N114)? mem[239] : 
                         (N116)? mem[303] : 
                         (N118)? mem[367] : 
                         (N120)? mem[431] : 
                         (N122)? mem[495] : 
                         (N124)? mem[559] : 
                         (N126)? mem[623] : 
                         (N128)? mem[687] : 
                         (N130)? mem[751] : 
                         (N132)? mem[815] : 
                         (N134)? mem[879] : 
                         (N136)? mem[943] : 
                         (N138)? mem[1007] : 
                         (N109)? mem[1071] : 
                         (N111)? mem[1135] : 
                         (N113)? mem[1199] : 
                         (N115)? mem[1263] : 
                         (N117)? mem[1327] : 
                         (N119)? mem[1391] : 
                         (N121)? mem[1455] : 
                         (N123)? mem[1519] : 
                         (N125)? mem[1583] : 
                         (N127)? mem[1647] : 
                         (N129)? mem[1711] : 
                         (N131)? mem[1775] : 
                         (N133)? mem[1839] : 
                         (N135)? mem[1903] : 
                         (N137)? mem[1967] : 
                         (N139)? mem[2031] : 1'b0;
  assign r1_data_o[46] = (N108)? mem[46] : 
                         (N110)? mem[110] : 
                         (N112)? mem[174] : 
                         (N114)? mem[238] : 
                         (N116)? mem[302] : 
                         (N118)? mem[366] : 
                         (N120)? mem[430] : 
                         (N122)? mem[494] : 
                         (N124)? mem[558] : 
                         (N126)? mem[622] : 
                         (N128)? mem[686] : 
                         (N130)? mem[750] : 
                         (N132)? mem[814] : 
                         (N134)? mem[878] : 
                         (N136)? mem[942] : 
                         (N138)? mem[1006] : 
                         (N109)? mem[1070] : 
                         (N111)? mem[1134] : 
                         (N113)? mem[1198] : 
                         (N115)? mem[1262] : 
                         (N117)? mem[1326] : 
                         (N119)? mem[1390] : 
                         (N121)? mem[1454] : 
                         (N123)? mem[1518] : 
                         (N125)? mem[1582] : 
                         (N127)? mem[1646] : 
                         (N129)? mem[1710] : 
                         (N131)? mem[1774] : 
                         (N133)? mem[1838] : 
                         (N135)? mem[1902] : 
                         (N137)? mem[1966] : 
                         (N139)? mem[2030] : 1'b0;
  assign r1_data_o[45] = (N108)? mem[45] : 
                         (N110)? mem[109] : 
                         (N112)? mem[173] : 
                         (N114)? mem[237] : 
                         (N116)? mem[301] : 
                         (N118)? mem[365] : 
                         (N120)? mem[429] : 
                         (N122)? mem[493] : 
                         (N124)? mem[557] : 
                         (N126)? mem[621] : 
                         (N128)? mem[685] : 
                         (N130)? mem[749] : 
                         (N132)? mem[813] : 
                         (N134)? mem[877] : 
                         (N136)? mem[941] : 
                         (N138)? mem[1005] : 
                         (N109)? mem[1069] : 
                         (N111)? mem[1133] : 
                         (N113)? mem[1197] : 
                         (N115)? mem[1261] : 
                         (N117)? mem[1325] : 
                         (N119)? mem[1389] : 
                         (N121)? mem[1453] : 
                         (N123)? mem[1517] : 
                         (N125)? mem[1581] : 
                         (N127)? mem[1645] : 
                         (N129)? mem[1709] : 
                         (N131)? mem[1773] : 
                         (N133)? mem[1837] : 
                         (N135)? mem[1901] : 
                         (N137)? mem[1965] : 
                         (N139)? mem[2029] : 1'b0;
  assign r1_data_o[44] = (N108)? mem[44] : 
                         (N110)? mem[108] : 
                         (N112)? mem[172] : 
                         (N114)? mem[236] : 
                         (N116)? mem[300] : 
                         (N118)? mem[364] : 
                         (N120)? mem[428] : 
                         (N122)? mem[492] : 
                         (N124)? mem[556] : 
                         (N126)? mem[620] : 
                         (N128)? mem[684] : 
                         (N130)? mem[748] : 
                         (N132)? mem[812] : 
                         (N134)? mem[876] : 
                         (N136)? mem[940] : 
                         (N138)? mem[1004] : 
                         (N109)? mem[1068] : 
                         (N111)? mem[1132] : 
                         (N113)? mem[1196] : 
                         (N115)? mem[1260] : 
                         (N117)? mem[1324] : 
                         (N119)? mem[1388] : 
                         (N121)? mem[1452] : 
                         (N123)? mem[1516] : 
                         (N125)? mem[1580] : 
                         (N127)? mem[1644] : 
                         (N129)? mem[1708] : 
                         (N131)? mem[1772] : 
                         (N133)? mem[1836] : 
                         (N135)? mem[1900] : 
                         (N137)? mem[1964] : 
                         (N139)? mem[2028] : 1'b0;
  assign r1_data_o[43] = (N108)? mem[43] : 
                         (N110)? mem[107] : 
                         (N112)? mem[171] : 
                         (N114)? mem[235] : 
                         (N116)? mem[299] : 
                         (N118)? mem[363] : 
                         (N120)? mem[427] : 
                         (N122)? mem[491] : 
                         (N124)? mem[555] : 
                         (N126)? mem[619] : 
                         (N128)? mem[683] : 
                         (N130)? mem[747] : 
                         (N132)? mem[811] : 
                         (N134)? mem[875] : 
                         (N136)? mem[939] : 
                         (N138)? mem[1003] : 
                         (N109)? mem[1067] : 
                         (N111)? mem[1131] : 
                         (N113)? mem[1195] : 
                         (N115)? mem[1259] : 
                         (N117)? mem[1323] : 
                         (N119)? mem[1387] : 
                         (N121)? mem[1451] : 
                         (N123)? mem[1515] : 
                         (N125)? mem[1579] : 
                         (N127)? mem[1643] : 
                         (N129)? mem[1707] : 
                         (N131)? mem[1771] : 
                         (N133)? mem[1835] : 
                         (N135)? mem[1899] : 
                         (N137)? mem[1963] : 
                         (N139)? mem[2027] : 1'b0;
  assign r1_data_o[42] = (N108)? mem[42] : 
                         (N110)? mem[106] : 
                         (N112)? mem[170] : 
                         (N114)? mem[234] : 
                         (N116)? mem[298] : 
                         (N118)? mem[362] : 
                         (N120)? mem[426] : 
                         (N122)? mem[490] : 
                         (N124)? mem[554] : 
                         (N126)? mem[618] : 
                         (N128)? mem[682] : 
                         (N130)? mem[746] : 
                         (N132)? mem[810] : 
                         (N134)? mem[874] : 
                         (N136)? mem[938] : 
                         (N138)? mem[1002] : 
                         (N109)? mem[1066] : 
                         (N111)? mem[1130] : 
                         (N113)? mem[1194] : 
                         (N115)? mem[1258] : 
                         (N117)? mem[1322] : 
                         (N119)? mem[1386] : 
                         (N121)? mem[1450] : 
                         (N123)? mem[1514] : 
                         (N125)? mem[1578] : 
                         (N127)? mem[1642] : 
                         (N129)? mem[1706] : 
                         (N131)? mem[1770] : 
                         (N133)? mem[1834] : 
                         (N135)? mem[1898] : 
                         (N137)? mem[1962] : 
                         (N139)? mem[2026] : 1'b0;
  assign r1_data_o[41] = (N108)? mem[41] : 
                         (N110)? mem[105] : 
                         (N112)? mem[169] : 
                         (N114)? mem[233] : 
                         (N116)? mem[297] : 
                         (N118)? mem[361] : 
                         (N120)? mem[425] : 
                         (N122)? mem[489] : 
                         (N124)? mem[553] : 
                         (N126)? mem[617] : 
                         (N128)? mem[681] : 
                         (N130)? mem[745] : 
                         (N132)? mem[809] : 
                         (N134)? mem[873] : 
                         (N136)? mem[937] : 
                         (N138)? mem[1001] : 
                         (N109)? mem[1065] : 
                         (N111)? mem[1129] : 
                         (N113)? mem[1193] : 
                         (N115)? mem[1257] : 
                         (N117)? mem[1321] : 
                         (N119)? mem[1385] : 
                         (N121)? mem[1449] : 
                         (N123)? mem[1513] : 
                         (N125)? mem[1577] : 
                         (N127)? mem[1641] : 
                         (N129)? mem[1705] : 
                         (N131)? mem[1769] : 
                         (N133)? mem[1833] : 
                         (N135)? mem[1897] : 
                         (N137)? mem[1961] : 
                         (N139)? mem[2025] : 1'b0;
  assign r1_data_o[40] = (N108)? mem[40] : 
                         (N110)? mem[104] : 
                         (N112)? mem[168] : 
                         (N114)? mem[232] : 
                         (N116)? mem[296] : 
                         (N118)? mem[360] : 
                         (N120)? mem[424] : 
                         (N122)? mem[488] : 
                         (N124)? mem[552] : 
                         (N126)? mem[616] : 
                         (N128)? mem[680] : 
                         (N130)? mem[744] : 
                         (N132)? mem[808] : 
                         (N134)? mem[872] : 
                         (N136)? mem[936] : 
                         (N138)? mem[1000] : 
                         (N109)? mem[1064] : 
                         (N111)? mem[1128] : 
                         (N113)? mem[1192] : 
                         (N115)? mem[1256] : 
                         (N117)? mem[1320] : 
                         (N119)? mem[1384] : 
                         (N121)? mem[1448] : 
                         (N123)? mem[1512] : 
                         (N125)? mem[1576] : 
                         (N127)? mem[1640] : 
                         (N129)? mem[1704] : 
                         (N131)? mem[1768] : 
                         (N133)? mem[1832] : 
                         (N135)? mem[1896] : 
                         (N137)? mem[1960] : 
                         (N139)? mem[2024] : 1'b0;
  assign r1_data_o[39] = (N108)? mem[39] : 
                         (N110)? mem[103] : 
                         (N112)? mem[167] : 
                         (N114)? mem[231] : 
                         (N116)? mem[295] : 
                         (N118)? mem[359] : 
                         (N120)? mem[423] : 
                         (N122)? mem[487] : 
                         (N124)? mem[551] : 
                         (N126)? mem[615] : 
                         (N128)? mem[679] : 
                         (N130)? mem[743] : 
                         (N132)? mem[807] : 
                         (N134)? mem[871] : 
                         (N136)? mem[935] : 
                         (N138)? mem[999] : 
                         (N109)? mem[1063] : 
                         (N111)? mem[1127] : 
                         (N113)? mem[1191] : 
                         (N115)? mem[1255] : 
                         (N117)? mem[1319] : 
                         (N119)? mem[1383] : 
                         (N121)? mem[1447] : 
                         (N123)? mem[1511] : 
                         (N125)? mem[1575] : 
                         (N127)? mem[1639] : 
                         (N129)? mem[1703] : 
                         (N131)? mem[1767] : 
                         (N133)? mem[1831] : 
                         (N135)? mem[1895] : 
                         (N137)? mem[1959] : 
                         (N139)? mem[2023] : 1'b0;
  assign r1_data_o[38] = (N108)? mem[38] : 
                         (N110)? mem[102] : 
                         (N112)? mem[166] : 
                         (N114)? mem[230] : 
                         (N116)? mem[294] : 
                         (N118)? mem[358] : 
                         (N120)? mem[422] : 
                         (N122)? mem[486] : 
                         (N124)? mem[550] : 
                         (N126)? mem[614] : 
                         (N128)? mem[678] : 
                         (N130)? mem[742] : 
                         (N132)? mem[806] : 
                         (N134)? mem[870] : 
                         (N136)? mem[934] : 
                         (N138)? mem[998] : 
                         (N109)? mem[1062] : 
                         (N111)? mem[1126] : 
                         (N113)? mem[1190] : 
                         (N115)? mem[1254] : 
                         (N117)? mem[1318] : 
                         (N119)? mem[1382] : 
                         (N121)? mem[1446] : 
                         (N123)? mem[1510] : 
                         (N125)? mem[1574] : 
                         (N127)? mem[1638] : 
                         (N129)? mem[1702] : 
                         (N131)? mem[1766] : 
                         (N133)? mem[1830] : 
                         (N135)? mem[1894] : 
                         (N137)? mem[1958] : 
                         (N139)? mem[2022] : 1'b0;
  assign r1_data_o[37] = (N108)? mem[37] : 
                         (N110)? mem[101] : 
                         (N112)? mem[165] : 
                         (N114)? mem[229] : 
                         (N116)? mem[293] : 
                         (N118)? mem[357] : 
                         (N120)? mem[421] : 
                         (N122)? mem[485] : 
                         (N124)? mem[549] : 
                         (N126)? mem[613] : 
                         (N128)? mem[677] : 
                         (N130)? mem[741] : 
                         (N132)? mem[805] : 
                         (N134)? mem[869] : 
                         (N136)? mem[933] : 
                         (N138)? mem[997] : 
                         (N109)? mem[1061] : 
                         (N111)? mem[1125] : 
                         (N113)? mem[1189] : 
                         (N115)? mem[1253] : 
                         (N117)? mem[1317] : 
                         (N119)? mem[1381] : 
                         (N121)? mem[1445] : 
                         (N123)? mem[1509] : 
                         (N125)? mem[1573] : 
                         (N127)? mem[1637] : 
                         (N129)? mem[1701] : 
                         (N131)? mem[1765] : 
                         (N133)? mem[1829] : 
                         (N135)? mem[1893] : 
                         (N137)? mem[1957] : 
                         (N139)? mem[2021] : 1'b0;
  assign r1_data_o[36] = (N108)? mem[36] : 
                         (N110)? mem[100] : 
                         (N112)? mem[164] : 
                         (N114)? mem[228] : 
                         (N116)? mem[292] : 
                         (N118)? mem[356] : 
                         (N120)? mem[420] : 
                         (N122)? mem[484] : 
                         (N124)? mem[548] : 
                         (N126)? mem[612] : 
                         (N128)? mem[676] : 
                         (N130)? mem[740] : 
                         (N132)? mem[804] : 
                         (N134)? mem[868] : 
                         (N136)? mem[932] : 
                         (N138)? mem[996] : 
                         (N109)? mem[1060] : 
                         (N111)? mem[1124] : 
                         (N113)? mem[1188] : 
                         (N115)? mem[1252] : 
                         (N117)? mem[1316] : 
                         (N119)? mem[1380] : 
                         (N121)? mem[1444] : 
                         (N123)? mem[1508] : 
                         (N125)? mem[1572] : 
                         (N127)? mem[1636] : 
                         (N129)? mem[1700] : 
                         (N131)? mem[1764] : 
                         (N133)? mem[1828] : 
                         (N135)? mem[1892] : 
                         (N137)? mem[1956] : 
                         (N139)? mem[2020] : 1'b0;
  assign r1_data_o[35] = (N108)? mem[35] : 
                         (N110)? mem[99] : 
                         (N112)? mem[163] : 
                         (N114)? mem[227] : 
                         (N116)? mem[291] : 
                         (N118)? mem[355] : 
                         (N120)? mem[419] : 
                         (N122)? mem[483] : 
                         (N124)? mem[547] : 
                         (N126)? mem[611] : 
                         (N128)? mem[675] : 
                         (N130)? mem[739] : 
                         (N132)? mem[803] : 
                         (N134)? mem[867] : 
                         (N136)? mem[931] : 
                         (N138)? mem[995] : 
                         (N109)? mem[1059] : 
                         (N111)? mem[1123] : 
                         (N113)? mem[1187] : 
                         (N115)? mem[1251] : 
                         (N117)? mem[1315] : 
                         (N119)? mem[1379] : 
                         (N121)? mem[1443] : 
                         (N123)? mem[1507] : 
                         (N125)? mem[1571] : 
                         (N127)? mem[1635] : 
                         (N129)? mem[1699] : 
                         (N131)? mem[1763] : 
                         (N133)? mem[1827] : 
                         (N135)? mem[1891] : 
                         (N137)? mem[1955] : 
                         (N139)? mem[2019] : 1'b0;
  assign r1_data_o[34] = (N108)? mem[34] : 
                         (N110)? mem[98] : 
                         (N112)? mem[162] : 
                         (N114)? mem[226] : 
                         (N116)? mem[290] : 
                         (N118)? mem[354] : 
                         (N120)? mem[418] : 
                         (N122)? mem[482] : 
                         (N124)? mem[546] : 
                         (N126)? mem[610] : 
                         (N128)? mem[674] : 
                         (N130)? mem[738] : 
                         (N132)? mem[802] : 
                         (N134)? mem[866] : 
                         (N136)? mem[930] : 
                         (N138)? mem[994] : 
                         (N109)? mem[1058] : 
                         (N111)? mem[1122] : 
                         (N113)? mem[1186] : 
                         (N115)? mem[1250] : 
                         (N117)? mem[1314] : 
                         (N119)? mem[1378] : 
                         (N121)? mem[1442] : 
                         (N123)? mem[1506] : 
                         (N125)? mem[1570] : 
                         (N127)? mem[1634] : 
                         (N129)? mem[1698] : 
                         (N131)? mem[1762] : 
                         (N133)? mem[1826] : 
                         (N135)? mem[1890] : 
                         (N137)? mem[1954] : 
                         (N139)? mem[2018] : 1'b0;
  assign r1_data_o[33] = (N108)? mem[33] : 
                         (N110)? mem[97] : 
                         (N112)? mem[161] : 
                         (N114)? mem[225] : 
                         (N116)? mem[289] : 
                         (N118)? mem[353] : 
                         (N120)? mem[417] : 
                         (N122)? mem[481] : 
                         (N124)? mem[545] : 
                         (N126)? mem[609] : 
                         (N128)? mem[673] : 
                         (N130)? mem[737] : 
                         (N132)? mem[801] : 
                         (N134)? mem[865] : 
                         (N136)? mem[929] : 
                         (N138)? mem[993] : 
                         (N109)? mem[1057] : 
                         (N111)? mem[1121] : 
                         (N113)? mem[1185] : 
                         (N115)? mem[1249] : 
                         (N117)? mem[1313] : 
                         (N119)? mem[1377] : 
                         (N121)? mem[1441] : 
                         (N123)? mem[1505] : 
                         (N125)? mem[1569] : 
                         (N127)? mem[1633] : 
                         (N129)? mem[1697] : 
                         (N131)? mem[1761] : 
                         (N133)? mem[1825] : 
                         (N135)? mem[1889] : 
                         (N137)? mem[1953] : 
                         (N139)? mem[2017] : 1'b0;
  assign r1_data_o[32] = (N108)? mem[32] : 
                         (N110)? mem[96] : 
                         (N112)? mem[160] : 
                         (N114)? mem[224] : 
                         (N116)? mem[288] : 
                         (N118)? mem[352] : 
                         (N120)? mem[416] : 
                         (N122)? mem[480] : 
                         (N124)? mem[544] : 
                         (N126)? mem[608] : 
                         (N128)? mem[672] : 
                         (N130)? mem[736] : 
                         (N132)? mem[800] : 
                         (N134)? mem[864] : 
                         (N136)? mem[928] : 
                         (N138)? mem[992] : 
                         (N109)? mem[1056] : 
                         (N111)? mem[1120] : 
                         (N113)? mem[1184] : 
                         (N115)? mem[1248] : 
                         (N117)? mem[1312] : 
                         (N119)? mem[1376] : 
                         (N121)? mem[1440] : 
                         (N123)? mem[1504] : 
                         (N125)? mem[1568] : 
                         (N127)? mem[1632] : 
                         (N129)? mem[1696] : 
                         (N131)? mem[1760] : 
                         (N133)? mem[1824] : 
                         (N135)? mem[1888] : 
                         (N137)? mem[1952] : 
                         (N139)? mem[2016] : 1'b0;
  assign r1_data_o[31] = (N108)? mem[31] : 
                         (N110)? mem[95] : 
                         (N112)? mem[159] : 
                         (N114)? mem[223] : 
                         (N116)? mem[287] : 
                         (N118)? mem[351] : 
                         (N120)? mem[415] : 
                         (N122)? mem[479] : 
                         (N124)? mem[543] : 
                         (N126)? mem[607] : 
                         (N128)? mem[671] : 
                         (N130)? mem[735] : 
                         (N132)? mem[799] : 
                         (N134)? mem[863] : 
                         (N136)? mem[927] : 
                         (N138)? mem[991] : 
                         (N109)? mem[1055] : 
                         (N111)? mem[1119] : 
                         (N113)? mem[1183] : 
                         (N115)? mem[1247] : 
                         (N117)? mem[1311] : 
                         (N119)? mem[1375] : 
                         (N121)? mem[1439] : 
                         (N123)? mem[1503] : 
                         (N125)? mem[1567] : 
                         (N127)? mem[1631] : 
                         (N129)? mem[1695] : 
                         (N131)? mem[1759] : 
                         (N133)? mem[1823] : 
                         (N135)? mem[1887] : 
                         (N137)? mem[1951] : 
                         (N139)? mem[2015] : 1'b0;
  assign r1_data_o[30] = (N108)? mem[30] : 
                         (N110)? mem[94] : 
                         (N112)? mem[158] : 
                         (N114)? mem[222] : 
                         (N116)? mem[286] : 
                         (N118)? mem[350] : 
                         (N120)? mem[414] : 
                         (N122)? mem[478] : 
                         (N124)? mem[542] : 
                         (N126)? mem[606] : 
                         (N128)? mem[670] : 
                         (N130)? mem[734] : 
                         (N132)? mem[798] : 
                         (N134)? mem[862] : 
                         (N136)? mem[926] : 
                         (N138)? mem[990] : 
                         (N109)? mem[1054] : 
                         (N111)? mem[1118] : 
                         (N113)? mem[1182] : 
                         (N115)? mem[1246] : 
                         (N117)? mem[1310] : 
                         (N119)? mem[1374] : 
                         (N121)? mem[1438] : 
                         (N123)? mem[1502] : 
                         (N125)? mem[1566] : 
                         (N127)? mem[1630] : 
                         (N129)? mem[1694] : 
                         (N131)? mem[1758] : 
                         (N133)? mem[1822] : 
                         (N135)? mem[1886] : 
                         (N137)? mem[1950] : 
                         (N139)? mem[2014] : 1'b0;
  assign r1_data_o[29] = (N108)? mem[29] : 
                         (N110)? mem[93] : 
                         (N112)? mem[157] : 
                         (N114)? mem[221] : 
                         (N116)? mem[285] : 
                         (N118)? mem[349] : 
                         (N120)? mem[413] : 
                         (N122)? mem[477] : 
                         (N124)? mem[541] : 
                         (N126)? mem[605] : 
                         (N128)? mem[669] : 
                         (N130)? mem[733] : 
                         (N132)? mem[797] : 
                         (N134)? mem[861] : 
                         (N136)? mem[925] : 
                         (N138)? mem[989] : 
                         (N109)? mem[1053] : 
                         (N111)? mem[1117] : 
                         (N113)? mem[1181] : 
                         (N115)? mem[1245] : 
                         (N117)? mem[1309] : 
                         (N119)? mem[1373] : 
                         (N121)? mem[1437] : 
                         (N123)? mem[1501] : 
                         (N125)? mem[1565] : 
                         (N127)? mem[1629] : 
                         (N129)? mem[1693] : 
                         (N131)? mem[1757] : 
                         (N133)? mem[1821] : 
                         (N135)? mem[1885] : 
                         (N137)? mem[1949] : 
                         (N139)? mem[2013] : 1'b0;
  assign r1_data_o[28] = (N108)? mem[28] : 
                         (N110)? mem[92] : 
                         (N112)? mem[156] : 
                         (N114)? mem[220] : 
                         (N116)? mem[284] : 
                         (N118)? mem[348] : 
                         (N120)? mem[412] : 
                         (N122)? mem[476] : 
                         (N124)? mem[540] : 
                         (N126)? mem[604] : 
                         (N128)? mem[668] : 
                         (N130)? mem[732] : 
                         (N132)? mem[796] : 
                         (N134)? mem[860] : 
                         (N136)? mem[924] : 
                         (N138)? mem[988] : 
                         (N109)? mem[1052] : 
                         (N111)? mem[1116] : 
                         (N113)? mem[1180] : 
                         (N115)? mem[1244] : 
                         (N117)? mem[1308] : 
                         (N119)? mem[1372] : 
                         (N121)? mem[1436] : 
                         (N123)? mem[1500] : 
                         (N125)? mem[1564] : 
                         (N127)? mem[1628] : 
                         (N129)? mem[1692] : 
                         (N131)? mem[1756] : 
                         (N133)? mem[1820] : 
                         (N135)? mem[1884] : 
                         (N137)? mem[1948] : 
                         (N139)? mem[2012] : 1'b0;
  assign r1_data_o[27] = (N108)? mem[27] : 
                         (N110)? mem[91] : 
                         (N112)? mem[155] : 
                         (N114)? mem[219] : 
                         (N116)? mem[283] : 
                         (N118)? mem[347] : 
                         (N120)? mem[411] : 
                         (N122)? mem[475] : 
                         (N124)? mem[539] : 
                         (N126)? mem[603] : 
                         (N128)? mem[667] : 
                         (N130)? mem[731] : 
                         (N132)? mem[795] : 
                         (N134)? mem[859] : 
                         (N136)? mem[923] : 
                         (N138)? mem[987] : 
                         (N109)? mem[1051] : 
                         (N111)? mem[1115] : 
                         (N113)? mem[1179] : 
                         (N115)? mem[1243] : 
                         (N117)? mem[1307] : 
                         (N119)? mem[1371] : 
                         (N121)? mem[1435] : 
                         (N123)? mem[1499] : 
                         (N125)? mem[1563] : 
                         (N127)? mem[1627] : 
                         (N129)? mem[1691] : 
                         (N131)? mem[1755] : 
                         (N133)? mem[1819] : 
                         (N135)? mem[1883] : 
                         (N137)? mem[1947] : 
                         (N139)? mem[2011] : 1'b0;
  assign r1_data_o[26] = (N108)? mem[26] : 
                         (N110)? mem[90] : 
                         (N112)? mem[154] : 
                         (N114)? mem[218] : 
                         (N116)? mem[282] : 
                         (N118)? mem[346] : 
                         (N120)? mem[410] : 
                         (N122)? mem[474] : 
                         (N124)? mem[538] : 
                         (N126)? mem[602] : 
                         (N128)? mem[666] : 
                         (N130)? mem[730] : 
                         (N132)? mem[794] : 
                         (N134)? mem[858] : 
                         (N136)? mem[922] : 
                         (N138)? mem[986] : 
                         (N109)? mem[1050] : 
                         (N111)? mem[1114] : 
                         (N113)? mem[1178] : 
                         (N115)? mem[1242] : 
                         (N117)? mem[1306] : 
                         (N119)? mem[1370] : 
                         (N121)? mem[1434] : 
                         (N123)? mem[1498] : 
                         (N125)? mem[1562] : 
                         (N127)? mem[1626] : 
                         (N129)? mem[1690] : 
                         (N131)? mem[1754] : 
                         (N133)? mem[1818] : 
                         (N135)? mem[1882] : 
                         (N137)? mem[1946] : 
                         (N139)? mem[2010] : 1'b0;
  assign r1_data_o[25] = (N108)? mem[25] : 
                         (N110)? mem[89] : 
                         (N112)? mem[153] : 
                         (N114)? mem[217] : 
                         (N116)? mem[281] : 
                         (N118)? mem[345] : 
                         (N120)? mem[409] : 
                         (N122)? mem[473] : 
                         (N124)? mem[537] : 
                         (N126)? mem[601] : 
                         (N128)? mem[665] : 
                         (N130)? mem[729] : 
                         (N132)? mem[793] : 
                         (N134)? mem[857] : 
                         (N136)? mem[921] : 
                         (N138)? mem[985] : 
                         (N109)? mem[1049] : 
                         (N111)? mem[1113] : 
                         (N113)? mem[1177] : 
                         (N115)? mem[1241] : 
                         (N117)? mem[1305] : 
                         (N119)? mem[1369] : 
                         (N121)? mem[1433] : 
                         (N123)? mem[1497] : 
                         (N125)? mem[1561] : 
                         (N127)? mem[1625] : 
                         (N129)? mem[1689] : 
                         (N131)? mem[1753] : 
                         (N133)? mem[1817] : 
                         (N135)? mem[1881] : 
                         (N137)? mem[1945] : 
                         (N139)? mem[2009] : 1'b0;
  assign r1_data_o[24] = (N108)? mem[24] : 
                         (N110)? mem[88] : 
                         (N112)? mem[152] : 
                         (N114)? mem[216] : 
                         (N116)? mem[280] : 
                         (N118)? mem[344] : 
                         (N120)? mem[408] : 
                         (N122)? mem[472] : 
                         (N124)? mem[536] : 
                         (N126)? mem[600] : 
                         (N128)? mem[664] : 
                         (N130)? mem[728] : 
                         (N132)? mem[792] : 
                         (N134)? mem[856] : 
                         (N136)? mem[920] : 
                         (N138)? mem[984] : 
                         (N109)? mem[1048] : 
                         (N111)? mem[1112] : 
                         (N113)? mem[1176] : 
                         (N115)? mem[1240] : 
                         (N117)? mem[1304] : 
                         (N119)? mem[1368] : 
                         (N121)? mem[1432] : 
                         (N123)? mem[1496] : 
                         (N125)? mem[1560] : 
                         (N127)? mem[1624] : 
                         (N129)? mem[1688] : 
                         (N131)? mem[1752] : 
                         (N133)? mem[1816] : 
                         (N135)? mem[1880] : 
                         (N137)? mem[1944] : 
                         (N139)? mem[2008] : 1'b0;
  assign r1_data_o[23] = (N108)? mem[23] : 
                         (N110)? mem[87] : 
                         (N112)? mem[151] : 
                         (N114)? mem[215] : 
                         (N116)? mem[279] : 
                         (N118)? mem[343] : 
                         (N120)? mem[407] : 
                         (N122)? mem[471] : 
                         (N124)? mem[535] : 
                         (N126)? mem[599] : 
                         (N128)? mem[663] : 
                         (N130)? mem[727] : 
                         (N132)? mem[791] : 
                         (N134)? mem[855] : 
                         (N136)? mem[919] : 
                         (N138)? mem[983] : 
                         (N109)? mem[1047] : 
                         (N111)? mem[1111] : 
                         (N113)? mem[1175] : 
                         (N115)? mem[1239] : 
                         (N117)? mem[1303] : 
                         (N119)? mem[1367] : 
                         (N121)? mem[1431] : 
                         (N123)? mem[1495] : 
                         (N125)? mem[1559] : 
                         (N127)? mem[1623] : 
                         (N129)? mem[1687] : 
                         (N131)? mem[1751] : 
                         (N133)? mem[1815] : 
                         (N135)? mem[1879] : 
                         (N137)? mem[1943] : 
                         (N139)? mem[2007] : 1'b0;
  assign r1_data_o[22] = (N108)? mem[22] : 
                         (N110)? mem[86] : 
                         (N112)? mem[150] : 
                         (N114)? mem[214] : 
                         (N116)? mem[278] : 
                         (N118)? mem[342] : 
                         (N120)? mem[406] : 
                         (N122)? mem[470] : 
                         (N124)? mem[534] : 
                         (N126)? mem[598] : 
                         (N128)? mem[662] : 
                         (N130)? mem[726] : 
                         (N132)? mem[790] : 
                         (N134)? mem[854] : 
                         (N136)? mem[918] : 
                         (N138)? mem[982] : 
                         (N109)? mem[1046] : 
                         (N111)? mem[1110] : 
                         (N113)? mem[1174] : 
                         (N115)? mem[1238] : 
                         (N117)? mem[1302] : 
                         (N119)? mem[1366] : 
                         (N121)? mem[1430] : 
                         (N123)? mem[1494] : 
                         (N125)? mem[1558] : 
                         (N127)? mem[1622] : 
                         (N129)? mem[1686] : 
                         (N131)? mem[1750] : 
                         (N133)? mem[1814] : 
                         (N135)? mem[1878] : 
                         (N137)? mem[1942] : 
                         (N139)? mem[2006] : 1'b0;
  assign r1_data_o[21] = (N108)? mem[21] : 
                         (N110)? mem[85] : 
                         (N112)? mem[149] : 
                         (N114)? mem[213] : 
                         (N116)? mem[277] : 
                         (N118)? mem[341] : 
                         (N120)? mem[405] : 
                         (N122)? mem[469] : 
                         (N124)? mem[533] : 
                         (N126)? mem[597] : 
                         (N128)? mem[661] : 
                         (N130)? mem[725] : 
                         (N132)? mem[789] : 
                         (N134)? mem[853] : 
                         (N136)? mem[917] : 
                         (N138)? mem[981] : 
                         (N109)? mem[1045] : 
                         (N111)? mem[1109] : 
                         (N113)? mem[1173] : 
                         (N115)? mem[1237] : 
                         (N117)? mem[1301] : 
                         (N119)? mem[1365] : 
                         (N121)? mem[1429] : 
                         (N123)? mem[1493] : 
                         (N125)? mem[1557] : 
                         (N127)? mem[1621] : 
                         (N129)? mem[1685] : 
                         (N131)? mem[1749] : 
                         (N133)? mem[1813] : 
                         (N135)? mem[1877] : 
                         (N137)? mem[1941] : 
                         (N139)? mem[2005] : 1'b0;
  assign r1_data_o[20] = (N108)? mem[20] : 
                         (N110)? mem[84] : 
                         (N112)? mem[148] : 
                         (N114)? mem[212] : 
                         (N116)? mem[276] : 
                         (N118)? mem[340] : 
                         (N120)? mem[404] : 
                         (N122)? mem[468] : 
                         (N124)? mem[532] : 
                         (N126)? mem[596] : 
                         (N128)? mem[660] : 
                         (N130)? mem[724] : 
                         (N132)? mem[788] : 
                         (N134)? mem[852] : 
                         (N136)? mem[916] : 
                         (N138)? mem[980] : 
                         (N109)? mem[1044] : 
                         (N111)? mem[1108] : 
                         (N113)? mem[1172] : 
                         (N115)? mem[1236] : 
                         (N117)? mem[1300] : 
                         (N119)? mem[1364] : 
                         (N121)? mem[1428] : 
                         (N123)? mem[1492] : 
                         (N125)? mem[1556] : 
                         (N127)? mem[1620] : 
                         (N129)? mem[1684] : 
                         (N131)? mem[1748] : 
                         (N133)? mem[1812] : 
                         (N135)? mem[1876] : 
                         (N137)? mem[1940] : 
                         (N139)? mem[2004] : 1'b0;
  assign r1_data_o[19] = (N108)? mem[19] : 
                         (N110)? mem[83] : 
                         (N112)? mem[147] : 
                         (N114)? mem[211] : 
                         (N116)? mem[275] : 
                         (N118)? mem[339] : 
                         (N120)? mem[403] : 
                         (N122)? mem[467] : 
                         (N124)? mem[531] : 
                         (N126)? mem[595] : 
                         (N128)? mem[659] : 
                         (N130)? mem[723] : 
                         (N132)? mem[787] : 
                         (N134)? mem[851] : 
                         (N136)? mem[915] : 
                         (N138)? mem[979] : 
                         (N109)? mem[1043] : 
                         (N111)? mem[1107] : 
                         (N113)? mem[1171] : 
                         (N115)? mem[1235] : 
                         (N117)? mem[1299] : 
                         (N119)? mem[1363] : 
                         (N121)? mem[1427] : 
                         (N123)? mem[1491] : 
                         (N125)? mem[1555] : 
                         (N127)? mem[1619] : 
                         (N129)? mem[1683] : 
                         (N131)? mem[1747] : 
                         (N133)? mem[1811] : 
                         (N135)? mem[1875] : 
                         (N137)? mem[1939] : 
                         (N139)? mem[2003] : 1'b0;
  assign r1_data_o[18] = (N108)? mem[18] : 
                         (N110)? mem[82] : 
                         (N112)? mem[146] : 
                         (N114)? mem[210] : 
                         (N116)? mem[274] : 
                         (N118)? mem[338] : 
                         (N120)? mem[402] : 
                         (N122)? mem[466] : 
                         (N124)? mem[530] : 
                         (N126)? mem[594] : 
                         (N128)? mem[658] : 
                         (N130)? mem[722] : 
                         (N132)? mem[786] : 
                         (N134)? mem[850] : 
                         (N136)? mem[914] : 
                         (N138)? mem[978] : 
                         (N109)? mem[1042] : 
                         (N111)? mem[1106] : 
                         (N113)? mem[1170] : 
                         (N115)? mem[1234] : 
                         (N117)? mem[1298] : 
                         (N119)? mem[1362] : 
                         (N121)? mem[1426] : 
                         (N123)? mem[1490] : 
                         (N125)? mem[1554] : 
                         (N127)? mem[1618] : 
                         (N129)? mem[1682] : 
                         (N131)? mem[1746] : 
                         (N133)? mem[1810] : 
                         (N135)? mem[1874] : 
                         (N137)? mem[1938] : 
                         (N139)? mem[2002] : 1'b0;
  assign r1_data_o[17] = (N108)? mem[17] : 
                         (N110)? mem[81] : 
                         (N112)? mem[145] : 
                         (N114)? mem[209] : 
                         (N116)? mem[273] : 
                         (N118)? mem[337] : 
                         (N120)? mem[401] : 
                         (N122)? mem[465] : 
                         (N124)? mem[529] : 
                         (N126)? mem[593] : 
                         (N128)? mem[657] : 
                         (N130)? mem[721] : 
                         (N132)? mem[785] : 
                         (N134)? mem[849] : 
                         (N136)? mem[913] : 
                         (N138)? mem[977] : 
                         (N109)? mem[1041] : 
                         (N111)? mem[1105] : 
                         (N113)? mem[1169] : 
                         (N115)? mem[1233] : 
                         (N117)? mem[1297] : 
                         (N119)? mem[1361] : 
                         (N121)? mem[1425] : 
                         (N123)? mem[1489] : 
                         (N125)? mem[1553] : 
                         (N127)? mem[1617] : 
                         (N129)? mem[1681] : 
                         (N131)? mem[1745] : 
                         (N133)? mem[1809] : 
                         (N135)? mem[1873] : 
                         (N137)? mem[1937] : 
                         (N139)? mem[2001] : 1'b0;
  assign r1_data_o[16] = (N108)? mem[16] : 
                         (N110)? mem[80] : 
                         (N112)? mem[144] : 
                         (N114)? mem[208] : 
                         (N116)? mem[272] : 
                         (N118)? mem[336] : 
                         (N120)? mem[400] : 
                         (N122)? mem[464] : 
                         (N124)? mem[528] : 
                         (N126)? mem[592] : 
                         (N128)? mem[656] : 
                         (N130)? mem[720] : 
                         (N132)? mem[784] : 
                         (N134)? mem[848] : 
                         (N136)? mem[912] : 
                         (N138)? mem[976] : 
                         (N109)? mem[1040] : 
                         (N111)? mem[1104] : 
                         (N113)? mem[1168] : 
                         (N115)? mem[1232] : 
                         (N117)? mem[1296] : 
                         (N119)? mem[1360] : 
                         (N121)? mem[1424] : 
                         (N123)? mem[1488] : 
                         (N125)? mem[1552] : 
                         (N127)? mem[1616] : 
                         (N129)? mem[1680] : 
                         (N131)? mem[1744] : 
                         (N133)? mem[1808] : 
                         (N135)? mem[1872] : 
                         (N137)? mem[1936] : 
                         (N139)? mem[2000] : 1'b0;
  assign r1_data_o[15] = (N108)? mem[15] : 
                         (N110)? mem[79] : 
                         (N112)? mem[143] : 
                         (N114)? mem[207] : 
                         (N116)? mem[271] : 
                         (N118)? mem[335] : 
                         (N120)? mem[399] : 
                         (N122)? mem[463] : 
                         (N124)? mem[527] : 
                         (N126)? mem[591] : 
                         (N128)? mem[655] : 
                         (N130)? mem[719] : 
                         (N132)? mem[783] : 
                         (N134)? mem[847] : 
                         (N136)? mem[911] : 
                         (N138)? mem[975] : 
                         (N109)? mem[1039] : 
                         (N111)? mem[1103] : 
                         (N113)? mem[1167] : 
                         (N115)? mem[1231] : 
                         (N117)? mem[1295] : 
                         (N119)? mem[1359] : 
                         (N121)? mem[1423] : 
                         (N123)? mem[1487] : 
                         (N125)? mem[1551] : 
                         (N127)? mem[1615] : 
                         (N129)? mem[1679] : 
                         (N131)? mem[1743] : 
                         (N133)? mem[1807] : 
                         (N135)? mem[1871] : 
                         (N137)? mem[1935] : 
                         (N139)? mem[1999] : 1'b0;
  assign r1_data_o[14] = (N108)? mem[14] : 
                         (N110)? mem[78] : 
                         (N112)? mem[142] : 
                         (N114)? mem[206] : 
                         (N116)? mem[270] : 
                         (N118)? mem[334] : 
                         (N120)? mem[398] : 
                         (N122)? mem[462] : 
                         (N124)? mem[526] : 
                         (N126)? mem[590] : 
                         (N128)? mem[654] : 
                         (N130)? mem[718] : 
                         (N132)? mem[782] : 
                         (N134)? mem[846] : 
                         (N136)? mem[910] : 
                         (N138)? mem[974] : 
                         (N109)? mem[1038] : 
                         (N111)? mem[1102] : 
                         (N113)? mem[1166] : 
                         (N115)? mem[1230] : 
                         (N117)? mem[1294] : 
                         (N119)? mem[1358] : 
                         (N121)? mem[1422] : 
                         (N123)? mem[1486] : 
                         (N125)? mem[1550] : 
                         (N127)? mem[1614] : 
                         (N129)? mem[1678] : 
                         (N131)? mem[1742] : 
                         (N133)? mem[1806] : 
                         (N135)? mem[1870] : 
                         (N137)? mem[1934] : 
                         (N139)? mem[1998] : 1'b0;
  assign r1_data_o[13] = (N108)? mem[13] : 
                         (N110)? mem[77] : 
                         (N112)? mem[141] : 
                         (N114)? mem[205] : 
                         (N116)? mem[269] : 
                         (N118)? mem[333] : 
                         (N120)? mem[397] : 
                         (N122)? mem[461] : 
                         (N124)? mem[525] : 
                         (N126)? mem[589] : 
                         (N128)? mem[653] : 
                         (N130)? mem[717] : 
                         (N132)? mem[781] : 
                         (N134)? mem[845] : 
                         (N136)? mem[909] : 
                         (N138)? mem[973] : 
                         (N109)? mem[1037] : 
                         (N111)? mem[1101] : 
                         (N113)? mem[1165] : 
                         (N115)? mem[1229] : 
                         (N117)? mem[1293] : 
                         (N119)? mem[1357] : 
                         (N121)? mem[1421] : 
                         (N123)? mem[1485] : 
                         (N125)? mem[1549] : 
                         (N127)? mem[1613] : 
                         (N129)? mem[1677] : 
                         (N131)? mem[1741] : 
                         (N133)? mem[1805] : 
                         (N135)? mem[1869] : 
                         (N137)? mem[1933] : 
                         (N139)? mem[1997] : 1'b0;
  assign r1_data_o[12] = (N108)? mem[12] : 
                         (N110)? mem[76] : 
                         (N112)? mem[140] : 
                         (N114)? mem[204] : 
                         (N116)? mem[268] : 
                         (N118)? mem[332] : 
                         (N120)? mem[396] : 
                         (N122)? mem[460] : 
                         (N124)? mem[524] : 
                         (N126)? mem[588] : 
                         (N128)? mem[652] : 
                         (N130)? mem[716] : 
                         (N132)? mem[780] : 
                         (N134)? mem[844] : 
                         (N136)? mem[908] : 
                         (N138)? mem[972] : 
                         (N109)? mem[1036] : 
                         (N111)? mem[1100] : 
                         (N113)? mem[1164] : 
                         (N115)? mem[1228] : 
                         (N117)? mem[1292] : 
                         (N119)? mem[1356] : 
                         (N121)? mem[1420] : 
                         (N123)? mem[1484] : 
                         (N125)? mem[1548] : 
                         (N127)? mem[1612] : 
                         (N129)? mem[1676] : 
                         (N131)? mem[1740] : 
                         (N133)? mem[1804] : 
                         (N135)? mem[1868] : 
                         (N137)? mem[1932] : 
                         (N139)? mem[1996] : 1'b0;
  assign r1_data_o[11] = (N108)? mem[11] : 
                         (N110)? mem[75] : 
                         (N112)? mem[139] : 
                         (N114)? mem[203] : 
                         (N116)? mem[267] : 
                         (N118)? mem[331] : 
                         (N120)? mem[395] : 
                         (N122)? mem[459] : 
                         (N124)? mem[523] : 
                         (N126)? mem[587] : 
                         (N128)? mem[651] : 
                         (N130)? mem[715] : 
                         (N132)? mem[779] : 
                         (N134)? mem[843] : 
                         (N136)? mem[907] : 
                         (N138)? mem[971] : 
                         (N109)? mem[1035] : 
                         (N111)? mem[1099] : 
                         (N113)? mem[1163] : 
                         (N115)? mem[1227] : 
                         (N117)? mem[1291] : 
                         (N119)? mem[1355] : 
                         (N121)? mem[1419] : 
                         (N123)? mem[1483] : 
                         (N125)? mem[1547] : 
                         (N127)? mem[1611] : 
                         (N129)? mem[1675] : 
                         (N131)? mem[1739] : 
                         (N133)? mem[1803] : 
                         (N135)? mem[1867] : 
                         (N137)? mem[1931] : 
                         (N139)? mem[1995] : 1'b0;
  assign r1_data_o[10] = (N108)? mem[10] : 
                         (N110)? mem[74] : 
                         (N112)? mem[138] : 
                         (N114)? mem[202] : 
                         (N116)? mem[266] : 
                         (N118)? mem[330] : 
                         (N120)? mem[394] : 
                         (N122)? mem[458] : 
                         (N124)? mem[522] : 
                         (N126)? mem[586] : 
                         (N128)? mem[650] : 
                         (N130)? mem[714] : 
                         (N132)? mem[778] : 
                         (N134)? mem[842] : 
                         (N136)? mem[906] : 
                         (N138)? mem[970] : 
                         (N109)? mem[1034] : 
                         (N111)? mem[1098] : 
                         (N113)? mem[1162] : 
                         (N115)? mem[1226] : 
                         (N117)? mem[1290] : 
                         (N119)? mem[1354] : 
                         (N121)? mem[1418] : 
                         (N123)? mem[1482] : 
                         (N125)? mem[1546] : 
                         (N127)? mem[1610] : 
                         (N129)? mem[1674] : 
                         (N131)? mem[1738] : 
                         (N133)? mem[1802] : 
                         (N135)? mem[1866] : 
                         (N137)? mem[1930] : 
                         (N139)? mem[1994] : 1'b0;
  assign r1_data_o[9] = (N108)? mem[9] : 
                        (N110)? mem[73] : 
                        (N112)? mem[137] : 
                        (N114)? mem[201] : 
                        (N116)? mem[265] : 
                        (N118)? mem[329] : 
                        (N120)? mem[393] : 
                        (N122)? mem[457] : 
                        (N124)? mem[521] : 
                        (N126)? mem[585] : 
                        (N128)? mem[649] : 
                        (N130)? mem[713] : 
                        (N132)? mem[777] : 
                        (N134)? mem[841] : 
                        (N136)? mem[905] : 
                        (N138)? mem[969] : 
                        (N109)? mem[1033] : 
                        (N111)? mem[1097] : 
                        (N113)? mem[1161] : 
                        (N115)? mem[1225] : 
                        (N117)? mem[1289] : 
                        (N119)? mem[1353] : 
                        (N121)? mem[1417] : 
                        (N123)? mem[1481] : 
                        (N125)? mem[1545] : 
                        (N127)? mem[1609] : 
                        (N129)? mem[1673] : 
                        (N131)? mem[1737] : 
                        (N133)? mem[1801] : 
                        (N135)? mem[1865] : 
                        (N137)? mem[1929] : 
                        (N139)? mem[1993] : 1'b0;
  assign r1_data_o[8] = (N108)? mem[8] : 
                        (N110)? mem[72] : 
                        (N112)? mem[136] : 
                        (N114)? mem[200] : 
                        (N116)? mem[264] : 
                        (N118)? mem[328] : 
                        (N120)? mem[392] : 
                        (N122)? mem[456] : 
                        (N124)? mem[520] : 
                        (N126)? mem[584] : 
                        (N128)? mem[648] : 
                        (N130)? mem[712] : 
                        (N132)? mem[776] : 
                        (N134)? mem[840] : 
                        (N136)? mem[904] : 
                        (N138)? mem[968] : 
                        (N109)? mem[1032] : 
                        (N111)? mem[1096] : 
                        (N113)? mem[1160] : 
                        (N115)? mem[1224] : 
                        (N117)? mem[1288] : 
                        (N119)? mem[1352] : 
                        (N121)? mem[1416] : 
                        (N123)? mem[1480] : 
                        (N125)? mem[1544] : 
                        (N127)? mem[1608] : 
                        (N129)? mem[1672] : 
                        (N131)? mem[1736] : 
                        (N133)? mem[1800] : 
                        (N135)? mem[1864] : 
                        (N137)? mem[1928] : 
                        (N139)? mem[1992] : 1'b0;
  assign r1_data_o[7] = (N108)? mem[7] : 
                        (N110)? mem[71] : 
                        (N112)? mem[135] : 
                        (N114)? mem[199] : 
                        (N116)? mem[263] : 
                        (N118)? mem[327] : 
                        (N120)? mem[391] : 
                        (N122)? mem[455] : 
                        (N124)? mem[519] : 
                        (N126)? mem[583] : 
                        (N128)? mem[647] : 
                        (N130)? mem[711] : 
                        (N132)? mem[775] : 
                        (N134)? mem[839] : 
                        (N136)? mem[903] : 
                        (N138)? mem[967] : 
                        (N109)? mem[1031] : 
                        (N111)? mem[1095] : 
                        (N113)? mem[1159] : 
                        (N115)? mem[1223] : 
                        (N117)? mem[1287] : 
                        (N119)? mem[1351] : 
                        (N121)? mem[1415] : 
                        (N123)? mem[1479] : 
                        (N125)? mem[1543] : 
                        (N127)? mem[1607] : 
                        (N129)? mem[1671] : 
                        (N131)? mem[1735] : 
                        (N133)? mem[1799] : 
                        (N135)? mem[1863] : 
                        (N137)? mem[1927] : 
                        (N139)? mem[1991] : 1'b0;
  assign r1_data_o[6] = (N108)? mem[6] : 
                        (N110)? mem[70] : 
                        (N112)? mem[134] : 
                        (N114)? mem[198] : 
                        (N116)? mem[262] : 
                        (N118)? mem[326] : 
                        (N120)? mem[390] : 
                        (N122)? mem[454] : 
                        (N124)? mem[518] : 
                        (N126)? mem[582] : 
                        (N128)? mem[646] : 
                        (N130)? mem[710] : 
                        (N132)? mem[774] : 
                        (N134)? mem[838] : 
                        (N136)? mem[902] : 
                        (N138)? mem[966] : 
                        (N109)? mem[1030] : 
                        (N111)? mem[1094] : 
                        (N113)? mem[1158] : 
                        (N115)? mem[1222] : 
                        (N117)? mem[1286] : 
                        (N119)? mem[1350] : 
                        (N121)? mem[1414] : 
                        (N123)? mem[1478] : 
                        (N125)? mem[1542] : 
                        (N127)? mem[1606] : 
                        (N129)? mem[1670] : 
                        (N131)? mem[1734] : 
                        (N133)? mem[1798] : 
                        (N135)? mem[1862] : 
                        (N137)? mem[1926] : 
                        (N139)? mem[1990] : 1'b0;
  assign r1_data_o[5] = (N108)? mem[5] : 
                        (N110)? mem[69] : 
                        (N112)? mem[133] : 
                        (N114)? mem[197] : 
                        (N116)? mem[261] : 
                        (N118)? mem[325] : 
                        (N120)? mem[389] : 
                        (N122)? mem[453] : 
                        (N124)? mem[517] : 
                        (N126)? mem[581] : 
                        (N128)? mem[645] : 
                        (N130)? mem[709] : 
                        (N132)? mem[773] : 
                        (N134)? mem[837] : 
                        (N136)? mem[901] : 
                        (N138)? mem[965] : 
                        (N109)? mem[1029] : 
                        (N111)? mem[1093] : 
                        (N113)? mem[1157] : 
                        (N115)? mem[1221] : 
                        (N117)? mem[1285] : 
                        (N119)? mem[1349] : 
                        (N121)? mem[1413] : 
                        (N123)? mem[1477] : 
                        (N125)? mem[1541] : 
                        (N127)? mem[1605] : 
                        (N129)? mem[1669] : 
                        (N131)? mem[1733] : 
                        (N133)? mem[1797] : 
                        (N135)? mem[1861] : 
                        (N137)? mem[1925] : 
                        (N139)? mem[1989] : 1'b0;
  assign r1_data_o[4] = (N108)? mem[4] : 
                        (N110)? mem[68] : 
                        (N112)? mem[132] : 
                        (N114)? mem[196] : 
                        (N116)? mem[260] : 
                        (N118)? mem[324] : 
                        (N120)? mem[388] : 
                        (N122)? mem[452] : 
                        (N124)? mem[516] : 
                        (N126)? mem[580] : 
                        (N128)? mem[644] : 
                        (N130)? mem[708] : 
                        (N132)? mem[772] : 
                        (N134)? mem[836] : 
                        (N136)? mem[900] : 
                        (N138)? mem[964] : 
                        (N109)? mem[1028] : 
                        (N111)? mem[1092] : 
                        (N113)? mem[1156] : 
                        (N115)? mem[1220] : 
                        (N117)? mem[1284] : 
                        (N119)? mem[1348] : 
                        (N121)? mem[1412] : 
                        (N123)? mem[1476] : 
                        (N125)? mem[1540] : 
                        (N127)? mem[1604] : 
                        (N129)? mem[1668] : 
                        (N131)? mem[1732] : 
                        (N133)? mem[1796] : 
                        (N135)? mem[1860] : 
                        (N137)? mem[1924] : 
                        (N139)? mem[1988] : 1'b0;
  assign r1_data_o[3] = (N108)? mem[3] : 
                        (N110)? mem[67] : 
                        (N112)? mem[131] : 
                        (N114)? mem[195] : 
                        (N116)? mem[259] : 
                        (N118)? mem[323] : 
                        (N120)? mem[387] : 
                        (N122)? mem[451] : 
                        (N124)? mem[515] : 
                        (N126)? mem[579] : 
                        (N128)? mem[643] : 
                        (N130)? mem[707] : 
                        (N132)? mem[771] : 
                        (N134)? mem[835] : 
                        (N136)? mem[899] : 
                        (N138)? mem[963] : 
                        (N109)? mem[1027] : 
                        (N111)? mem[1091] : 
                        (N113)? mem[1155] : 
                        (N115)? mem[1219] : 
                        (N117)? mem[1283] : 
                        (N119)? mem[1347] : 
                        (N121)? mem[1411] : 
                        (N123)? mem[1475] : 
                        (N125)? mem[1539] : 
                        (N127)? mem[1603] : 
                        (N129)? mem[1667] : 
                        (N131)? mem[1731] : 
                        (N133)? mem[1795] : 
                        (N135)? mem[1859] : 
                        (N137)? mem[1923] : 
                        (N139)? mem[1987] : 1'b0;
  assign r1_data_o[2] = (N108)? mem[2] : 
                        (N110)? mem[66] : 
                        (N112)? mem[130] : 
                        (N114)? mem[194] : 
                        (N116)? mem[258] : 
                        (N118)? mem[322] : 
                        (N120)? mem[386] : 
                        (N122)? mem[450] : 
                        (N124)? mem[514] : 
                        (N126)? mem[578] : 
                        (N128)? mem[642] : 
                        (N130)? mem[706] : 
                        (N132)? mem[770] : 
                        (N134)? mem[834] : 
                        (N136)? mem[898] : 
                        (N138)? mem[962] : 
                        (N109)? mem[1026] : 
                        (N111)? mem[1090] : 
                        (N113)? mem[1154] : 
                        (N115)? mem[1218] : 
                        (N117)? mem[1282] : 
                        (N119)? mem[1346] : 
                        (N121)? mem[1410] : 
                        (N123)? mem[1474] : 
                        (N125)? mem[1538] : 
                        (N127)? mem[1602] : 
                        (N129)? mem[1666] : 
                        (N131)? mem[1730] : 
                        (N133)? mem[1794] : 
                        (N135)? mem[1858] : 
                        (N137)? mem[1922] : 
                        (N139)? mem[1986] : 1'b0;
  assign r1_data_o[1] = (N108)? mem[1] : 
                        (N110)? mem[65] : 
                        (N112)? mem[129] : 
                        (N114)? mem[193] : 
                        (N116)? mem[257] : 
                        (N118)? mem[321] : 
                        (N120)? mem[385] : 
                        (N122)? mem[449] : 
                        (N124)? mem[513] : 
                        (N126)? mem[577] : 
                        (N128)? mem[641] : 
                        (N130)? mem[705] : 
                        (N132)? mem[769] : 
                        (N134)? mem[833] : 
                        (N136)? mem[897] : 
                        (N138)? mem[961] : 
                        (N109)? mem[1025] : 
                        (N111)? mem[1089] : 
                        (N113)? mem[1153] : 
                        (N115)? mem[1217] : 
                        (N117)? mem[1281] : 
                        (N119)? mem[1345] : 
                        (N121)? mem[1409] : 
                        (N123)? mem[1473] : 
                        (N125)? mem[1537] : 
                        (N127)? mem[1601] : 
                        (N129)? mem[1665] : 
                        (N131)? mem[1729] : 
                        (N133)? mem[1793] : 
                        (N135)? mem[1857] : 
                        (N137)? mem[1921] : 
                        (N139)? mem[1985] : 1'b0;
  assign r1_data_o[0] = (N108)? mem[0] : 
                        (N110)? mem[64] : 
                        (N112)? mem[128] : 
                        (N114)? mem[192] : 
                        (N116)? mem[256] : 
                        (N118)? mem[320] : 
                        (N120)? mem[384] : 
                        (N122)? mem[448] : 
                        (N124)? mem[512] : 
                        (N126)? mem[576] : 
                        (N128)? mem[640] : 
                        (N130)? mem[704] : 
                        (N132)? mem[768] : 
                        (N134)? mem[832] : 
                        (N136)? mem[896] : 
                        (N138)? mem[960] : 
                        (N109)? mem[1024] : 
                        (N111)? mem[1088] : 
                        (N113)? mem[1152] : 
                        (N115)? mem[1216] : 
                        (N117)? mem[1280] : 
                        (N119)? mem[1344] : 
                        (N121)? mem[1408] : 
                        (N123)? mem[1472] : 
                        (N125)? mem[1536] : 
                        (N127)? mem[1600] : 
                        (N129)? mem[1664] : 
                        (N131)? mem[1728] : 
                        (N133)? mem[1792] : 
                        (N135)? mem[1856] : 
                        (N137)? mem[1920] : 
                        (N139)? mem[1984] : 1'b0;
  assign N205 = w_addr_i[3] & w_addr_i[4];
  assign N206 = N0 & w_addr_i[4];
  assign N0 = ~w_addr_i[3];
  assign N207 = w_addr_i[3] & N1;
  assign N1 = ~w_addr_i[4];
  assign N208 = N2 & N3;
  assign N2 = ~w_addr_i[3];
  assign N3 = ~w_addr_i[4];
  assign N209 = ~w_addr_i[2];
  assign N210 = w_addr_i[0] & w_addr_i[1];
  assign N211 = N4 & w_addr_i[1];
  assign N4 = ~w_addr_i[0];
  assign N212 = w_addr_i[0] & N5;
  assign N5 = ~w_addr_i[1];
  assign N213 = N6 & N7;
  assign N6 = ~w_addr_i[0];
  assign N7 = ~w_addr_i[1];
  assign N214 = w_addr_i[2] & N210;
  assign N215 = w_addr_i[2] & N211;
  assign N216 = w_addr_i[2] & N212;
  assign N217 = w_addr_i[2] & N213;
  assign N218 = N209 & N210;
  assign N219 = N209 & N211;
  assign N220 = N209 & N212;
  assign N221 = N209 & N213;
  assign N172 = N205 & N214;
  assign N171 = N205 & N215;
  assign N170 = N205 & N216;
  assign N169 = N205 & N217;
  assign N168 = N205 & N218;
  assign N167 = N205 & N219;
  assign N166 = N205 & N220;
  assign N165 = N205 & N221;
  assign N164 = N206 & N214;
  assign N163 = N206 & N215;
  assign N162 = N206 & N216;
  assign N161 = N206 & N217;
  assign N160 = N206 & N218;
  assign N159 = N206 & N219;
  assign N158 = N206 & N220;
  assign N157 = N206 & N221;
  assign N156 = N207 & N214;
  assign N155 = N207 & N215;
  assign N154 = N207 & N216;
  assign N153 = N207 & N217;
  assign N152 = N207 & N218;
  assign N151 = N207 & N219;
  assign N150 = N207 & N220;
  assign N149 = N207 & N221;
  assign N148 = N208 & N214;
  assign N147 = N208 & N215;
  assign N146 = N208 & N216;
  assign N145 = N208 & N217;
  assign N144 = N208 & N218;
  assign N143 = N208 & N219;
  assign N142 = N208 & N220;
  assign N141 = N208 & N221;
  assign { N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173 } = (N8)? { N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141 } : 
                                                                                                                                                                                                              (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N140;
  assign N10 = ~r0_addr_r[0];
  assign N11 = ~r0_addr_r[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r0_addr_r[1];
  assign N14 = r0_addr_r[0] & N11;
  assign N15 = r0_addr_r[0] & r0_addr_r[1];
  assign N16 = ~r0_addr_r[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r0_addr_r[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r0_addr_r[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r0_addr_r[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r0_addr_r[2];
  assign N25 = ~r0_addr_r[3];
  assign N26 = N17 & N25;
  assign N27 = N17 & r0_addr_r[3];
  assign N28 = N19 & N25;
  assign N29 = N19 & r0_addr_r[3];
  assign N30 = N21 & N25;
  assign N31 = N21 & r0_addr_r[3];
  assign N32 = N23 & N25;
  assign N33 = N23 & r0_addr_r[3];
  assign N34 = N18 & N25;
  assign N35 = N18 & r0_addr_r[3];
  assign N36 = N20 & N25;
  assign N37 = N20 & r0_addr_r[3];
  assign N38 = N22 & N25;
  assign N39 = N22 & r0_addr_r[3];
  assign N40 = N24 & N25;
  assign N41 = N24 & r0_addr_r[3];
  assign N42 = ~r0_addr_r[4];
  assign N43 = N26 & N42;
  assign N44 = N26 & r0_addr_r[4];
  assign N45 = N28 & N42;
  assign N46 = N28 & r0_addr_r[4];
  assign N47 = N30 & N42;
  assign N48 = N30 & r0_addr_r[4];
  assign N49 = N32 & N42;
  assign N50 = N32 & r0_addr_r[4];
  assign N51 = N34 & N42;
  assign N52 = N34 & r0_addr_r[4];
  assign N53 = N36 & N42;
  assign N54 = N36 & r0_addr_r[4];
  assign N55 = N38 & N42;
  assign N56 = N38 & r0_addr_r[4];
  assign N57 = N40 & N42;
  assign N58 = N40 & r0_addr_r[4];
  assign N59 = N27 & N42;
  assign N60 = N27 & r0_addr_r[4];
  assign N61 = N29 & N42;
  assign N62 = N29 & r0_addr_r[4];
  assign N63 = N31 & N42;
  assign N64 = N31 & r0_addr_r[4];
  assign N65 = N33 & N42;
  assign N66 = N33 & r0_addr_r[4];
  assign N67 = N35 & N42;
  assign N68 = N35 & r0_addr_r[4];
  assign N69 = N37 & N42;
  assign N70 = N37 & r0_addr_r[4];
  assign N71 = N39 & N42;
  assign N72 = N39 & r0_addr_r[4];
  assign N73 = N41 & N42;
  assign N74 = N41 & r0_addr_r[4];
  assign N75 = ~r1_addr_r[0];
  assign N76 = ~r1_addr_r[1];
  assign N77 = N75 & N76;
  assign N78 = N75 & r1_addr_r[1];
  assign N79 = r1_addr_r[0] & N76;
  assign N80 = r1_addr_r[0] & r1_addr_r[1];
  assign N81 = ~r1_addr_r[2];
  assign N82 = N77 & N81;
  assign N83 = N77 & r1_addr_r[2];
  assign N84 = N79 & N81;
  assign N85 = N79 & r1_addr_r[2];
  assign N86 = N78 & N81;
  assign N87 = N78 & r1_addr_r[2];
  assign N88 = N80 & N81;
  assign N89 = N80 & r1_addr_r[2];
  assign N90 = ~r1_addr_r[3];
  assign N91 = N82 & N90;
  assign N92 = N82 & r1_addr_r[3];
  assign N93 = N84 & N90;
  assign N94 = N84 & r1_addr_r[3];
  assign N95 = N86 & N90;
  assign N96 = N86 & r1_addr_r[3];
  assign N97 = N88 & N90;
  assign N98 = N88 & r1_addr_r[3];
  assign N99 = N83 & N90;
  assign N100 = N83 & r1_addr_r[3];
  assign N101 = N85 & N90;
  assign N102 = N85 & r1_addr_r[3];
  assign N103 = N87 & N90;
  assign N104 = N87 & r1_addr_r[3];
  assign N105 = N89 & N90;
  assign N106 = N89 & r1_addr_r[3];
  assign N107 = ~r1_addr_r[4];
  assign N108 = N91 & N107;
  assign N109 = N91 & r1_addr_r[4];
  assign N110 = N93 & N107;
  assign N111 = N93 & r1_addr_r[4];
  assign N112 = N95 & N107;
  assign N113 = N95 & r1_addr_r[4];
  assign N114 = N97 & N107;
  assign N115 = N97 & r1_addr_r[4];
  assign N116 = N99 & N107;
  assign N117 = N99 & r1_addr_r[4];
  assign N118 = N101 & N107;
  assign N119 = N101 & r1_addr_r[4];
  assign N120 = N103 & N107;
  assign N121 = N103 & r1_addr_r[4];
  assign N122 = N105 & N107;
  assign N123 = N105 & r1_addr_r[4];
  assign N124 = N92 & N107;
  assign N125 = N92 & r1_addr_r[4];
  assign N126 = N94 & N107;
  assign N127 = N94 & r1_addr_r[4];
  assign N128 = N96 & N107;
  assign N129 = N96 & r1_addr_r[4];
  assign N130 = N98 & N107;
  assign N131 = N98 & r1_addr_r[4];
  assign N132 = N100 & N107;
  assign N133 = N100 & r1_addr_r[4];
  assign N134 = N102 & N107;
  assign N135 = N102 & r1_addr_r[4];
  assign N136 = N104 & N107;
  assign N137 = N104 & r1_addr_r[4];
  assign N138 = N106 & N107;
  assign N139 = N106 & r1_addr_r[4];
  assign N140 = ~w_v_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { r0_addr_r[4:0] } <= { r0_addr_i[4:0] };
      { r1_addr_r[4:0] } <= { r1_addr_i[4:0] };
    end 
    if(N204) begin
      { mem[2047:1984] } <= { w_data_i[63:0] };
    end 
    if(N203) begin
      { mem[1983:1920] } <= { w_data_i[63:0] };
    end 
    if(N202) begin
      { mem[1919:1856] } <= { w_data_i[63:0] };
    end 
    if(N201) begin
      { mem[1855:1792] } <= { w_data_i[63:0] };
    end 
    if(N200) begin
      { mem[1791:1728] } <= { w_data_i[63:0] };
    end 
    if(N199) begin
      { mem[1727:1664] } <= { w_data_i[63:0] };
    end 
    if(N198) begin
      { mem[1663:1600] } <= { w_data_i[63:0] };
    end 
    if(N197) begin
      { mem[1599:1536] } <= { w_data_i[63:0] };
    end 
    if(N196) begin
      { mem[1535:1472] } <= { w_data_i[63:0] };
    end 
    if(N195) begin
      { mem[1471:1408] } <= { w_data_i[63:0] };
    end 
    if(N194) begin
      { mem[1407:1344] } <= { w_data_i[63:0] };
    end 
    if(N193) begin
      { mem[1343:1280] } <= { w_data_i[63:0] };
    end 
    if(N192) begin
      { mem[1279:1216] } <= { w_data_i[63:0] };
    end 
    if(N191) begin
      { mem[1215:1152] } <= { w_data_i[63:0] };
    end 
    if(N190) begin
      { mem[1151:1088] } <= { w_data_i[63:0] };
    end 
    if(N189) begin
      { mem[1087:1024] } <= { w_data_i[63:0] };
    end 
    if(N188) begin
      { mem[1023:960] } <= { w_data_i[63:0] };
    end 
    if(N187) begin
      { mem[959:896] } <= { w_data_i[63:0] };
    end 
    if(N186) begin
      { mem[895:832] } <= { w_data_i[63:0] };
    end 
    if(N185) begin
      { mem[831:768] } <= { w_data_i[63:0] };
    end 
    if(N184) begin
      { mem[767:704] } <= { w_data_i[63:0] };
    end 
    if(N183) begin
      { mem[703:640] } <= { w_data_i[63:0] };
    end 
    if(N182) begin
      { mem[639:576] } <= { w_data_i[63:0] };
    end 
    if(N181) begin
      { mem[575:512] } <= { w_data_i[63:0] };
    end 
    if(N180) begin
      { mem[511:448] } <= { w_data_i[63:0] };
    end 
    if(N179) begin
      { mem[447:384] } <= { w_data_i[63:0] };
    end 
    if(N178) begin
      { mem[383:320] } <= { w_data_i[63:0] };
    end 
    if(N177) begin
      { mem[319:256] } <= { w_data_i[63:0] };
    end 
    if(N176) begin
      { mem[255:192] } <= { w_data_i[63:0] };
    end 
    if(N175) begin
      { mem[191:128] } <= { w_data_i[63:0] };
    end 
    if(N174) begin
      { mem[127:64] } <= { w_data_i[63:0] };
    end 
    if(N173) begin
      { mem[63:0] } <= { w_data_i[63:0] };
    end 
  end


endmodule