module bsg_dff_reset_width_p65_harden_p0
(
  clock_i,
  data_i,
  reset_i,
  data_o
);

  input [64:0] data_i;
  output [64:0] data_o;
  input clock_i;
  input reset_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67;
  reg [64:0] data_o;

  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[64] <= N67;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[63] <= N66;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[62] <= N65;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[61] <= N64;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[60] <= N63;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[59] <= N62;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[58] <= N61;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[57] <= N60;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[56] <= N59;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[55] <= N58;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[54] <= N57;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[53] <= N56;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[52] <= N55;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[51] <= N54;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[50] <= N53;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[49] <= N52;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[48] <= N51;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[47] <= N50;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[46] <= N49;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[45] <= N48;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[44] <= N47;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[43] <= N46;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[42] <= N45;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[41] <= N44;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[40] <= N43;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[39] <= N42;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[38] <= N41;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[37] <= N40;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[36] <= N39;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[35] <= N38;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[34] <= N37;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[33] <= N36;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[32] <= N35;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[31] <= N34;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[30] <= N33;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[29] <= N32;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[28] <= N31;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[27] <= N30;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[26] <= N29;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[25] <= N28;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[24] <= N27;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[23] <= N26;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[22] <= N25;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[21] <= N24;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[20] <= N23;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[19] <= N22;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[18] <= N21;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[17] <= N20;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[16] <= N19;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[15] <= N18;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[14] <= N17;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[13] <= N16;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[12] <= N15;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[11] <= N14;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[10] <= N13;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[9] <= N12;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[8] <= N11;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[7] <= N10;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[6] <= N9;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[5] <= N8;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[4] <= N7;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[3] <= N6;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[2] <= N5;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[1] <= N4;
    end 
  end


  always @(posedge clock_i) begin
    if(1'b1) begin
      data_o[0] <= N3;
    end 
  end

  assign { N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4, N3 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                            (N1)? data_i : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign N2 = ~reset_i;

endmodule