module bsg_mux_one_hot_width_p62_els_p4
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [247:0] data_i;
  input [3:0] sel_one_hot_i;
  output [61:0] data_o;
  wire [61:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123;
  wire [247:0] data_masked;
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[1];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[1];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[1];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[1];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[1];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[1];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[1];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[1];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[1];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[1];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[1];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[1];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[1];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[1];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[1];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[1];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[1];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[1];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[1];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[1];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[1];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[1];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[1];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[1];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[1];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[1];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[1];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[1];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[1];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[1];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[1];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[1];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[1];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[1];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[1];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[1];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[1];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[1];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[1];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[1];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[1];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[1];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[1];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[1];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[1];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[1];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[1];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[1];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[1];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[1];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[1];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[1];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[1];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[1];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[1];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[1];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[1];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[1];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[1];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[1];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[1];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[2];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[2];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[2];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[2];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[2];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[2];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[2];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[2];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[2];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[2];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[2];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[2];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[2];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[2];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[2];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[2];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[2];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[2];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[2];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[2];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[2];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[2];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[2];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[2];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[2];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[2];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[2];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[2];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[2];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[2];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[2];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[2];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[2];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[2];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[2];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[2];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[2];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[2];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[2];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[2];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[2];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[2];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[2];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[2];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[2];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[2];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[2];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[2];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[2];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[2];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[2];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[2];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[2];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[2];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[2];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[2];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[2];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[2];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[2];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[2];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[2];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[2];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[3];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[3];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[3];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[3];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[3];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[3];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[3];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[3];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[3];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[3];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[3];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[3];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[3];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[3];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[3];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[3];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[3];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[3];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[3];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[3];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[3];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[3];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[3];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[3];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[3];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[3];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[3];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[3];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[3];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[3];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[3];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[3];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[3];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[3];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[3];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[3];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[3];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[3];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[3];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[3];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[3];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[3];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[3];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[3];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[3];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[3];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[3];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[3];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[3];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[3];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[3];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[3];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[3];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[3];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[3];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[3];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[3];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[3];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[3];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[3];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[3];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[3];
  assign data_o[0] = N1 | data_masked[0];
  assign N1 = N0 | data_masked[62];
  assign N0 = data_masked[186] | data_masked[124];
  assign data_o[1] = N3 | data_masked[1];
  assign N3 = N2 | data_masked[63];
  assign N2 = data_masked[187] | data_masked[125];
  assign data_o[2] = N5 | data_masked[2];
  assign N5 = N4 | data_masked[64];
  assign N4 = data_masked[188] | data_masked[126];
  assign data_o[3] = N7 | data_masked[3];
  assign N7 = N6 | data_masked[65];
  assign N6 = data_masked[189] | data_masked[127];
  assign data_o[4] = N9 | data_masked[4];
  assign N9 = N8 | data_masked[66];
  assign N8 = data_masked[190] | data_masked[128];
  assign data_o[5] = N11 | data_masked[5];
  assign N11 = N10 | data_masked[67];
  assign N10 = data_masked[191] | data_masked[129];
  assign data_o[6] = N13 | data_masked[6];
  assign N13 = N12 | data_masked[68];
  assign N12 = data_masked[192] | data_masked[130];
  assign data_o[7] = N15 | data_masked[7];
  assign N15 = N14 | data_masked[69];
  assign N14 = data_masked[193] | data_masked[131];
  assign data_o[8] = N17 | data_masked[8];
  assign N17 = N16 | data_masked[70];
  assign N16 = data_masked[194] | data_masked[132];
  assign data_o[9] = N19 | data_masked[9];
  assign N19 = N18 | data_masked[71];
  assign N18 = data_masked[195] | data_masked[133];
  assign data_o[10] = N21 | data_masked[10];
  assign N21 = N20 | data_masked[72];
  assign N20 = data_masked[196] | data_masked[134];
  assign data_o[11] = N23 | data_masked[11];
  assign N23 = N22 | data_masked[73];
  assign N22 = data_masked[197] | data_masked[135];
  assign data_o[12] = N25 | data_masked[12];
  assign N25 = N24 | data_masked[74];
  assign N24 = data_masked[198] | data_masked[136];
  assign data_o[13] = N27 | data_masked[13];
  assign N27 = N26 | data_masked[75];
  assign N26 = data_masked[199] | data_masked[137];
  assign data_o[14] = N29 | data_masked[14];
  assign N29 = N28 | data_masked[76];
  assign N28 = data_masked[200] | data_masked[138];
  assign data_o[15] = N31 | data_masked[15];
  assign N31 = N30 | data_masked[77];
  assign N30 = data_masked[201] | data_masked[139];
  assign data_o[16] = N33 | data_masked[16];
  assign N33 = N32 | data_masked[78];
  assign N32 = data_masked[202] | data_masked[140];
  assign data_o[17] = N35 | data_masked[17];
  assign N35 = N34 | data_masked[79];
  assign N34 = data_masked[203] | data_masked[141];
  assign data_o[18] = N37 | data_masked[18];
  assign N37 = N36 | data_masked[80];
  assign N36 = data_masked[204] | data_masked[142];
  assign data_o[19] = N39 | data_masked[19];
  assign N39 = N38 | data_masked[81];
  assign N38 = data_masked[205] | data_masked[143];
  assign data_o[20] = N41 | data_masked[20];
  assign N41 = N40 | data_masked[82];
  assign N40 = data_masked[206] | data_masked[144];
  assign data_o[21] = N43 | data_masked[21];
  assign N43 = N42 | data_masked[83];
  assign N42 = data_masked[207] | data_masked[145];
  assign data_o[22] = N45 | data_masked[22];
  assign N45 = N44 | data_masked[84];
  assign N44 = data_masked[208] | data_masked[146];
  assign data_o[23] = N47 | data_masked[23];
  assign N47 = N46 | data_masked[85];
  assign N46 = data_masked[209] | data_masked[147];
  assign data_o[24] = N49 | data_masked[24];
  assign N49 = N48 | data_masked[86];
  assign N48 = data_masked[210] | data_masked[148];
  assign data_o[25] = N51 | data_masked[25];
  assign N51 = N50 | data_masked[87];
  assign N50 = data_masked[211] | data_masked[149];
  assign data_o[26] = N53 | data_masked[26];
  assign N53 = N52 | data_masked[88];
  assign N52 = data_masked[212] | data_masked[150];
  assign data_o[27] = N55 | data_masked[27];
  assign N55 = N54 | data_masked[89];
  assign N54 = data_masked[213] | data_masked[151];
  assign data_o[28] = N57 | data_masked[28];
  assign N57 = N56 | data_masked[90];
  assign N56 = data_masked[214] | data_masked[152];
  assign data_o[29] = N59 | data_masked[29];
  assign N59 = N58 | data_masked[91];
  assign N58 = data_masked[215] | data_masked[153];
  assign data_o[30] = N61 | data_masked[30];
  assign N61 = N60 | data_masked[92];
  assign N60 = data_masked[216] | data_masked[154];
  assign data_o[31] = N63 | data_masked[31];
  assign N63 = N62 | data_masked[93];
  assign N62 = data_masked[217] | data_masked[155];
  assign data_o[32] = N65 | data_masked[32];
  assign N65 = N64 | data_masked[94];
  assign N64 = data_masked[218] | data_masked[156];
  assign data_o[33] = N67 | data_masked[33];
  assign N67 = N66 | data_masked[95];
  assign N66 = data_masked[219] | data_masked[157];
  assign data_o[34] = N69 | data_masked[34];
  assign N69 = N68 | data_masked[96];
  assign N68 = data_masked[220] | data_masked[158];
  assign data_o[35] = N71 | data_masked[35];
  assign N71 = N70 | data_masked[97];
  assign N70 = data_masked[221] | data_masked[159];
  assign data_o[36] = N73 | data_masked[36];
  assign N73 = N72 | data_masked[98];
  assign N72 = data_masked[222] | data_masked[160];
  assign data_o[37] = N75 | data_masked[37];
  assign N75 = N74 | data_masked[99];
  assign N74 = data_masked[223] | data_masked[161];
  assign data_o[38] = N77 | data_masked[38];
  assign N77 = N76 | data_masked[100];
  assign N76 = data_masked[224] | data_masked[162];
  assign data_o[39] = N79 | data_masked[39];
  assign N79 = N78 | data_masked[101];
  assign N78 = data_masked[225] | data_masked[163];
  assign data_o[40] = N81 | data_masked[40];
  assign N81 = N80 | data_masked[102];
  assign N80 = data_masked[226] | data_masked[164];
  assign data_o[41] = N83 | data_masked[41];
  assign N83 = N82 | data_masked[103];
  assign N82 = data_masked[227] | data_masked[165];
  assign data_o[42] = N85 | data_masked[42];
  assign N85 = N84 | data_masked[104];
  assign N84 = data_masked[228] | data_masked[166];
  assign data_o[43] = N87 | data_masked[43];
  assign N87 = N86 | data_masked[105];
  assign N86 = data_masked[229] | data_masked[167];
  assign data_o[44] = N89 | data_masked[44];
  assign N89 = N88 | data_masked[106];
  assign N88 = data_masked[230] | data_masked[168];
  assign data_o[45] = N91 | data_masked[45];
  assign N91 = N90 | data_masked[107];
  assign N90 = data_masked[231] | data_masked[169];
  assign data_o[46] = N93 | data_masked[46];
  assign N93 = N92 | data_masked[108];
  assign N92 = data_masked[232] | data_masked[170];
  assign data_o[47] = N95 | data_masked[47];
  assign N95 = N94 | data_masked[109];
  assign N94 = data_masked[233] | data_masked[171];
  assign data_o[48] = N97 | data_masked[48];
  assign N97 = N96 | data_masked[110];
  assign N96 = data_masked[234] | data_masked[172];
  assign data_o[49] = N99 | data_masked[49];
  assign N99 = N98 | data_masked[111];
  assign N98 = data_masked[235] | data_masked[173];
  assign data_o[50] = N101 | data_masked[50];
  assign N101 = N100 | data_masked[112];
  assign N100 = data_masked[236] | data_masked[174];
  assign data_o[51] = N103 | data_masked[51];
  assign N103 = N102 | data_masked[113];
  assign N102 = data_masked[237] | data_masked[175];
  assign data_o[52] = N105 | data_masked[52];
  assign N105 = N104 | data_masked[114];
  assign N104 = data_masked[238] | data_masked[176];
  assign data_o[53] = N107 | data_masked[53];
  assign N107 = N106 | data_masked[115];
  assign N106 = data_masked[239] | data_masked[177];
  assign data_o[54] = N109 | data_masked[54];
  assign N109 = N108 | data_masked[116];
  assign N108 = data_masked[240] | data_masked[178];
  assign data_o[55] = N111 | data_masked[55];
  assign N111 = N110 | data_masked[117];
  assign N110 = data_masked[241] | data_masked[179];
  assign data_o[56] = N113 | data_masked[56];
  assign N113 = N112 | data_masked[118];
  assign N112 = data_masked[242] | data_masked[180];
  assign data_o[57] = N115 | data_masked[57];
  assign N115 = N114 | data_masked[119];
  assign N114 = data_masked[243] | data_masked[181];
  assign data_o[58] = N117 | data_masked[58];
  assign N117 = N116 | data_masked[120];
  assign N116 = data_masked[244] | data_masked[182];
  assign data_o[59] = N119 | data_masked[59];
  assign N119 = N118 | data_masked[121];
  assign N118 = data_masked[245] | data_masked[183];
  assign data_o[60] = N121 | data_masked[60];
  assign N121 = N120 | data_masked[122];
  assign N120 = data_masked[246] | data_masked[184];
  assign data_o[61] = N123 | data_masked[61];
  assign N123 = N122 | data_masked[123];
  assign N122 = data_masked[247] | data_masked[185];

endmodule