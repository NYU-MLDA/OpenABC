module ALU( // @[:freechips.rocketchip.system.TinyConfig.fir@123304.2]
  input  [3:0]  io_fn, // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
  input  [31:0] io_in2, // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
  input  [31:0] io_in1, // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
  output [31:0] io_out, // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
  output [31:0] io_adder_out, // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
  output        io_cmp_out // @[:freechips.rocketchip.system.TinyConfig.fir@123307.4]
);
  wire  _T; // @[ALU.scala 40:29:freechips.rocketchip.system.TinyConfig.fir@123312.4]
  wire [31:0] _T_1; // @[ALU.scala 62:35:freechips.rocketchip.system.TinyConfig.fir@123313.4]
  wire [31:0] in2_inv; // @[ALU.scala 62:20:freechips.rocketchip.system.TinyConfig.fir@123314.4]
  wire [31:0] in1_xor_in2; // @[ALU.scala 63:28:freechips.rocketchip.system.TinyConfig.fir@123315.4]
  wire [31:0] _T_3; // @[ALU.scala 64:26:freechips.rocketchip.system.TinyConfig.fir@123317.4]
  wire [31:0] _GEN_0; // @[ALU.scala 64:36:freechips.rocketchip.system.TinyConfig.fir@123319.4]
  wire  _T_7; // @[ALU.scala 68:15:freechips.rocketchip.system.TinyConfig.fir@123322.4]
  wire  _T_8; // @[ALU.scala 68:34:freechips.rocketchip.system.TinyConfig.fir@123323.4]
  wire  _T_9; // @[ALU.scala 68:24:freechips.rocketchip.system.TinyConfig.fir@123324.4]
  wire  _T_10; // @[ALU.scala 68:56:freechips.rocketchip.system.TinyConfig.fir@123325.4]
  wire  _T_11; // @[ALU.scala 42:35:freechips.rocketchip.system.TinyConfig.fir@123326.4]
  wire  _T_14; // @[ALU.scala 69:8:freechips.rocketchip.system.TinyConfig.fir@123329.4]
  wire  slt; // @[ALU.scala 68:8:freechips.rocketchip.system.TinyConfig.fir@123330.4]
  wire  _T_15; // @[ALU.scala 43:35:freechips.rocketchip.system.TinyConfig.fir@123331.4]
  wire  _T_17; // @[ALU.scala 44:26:freechips.rocketchip.system.TinyConfig.fir@123333.4]
  wire  _T_18; // @[ALU.scala 70:68:freechips.rocketchip.system.TinyConfig.fir@123334.4]
  wire  _T_19; // @[ALU.scala 70:41:freechips.rocketchip.system.TinyConfig.fir@123335.4]
  wire [4:0] shamt; // @[ALU.scala 74:28:freechips.rocketchip.system.TinyConfig.fir@123338.4]
  wire  _T_21; // @[ALU.scala 82:24:freechips.rocketchip.system.TinyConfig.fir@123339.4]
  wire  _T_22; // @[ALU.scala 82:44:freechips.rocketchip.system.TinyConfig.fir@123340.4]
  wire  _T_23; // @[ALU.scala 82:35:freechips.rocketchip.system.TinyConfig.fir@123341.4]
  wire [15:0] _T_26; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123344.4]
  wire [31:0] _T_27; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123345.4]
  wire [15:0] _T_28; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123346.4]
  wire [31:0] _T_29; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123347.4]
  wire [31:0] _T_31; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123349.4]
  wire [31:0] _T_32; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123350.4]
  wire [23:0] _T_36; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123354.4]
  wire [31:0] _GEN_1; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123355.4]
  wire [31:0] _T_37; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123355.4]
  wire [23:0] _T_38; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123356.4]
  wire [31:0] _T_39; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123357.4]
  wire [31:0] _T_41; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123359.4]
  wire [31:0] _T_42; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123360.4]
  wire [27:0] _T_46; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123364.4]
  wire [31:0] _GEN_2; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123365.4]
  wire [31:0] _T_47; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123365.4]
  wire [27:0] _T_48; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123366.4]
  wire [31:0] _T_49; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123367.4]
  wire [31:0] _T_51; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123369.4]
  wire [31:0] _T_52; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123370.4]
  wire [29:0] _T_56; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123374.4]
  wire [31:0] _GEN_3; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123375.4]
  wire [31:0] _T_57; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123375.4]
  wire [29:0] _T_58; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123376.4]
  wire [31:0] _T_59; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123377.4]
  wire [31:0] _T_61; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123379.4]
  wire [31:0] _T_62; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123380.4]
  wire [30:0] _T_66; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123384.4]
  wire [31:0] _GEN_4; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123385.4]
  wire [31:0] _T_67; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123385.4]
  wire [30:0] _T_68; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123386.4]
  wire [31:0] _T_69; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123387.4]
  wire [31:0] _T_71; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123389.4]
  wire [31:0] _T_72; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123390.4]
  wire [31:0] shin; // @[ALU.scala 82:17:freechips.rocketchip.system.TinyConfig.fir@123391.4]
  wire  _T_74; // @[ALU.scala 83:41:freechips.rocketchip.system.TinyConfig.fir@123393.4]
  wire  _T_75; // @[ALU.scala 83:35:freechips.rocketchip.system.TinyConfig.fir@123394.4]
  wire [32:0] _T_76; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@123395.4]
  wire [32:0] _T_77; // @[ALU.scala 83:57:freechips.rocketchip.system.TinyConfig.fir@123396.4]
  wire [32:0] _T_78; // @[ALU.scala 83:64:freechips.rocketchip.system.TinyConfig.fir@123397.4]
  wire [31:0] shout_r; // @[ALU.scala 83:73:freechips.rocketchip.system.TinyConfig.fir@123398.4]
  wire [15:0] _T_81; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123401.4]
  wire [31:0] _T_82; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123402.4]
  wire [15:0] _T_83; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123403.4]
  wire [31:0] _T_84; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123404.4]
  wire [31:0] _T_86; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123406.4]
  wire [31:0] _T_87; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123407.4]
  wire [23:0] _T_91; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123411.4]
  wire [31:0] _GEN_5; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123412.4]
  wire [31:0] _T_92; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123412.4]
  wire [23:0] _T_93; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123413.4]
  wire [31:0] _T_94; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123414.4]
  wire [31:0] _T_96; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123416.4]
  wire [31:0] _T_97; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123417.4]
  wire [27:0] _T_101; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123421.4]
  wire [31:0] _GEN_6; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123422.4]
  wire [31:0] _T_102; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123422.4]
  wire [27:0] _T_103; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123423.4]
  wire [31:0] _T_104; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123424.4]
  wire [31:0] _T_106; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123426.4]
  wire [31:0] _T_107; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123427.4]
  wire [29:0] _T_111; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123431.4]
  wire [31:0] _GEN_7; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123432.4]
  wire [31:0] _T_112; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123432.4]
  wire [29:0] _T_113; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123433.4]
  wire [31:0] _T_114; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123434.4]
  wire [31:0] _T_116; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123436.4]
  wire [31:0] _T_117; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123437.4]
  wire [30:0] _T_121; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123441.4]
  wire [31:0] _GEN_8; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123442.4]
  wire [31:0] _T_122; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123442.4]
  wire [30:0] _T_123; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123443.4]
  wire [31:0] _T_124; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123444.4]
  wire [31:0] _T_126; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123446.4]
  wire [31:0] shout_l; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123447.4]
  wire [31:0] _T_130; // @[ALU.scala 85:18:freechips.rocketchip.system.TinyConfig.fir@123451.4]
  wire  _T_131; // @[ALU.scala 86:25:freechips.rocketchip.system.TinyConfig.fir@123452.4]
  wire [31:0] _T_132; // @[ALU.scala 86:18:freechips.rocketchip.system.TinyConfig.fir@123453.4]
  wire [31:0] shout; // @[ALU.scala 85:74:freechips.rocketchip.system.TinyConfig.fir@123454.4]
  wire  _T_133; // @[ALU.scala 89:25:freechips.rocketchip.system.TinyConfig.fir@123455.4]
  wire  _T_134; // @[ALU.scala 89:45:freechips.rocketchip.system.TinyConfig.fir@123456.4]
  wire  _T_135; // @[ALU.scala 89:36:freechips.rocketchip.system.TinyConfig.fir@123457.4]
  wire [31:0] _T_136; // @[ALU.scala 89:18:freechips.rocketchip.system.TinyConfig.fir@123458.4]
  wire  _T_138; // @[ALU.scala 90:44:freechips.rocketchip.system.TinyConfig.fir@123460.4]
  wire  _T_139; // @[ALU.scala 90:35:freechips.rocketchip.system.TinyConfig.fir@123461.4]
  wire [31:0] _T_140; // @[ALU.scala 90:63:freechips.rocketchip.system.TinyConfig.fir@123462.4]
  wire [31:0] _T_141; // @[ALU.scala 90:18:freechips.rocketchip.system.TinyConfig.fir@123463.4]
  wire [31:0] logic_; // @[ALU.scala 89:78:freechips.rocketchip.system.TinyConfig.fir@123464.4]
  wire  _T_142; // @[ALU.scala 41:30:freechips.rocketchip.system.TinyConfig.fir@123465.4]
  wire  _T_143; // @[ALU.scala 91:35:freechips.rocketchip.system.TinyConfig.fir@123466.4]
  wire [31:0] _GEN_9; // @[ALU.scala 91:43:freechips.rocketchip.system.TinyConfig.fir@123467.4]
  wire [31:0] _T_144; // @[ALU.scala 91:43:freechips.rocketchip.system.TinyConfig.fir@123467.4]
  wire [31:0] shift_logic; // @[ALU.scala 91:51:freechips.rocketchip.system.TinyConfig.fir@123468.4]
  wire  _T_145; // @[ALU.scala 92:23:freechips.rocketchip.system.TinyConfig.fir@123469.4]
  wire  _T_146; // @[ALU.scala 92:43:freechips.rocketchip.system.TinyConfig.fir@123470.4]
  wire  _T_147; // @[ALU.scala 92:34:freechips.rocketchip.system.TinyConfig.fir@123471.4]
  assign _T = io_fn[3]; // @[ALU.scala 40:29:freechips.rocketchip.system.TinyConfig.fir@123312.4]
  assign _T_1 = ~ io_in2; // @[ALU.scala 62:35:freechips.rocketchip.system.TinyConfig.fir@123313.4]
  assign in2_inv = _T ? _T_1 : io_in2; // @[ALU.scala 62:20:freechips.rocketchip.system.TinyConfig.fir@123314.4]
  assign in1_xor_in2 = io_in1 ^ in2_inv; // @[ALU.scala 63:28:freechips.rocketchip.system.TinyConfig.fir@123315.4]
  assign _T_3 = io_in1 + in2_inv; // @[ALU.scala 64:26:freechips.rocketchip.system.TinyConfig.fir@123317.4]
  assign _GEN_0 = {{31'd0}, _T}; // @[ALU.scala 64:36:freechips.rocketchip.system.TinyConfig.fir@123319.4]
  assign _T_7 = io_in1[31]; // @[ALU.scala 68:15:freechips.rocketchip.system.TinyConfig.fir@123322.4]
  assign _T_8 = io_in2[31]; // @[ALU.scala 68:34:freechips.rocketchip.system.TinyConfig.fir@123323.4]
  assign _T_9 = _T_7 == _T_8; // @[ALU.scala 68:24:freechips.rocketchip.system.TinyConfig.fir@123324.4]
  assign _T_10 = io_adder_out[31]; // @[ALU.scala 68:56:freechips.rocketchip.system.TinyConfig.fir@123325.4]
  assign _T_11 = io_fn[1]; // @[ALU.scala 42:35:freechips.rocketchip.system.TinyConfig.fir@123326.4]
  assign _T_14 = _T_11 ? _T_8 : _T_7; // @[ALU.scala 69:8:freechips.rocketchip.system.TinyConfig.fir@123329.4]
  assign slt = _T_9 ? _T_10 : _T_14; // @[ALU.scala 68:8:freechips.rocketchip.system.TinyConfig.fir@123330.4]
  assign _T_15 = io_fn[0]; // @[ALU.scala 43:35:freechips.rocketchip.system.TinyConfig.fir@123331.4]
  assign _T_17 = _T == 1'h0; // @[ALU.scala 44:26:freechips.rocketchip.system.TinyConfig.fir@123333.4]
  assign _T_18 = in1_xor_in2 == 32'h0; // @[ALU.scala 70:68:freechips.rocketchip.system.TinyConfig.fir@123334.4]
  assign _T_19 = _T_17 ? _T_18 : slt; // @[ALU.scala 70:41:freechips.rocketchip.system.TinyConfig.fir@123335.4]
  assign shamt = io_in2[4:0]; // @[ALU.scala 74:28:freechips.rocketchip.system.TinyConfig.fir@123338.4]
  assign _T_21 = io_fn == 4'h5; // @[ALU.scala 82:24:freechips.rocketchip.system.TinyConfig.fir@123339.4]
  assign _T_22 = io_fn == 4'hb; // @[ALU.scala 82:44:freechips.rocketchip.system.TinyConfig.fir@123340.4]
  assign _T_23 = _T_21 | _T_22; // @[ALU.scala 82:35:freechips.rocketchip.system.TinyConfig.fir@123341.4]
  assign _T_26 = io_in1[31:16]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123344.4]
  assign _T_27 = {{16'd0}, _T_26}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123345.4]
  assign _T_28 = io_in1[15:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123346.4]
  assign _T_29 = {_T_28, 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123347.4]
  assign _T_31 = _T_29 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123349.4]
  assign _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123350.4]
  assign _T_36 = _T_32[31:8]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123354.4]
  assign _GEN_1 = {{8'd0}, _T_36}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123355.4]
  assign _T_37 = _GEN_1 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123355.4]
  assign _T_38 = _T_32[23:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123356.4]
  assign _T_39 = {_T_38, 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123357.4]
  assign _T_41 = _T_39 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123359.4]
  assign _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123360.4]
  assign _T_46 = _T_42[31:4]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123364.4]
  assign _GEN_2 = {{4'd0}, _T_46}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123365.4]
  assign _T_47 = _GEN_2 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123365.4]
  assign _T_48 = _T_42[27:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123366.4]
  assign _T_49 = {_T_48, 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123367.4]
  assign _T_51 = _T_49 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123369.4]
  assign _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123370.4]
  assign _T_56 = _T_52[31:2]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123374.4]
  assign _GEN_3 = {{2'd0}, _T_56}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123375.4]
  assign _T_57 = _GEN_3 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123375.4]
  assign _T_58 = _T_52[29:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123376.4]
  assign _T_59 = {_T_58, 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123377.4]
  assign _T_61 = _T_59 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123379.4]
  assign _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123380.4]
  assign _T_66 = _T_62[31:1]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123384.4]
  assign _GEN_4 = {{1'd0}, _T_66}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123385.4]
  assign _T_67 = _GEN_4 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123385.4]
  assign _T_68 = _T_62[30:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123386.4]
  assign _T_69 = {_T_68, 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123387.4]
  assign _T_71 = _T_69 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123389.4]
  assign _T_72 = _T_67 | _T_71; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123390.4]
  assign shin = _T_23 ? io_in1 : _T_72; // @[ALU.scala 82:17:freechips.rocketchip.system.TinyConfig.fir@123391.4]
  assign _T_74 = shin[31]; // @[ALU.scala 83:41:freechips.rocketchip.system.TinyConfig.fir@123393.4]
  assign _T_75 = _T & _T_74; // @[ALU.scala 83:35:freechips.rocketchip.system.TinyConfig.fir@123394.4]
  assign _T_76 = {_T_75,shin}; // @[Cat.scala 30:58:freechips.rocketchip.system.TinyConfig.fir@123395.4]
  assign _T_77 = $signed(_T_76); // @[ALU.scala 83:57:freechips.rocketchip.system.TinyConfig.fir@123396.4]
  assign _T_78 = $signed(_T_77) >>> shamt; // @[ALU.scala 83:64:freechips.rocketchip.system.TinyConfig.fir@123397.4]
  assign shout_r = _T_78[31:0]; // @[ALU.scala 83:73:freechips.rocketchip.system.TinyConfig.fir@123398.4]
  assign _T_81 = shout_r[31:16]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123401.4]
  assign _T_82 = {{16'd0}, _T_81}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123402.4]
  assign _T_83 = shout_r[15:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123403.4]
  assign _T_84 = {_T_83, 16'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123404.4]
  assign _T_86 = _T_84 & 32'hffff0000; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123406.4]
  assign _T_87 = _T_82 | _T_86; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123407.4]
  assign _T_91 = _T_87[31:8]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123411.4]
  assign _GEN_5 = {{8'd0}, _T_91}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123412.4]
  assign _T_92 = _GEN_5 & 32'hff00ff; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123412.4]
  assign _T_93 = _T_87[23:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123413.4]
  assign _T_94 = {_T_93, 8'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123414.4]
  assign _T_96 = _T_94 & 32'hff00ff00; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123416.4]
  assign _T_97 = _T_92 | _T_96; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123417.4]
  assign _T_101 = _T_97[31:4]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123421.4]
  assign _GEN_6 = {{4'd0}, _T_101}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123422.4]
  assign _T_102 = _GEN_6 & 32'hf0f0f0f; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123422.4]
  assign _T_103 = _T_97[27:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123423.4]
  assign _T_104 = {_T_103, 4'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123424.4]
  assign _T_106 = _T_104 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123426.4]
  assign _T_107 = _T_102 | _T_106; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123427.4]
  assign _T_111 = _T_107[31:2]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123431.4]
  assign _GEN_7 = {{2'd0}, _T_111}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123432.4]
  assign _T_112 = _GEN_7 & 32'h33333333; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123432.4]
  assign _T_113 = _T_107[29:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123433.4]
  assign _T_114 = {_T_113, 2'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123434.4]
  assign _T_116 = _T_114 & 32'hcccccccc; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123436.4]
  assign _T_117 = _T_112 | _T_116; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123437.4]
  assign _T_121 = _T_117[31:1]; // @[Bitwise.scala 103:21:freechips.rocketchip.system.TinyConfig.fir@123441.4]
  assign _GEN_8 = {{1'd0}, _T_121}; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123442.4]
  assign _T_122 = _GEN_8 & 32'h55555555; // @[Bitwise.scala 103:31:freechips.rocketchip.system.TinyConfig.fir@123442.4]
  assign _T_123 = _T_117[30:0]; // @[Bitwise.scala 103:46:freechips.rocketchip.system.TinyConfig.fir@123443.4]
  assign _T_124 = {_T_123, 1'h0}; // @[Bitwise.scala 103:65:freechips.rocketchip.system.TinyConfig.fir@123444.4]
  assign _T_126 = _T_124 & 32'haaaaaaaa; // @[Bitwise.scala 103:75:freechips.rocketchip.system.TinyConfig.fir@123446.4]
  assign shout_l = _T_122 | _T_126; // @[Bitwise.scala 103:39:freechips.rocketchip.system.TinyConfig.fir@123447.4]
  assign _T_130 = _T_23 ? shout_r : 32'h0; // @[ALU.scala 85:18:freechips.rocketchip.system.TinyConfig.fir@123451.4]
  assign _T_131 = io_fn == 4'h1; // @[ALU.scala 86:25:freechips.rocketchip.system.TinyConfig.fir@123452.4]
  assign _T_132 = _T_131 ? shout_l : 32'h0; // @[ALU.scala 86:18:freechips.rocketchip.system.TinyConfig.fir@123453.4]
  assign shout = _T_130 | _T_132; // @[ALU.scala 85:74:freechips.rocketchip.system.TinyConfig.fir@123454.4]
  assign _T_133 = io_fn == 4'h4; // @[ALU.scala 89:25:freechips.rocketchip.system.TinyConfig.fir@123455.4]
  assign _T_134 = io_fn == 4'h6; // @[ALU.scala 89:45:freechips.rocketchip.system.TinyConfig.fir@123456.4]
  assign _T_135 = _T_133 | _T_134; // @[ALU.scala 89:36:freechips.rocketchip.system.TinyConfig.fir@123457.4]
  assign _T_136 = _T_135 ? in1_xor_in2 : 32'h0; // @[ALU.scala 89:18:freechips.rocketchip.system.TinyConfig.fir@123458.4]
  assign _T_138 = io_fn == 4'h7; // @[ALU.scala 90:44:freechips.rocketchip.system.TinyConfig.fir@123460.4]
  assign _T_139 = _T_134 | _T_138; // @[ALU.scala 90:35:freechips.rocketchip.system.TinyConfig.fir@123461.4]
  assign _T_140 = io_in1 & io_in2; // @[ALU.scala 90:63:freechips.rocketchip.system.TinyConfig.fir@123462.4]
  assign _T_141 = _T_139 ? _T_140 : 32'h0; // @[ALU.scala 90:18:freechips.rocketchip.system.TinyConfig.fir@123463.4]
  assign logic_ = _T_136 | _T_141; // @[ALU.scala 89:78:freechips.rocketchip.system.TinyConfig.fir@123464.4]
  assign _T_142 = io_fn >= 4'hc; // @[ALU.scala 41:30:freechips.rocketchip.system.TinyConfig.fir@123465.4]
  assign _T_143 = _T_142 & slt; // @[ALU.scala 91:35:freechips.rocketchip.system.TinyConfig.fir@123466.4]
  assign _GEN_9 = {{31'd0}, _T_143}; // @[ALU.scala 91:43:freechips.rocketchip.system.TinyConfig.fir@123467.4]
  assign _T_144 = _GEN_9 | logic_; // @[ALU.scala 91:43:freechips.rocketchip.system.TinyConfig.fir@123467.4]
  assign shift_logic = _T_144 | shout; // @[ALU.scala 91:51:freechips.rocketchip.system.TinyConfig.fir@123468.4]
  assign _T_145 = io_fn == 4'h0; // @[ALU.scala 92:23:freechips.rocketchip.system.TinyConfig.fir@123469.4]
  assign _T_146 = io_fn == 4'ha; // @[ALU.scala 92:43:freechips.rocketchip.system.TinyConfig.fir@123470.4]
  assign _T_147 = _T_145 | _T_146; // @[ALU.scala 92:34:freechips.rocketchip.system.TinyConfig.fir@123471.4]
  assign io_out = _T_147 ? io_adder_out : shift_logic; // @[ALU.scala 94:10:freechips.rocketchip.system.TinyConfig.fir@123473.4]
  assign io_adder_out = _T_3 + _GEN_0; // @[ALU.scala 64:16:freechips.rocketchip.system.TinyConfig.fir@123321.4]
  assign io_cmp_out = _T_15 ^ _T_19; // @[ALU.scala 70:14:freechips.rocketchip.system.TinyConfig.fir@123337.4]
endmodule