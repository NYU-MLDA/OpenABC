module MulAddRecFN_postMul_0
(
  io_fromPreMul_highExpA,
  io_fromPreMul_isNaN_isQuietNaNA,
  io_fromPreMul_highExpB,
  io_fromPreMul_isNaN_isQuietNaNB,
  io_fromPreMul_signProd,
  io_fromPreMul_isZeroProd,
  io_fromPreMul_opSignC,
  io_fromPreMul_highExpC,
  io_fromPreMul_isNaN_isQuietNaNC,
  io_fromPreMul_isCDominant,
  io_fromPreMul_CAlignDist_0,
  io_fromPreMul_CAlignDist,
  io_fromPreMul_bit0AlignedNegSigC,
  io_fromPreMul_highAlignedNegSigC,
  io_fromPreMul_sExpSum,
  io_fromPreMul_roundingMode,
  io_mulAddResult,
  io_out,
  io_exceptionFlags
);

  input [2:0] io_fromPreMul_highExpA;
  input [2:0] io_fromPreMul_highExpB;
  input [2:0] io_fromPreMul_highExpC;
  input [6:0] io_fromPreMul_CAlignDist;
  input [25:0] io_fromPreMul_highAlignedNegSigC;
  input [10:0] io_fromPreMul_sExpSum;
  input [1:0] io_fromPreMul_roundingMode;
  input [48:0] io_mulAddResult;
  output [32:0] io_out;
  output [4:0] io_exceptionFlags;
  input io_fromPreMul_isNaN_isQuietNaNA;
  input io_fromPreMul_isNaN_isQuietNaNB;
  input io_fromPreMul_signProd;
  input io_fromPreMul_isZeroProd;
  input io_fromPreMul_opSignC;
  input io_fromPreMul_isNaN_isQuietNaNC;
  input io_fromPreMul_isCDominant;
  input io_fromPreMul_CAlignDist_0;
  input io_fromPreMul_bit0AlignedNegSigC;
  wire [32:0] io_out;
  wire [4:0] io_exceptionFlags,T395,T396,T397,T398,T399,T400,T401,T402,T403,T404,T405,T406,
  T407,T408,T409,T410,T475;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,T3,
  commonCase,inexactY,doIncrSig,N132,T215,anyRound,sigX3_27,T77_0,N133,N134,N135,N136,
  N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,
  N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
  N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,T32,N182,T34_5,
  T34_3,T34_1,T35_4,T35_2,T38_3,T38_2,T53_13,T53_11,T53_9,T53_7,T53_5,T53_3,T53_1,
  T54_12,T54_10,T54_8,T54_6,T54_4,T54_2,T57_11,T57_10,T57_7,T57_6,T57_3,T57_2,T58_9,
  T58_8,T58_5,T58_4,T61_7,T61_6,T61_5,T61_4,absSigSumExtraMask_1,T107_5,T107_3,
  T107_1,T108_4,T108_2,T111_3,T111_2,N183,N184,N185,T128_0,N186,T138,T148_0,T159,T168,
  T170,T178,T181,T187,T191,T189,allRound,T219,T221,T220,T223,T222,
  notSpecial_addZeros,addSpecial,mulSpecial,underflowY,T227,T228,sigX3Shift1,N187,roundEven,N188,
  T247,T244,T246,T245,T248,T249,T252,N189,T259,T253,roundDirectUp,signY,N190,
  isZeroY,N191,T255,doNegSignSum,N192,T256,T257,T262,T260,T261,T264,T263,T268,T265,T266,
  T267,T269,T270,T271,T276,N193,T279,T278,N194,N195,T305,notSigNaN_invalid,T302,
  T287,T288,T291,isInfC,T289,T297,T292,isInfA,isInfB,T293,T295,T300,T298,isNaNB,
  isNaNA,T304,T303,T308,isSigNaNC,isNaNC,T306,isSigNaNA,isSigNaNB,T309,T310,T313_0,
  T314,overflowY_roundMagUp,roundMagUp,T317,T315,T316,T320,T321,T325,N196,T326,
  totalUnderflowY,T331,T327,T328,notNaN_isInfOut,T336,T335,T337,pegMinFiniteMagOut,T342,
  notSpecial_isZeroOut,T355,T357,T356,T372,uncommonCaseSignOut,T362,T358,T359,
  T360,T361,T366,T363,T364,T365,T370,T367,T368,T369,T371,N197,N198,N199,N200,N201,
  N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,
  N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,
  N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,
  N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,
  N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,
  N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,
  N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,
  N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,
  N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,
  N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,
  N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,
  N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,
  N394,N395,N396,N397,N398,N399,N400,SV2V_UNCONNECTED_1,SV2V_UNCONNECTED_2,
  SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,
  SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,SV2V_UNCONNECTED_9,
  SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11,SV2V_UNCONNECTED_12,
  SV2V_UNCONNECTED_13,SV2V_UNCONNECTED_14,SV2V_UNCONNECTED_15,
  SV2V_UNCONNECTED_16,SV2V_UNCONNECTED_17,SV2V_UNCONNECTED_18,SV2V_UNCONNECTED_19,
  SV2V_UNCONNECTED_20,SV2V_UNCONNECTED_21,SV2V_UNCONNECTED_22,
  SV2V_UNCONNECTED_23,SV2V_UNCONNECTED_24,SV2V_UNCONNECTED_25,
  SV2V_UNCONNECTED_26,SV2V_UNCONNECTED_27,SV2V_UNCONNECTED_28,SV2V_UNCONNECTED_29,
  SV2V_UNCONNECTED_30,SV2V_UNCONNECTED_31,SV2V_UNCONNECTED_32,
  SV2V_UNCONNECTED_33,SV2V_UNCONNECTED_34,SV2V_UNCONNECTED_35,
  SV2V_UNCONNECTED_36,SV2V_UNCONNECTED_37,SV2V_UNCONNECTED_38,SV2V_UNCONNECTED_39,
  SV2V_UNCONNECTED_40,SV2V_UNCONNECTED_41,SV2V_UNCONNECTED_42,
  SV2V_UNCONNECTED_43,SV2V_UNCONNECTED_44,SV2V_UNCONNECTED_45,
  SV2V_UNCONNECTED_46,SV2V_UNCONNECTED_47,SV2V_UNCONNECTED_48,SV2V_UNCONNECTED_49,
  SV2V_UNCONNECTED_50,SV2V_UNCONNECTED_51,SV2V_UNCONNECTED_52,
  SV2V_UNCONNECTED_53,SV2V_UNCONNECTED_54,SV2V_UNCONNECTED_55,
  SV2V_UNCONNECTED_56,SV2V_UNCONNECTED_57,SV2V_UNCONNECTED_58,SV2V_UNCONNECTED_59,
  SV2V_UNCONNECTED_60,SV2V_UNCONNECTED_61,SV2V_UNCONNECTED_62,
  SV2V_UNCONNECTED_63,SV2V_UNCONNECTED_64,SV2V_UNCONNECTED_65,
  SV2V_UNCONNECTED_66,SV2V_UNCONNECTED_67,SV2V_UNCONNECTED_68,SV2V_UNCONNECTED_69,
  SV2V_UNCONNECTED_70,SV2V_UNCONNECTED_71,SV2V_UNCONNECTED_72,
  SV2V_UNCONNECTED_73,SV2V_UNCONNECTED_74,SV2V_UNCONNECTED_75,
  SV2V_UNCONNECTED_76,SV2V_UNCONNECTED_77,SV2V_UNCONNECTED_78,SV2V_UNCONNECTED_79,
  SV2V_UNCONNECTED_80,SV2V_UNCONNECTED_81,SV2V_UNCONNECTED_82,
  SV2V_UNCONNECTED_83,SV2V_UNCONNECTED_84,SV2V_UNCONNECTED_85,
  SV2V_UNCONNECTED_86,SV2V_UNCONNECTED_87,SV2V_UNCONNECTED_88,SV2V_UNCONNECTED_89,
  SV2V_UNCONNECTED_90,SV2V_UNCONNECTED_91,SV2V_UNCONNECTED_92,
  SV2V_UNCONNECTED_93,SV2V_UNCONNECTED_94,SV2V_UNCONNECTED_95,
  SV2V_UNCONNECTED_96,SV2V_UNCONNECTED_97,SV2V_UNCONNECTED_98,SV2V_UNCONNECTED_99,
  SV2V_UNCONNECTED_100,SV2V_UNCONNECTED_101,SV2V_UNCONNECTED_102,
  SV2V_UNCONNECTED_103,SV2V_UNCONNECTED_104,SV2V_UNCONNECTED_105,
  SV2V_UNCONNECTED_106,SV2V_UNCONNECTED_107,SV2V_UNCONNECTED_108,
  SV2V_UNCONNECTED_109,SV2V_UNCONNECTED_110,SV2V_UNCONNECTED_111,
  SV2V_UNCONNECTED_112,SV2V_UNCONNECTED_113,SV2V_UNCONNECTED_114,SV2V_UNCONNECTED_115,
  SV2V_UNCONNECTED_116,SV2V_UNCONNECTED_117,SV2V_UNCONNECTED_118,
  SV2V_UNCONNECTED_119,SV2V_UNCONNECTED_120,SV2V_UNCONNECTED_121,
  SV2V_UNCONNECTED_122,SV2V_UNCONNECTED_123,SV2V_UNCONNECTED_124,
  SV2V_UNCONNECTED_125,SV2V_UNCONNECTED_126,SV2V_UNCONNECTED_127,
  SV2V_UNCONNECTED_128,SV2V_UNCONNECTED_129,SV2V_UNCONNECTED_130,SV2V_UNCONNECTED_131,
  SV2V_UNCONNECTED_132,SV2V_UNCONNECTED_133,SV2V_UNCONNECTED_134,
  SV2V_UNCONNECTED_135,SV2V_UNCONNECTED_136,SV2V_UNCONNECTED_137,
  SV2V_UNCONNECTED_138,SV2V_UNCONNECTED_139,SV2V_UNCONNECTED_140,
  SV2V_UNCONNECTED_141,SV2V_UNCONNECTED_142,SV2V_UNCONNECTED_143,
  SV2V_UNCONNECTED_144,SV2V_UNCONNECTED_145,SV2V_UNCONNECTED_146,SV2V_UNCONNECTED_147,
  SV2V_UNCONNECTED_148,SV2V_UNCONNECTED_149,SV2V_UNCONNECTED_150,
  SV2V_UNCONNECTED_151,SV2V_UNCONNECTED_152,SV2V_UNCONNECTED_153,
  SV2V_UNCONNECTED_154,SV2V_UNCONNECTED_155,SV2V_UNCONNECTED_156,
  SV2V_UNCONNECTED_157,SV2V_UNCONNECTED_158,SV2V_UNCONNECTED_159,
  SV2V_UNCONNECTED_160,SV2V_UNCONNECTED_161,SV2V_UNCONNECTED_162,SV2V_UNCONNECTED_163,
  SV2V_UNCONNECTED_164,SV2V_UNCONNECTED_165,SV2V_UNCONNECTED_166,
  SV2V_UNCONNECTED_167,SV2V_UNCONNECTED_168,SV2V_UNCONNECTED_169,
  SV2V_UNCONNECTED_170,SV2V_UNCONNECTED_171,SV2V_UNCONNECTED_172,
  SV2V_UNCONNECTED_173,SV2V_UNCONNECTED_174,SV2V_UNCONNECTED_175,
  SV2V_UNCONNECTED_176,SV2V_UNCONNECTED_177,SV2V_UNCONNECTED_178,SV2V_UNCONNECTED_179,
  SV2V_UNCONNECTED_180,SV2V_UNCONNECTED_181,SV2V_UNCONNECTED_182,
  SV2V_UNCONNECTED_183,SV2V_UNCONNECTED_184,SV2V_UNCONNECTED_185,
  SV2V_UNCONNECTED_186,SV2V_UNCONNECTED_187,SV2V_UNCONNECTED_188,
  SV2V_UNCONNECTED_189,SV2V_UNCONNECTED_190,SV2V_UNCONNECTED_191,
  SV2V_UNCONNECTED_192,SV2V_UNCONNECTED_193,SV2V_UNCONNECTED_194,SV2V_UNCONNECTED_195,
  SV2V_UNCONNECTED_196,SV2V_UNCONNECTED_197,SV2V_UNCONNECTED_198,
  SV2V_UNCONNECTED_199,SV2V_UNCONNECTED_200,SV2V_UNCONNECTED_201,
  SV2V_UNCONNECTED_202,SV2V_UNCONNECTED_203,SV2V_UNCONNECTED_204,
  SV2V_UNCONNECTED_205,SV2V_UNCONNECTED_206,SV2V_UNCONNECTED_207,
  SV2V_UNCONNECTED_208,SV2V_UNCONNECTED_209,SV2V_UNCONNECTED_210,SV2V_UNCONNECTED_211,
  SV2V_UNCONNECTED_212,SV2V_UNCONNECTED_213,SV2V_UNCONNECTED_214,
  SV2V_UNCONNECTED_215,SV2V_UNCONNECTED_216,SV2V_UNCONNECTED_217,
  SV2V_UNCONNECTED_218,SV2V_UNCONNECTED_219,SV2V_UNCONNECTED_220,
  SV2V_UNCONNECTED_221,SV2V_UNCONNECTED_222,SV2V_UNCONNECTED_223,
  SV2V_UNCONNECTED_224,SV2V_UNCONNECTED_225,SV2V_UNCONNECTED_226,SV2V_UNCONNECTED_227,
  SV2V_UNCONNECTED_228,SV2V_UNCONNECTED_229,SV2V_UNCONNECTED_230,
  SV2V_UNCONNECTED_231,SV2V_UNCONNECTED_232,SV2V_UNCONNECTED_233,
  SV2V_UNCONNECTED_234,SV2V_UNCONNECTED_235,SV2V_UNCONNECTED_236,
  SV2V_UNCONNECTED_237,SV2V_UNCONNECTED_238,SV2V_UNCONNECTED_239,
  SV2V_UNCONNECTED_240,SV2V_UNCONNECTED_241,SV2V_UNCONNECTED_242,SV2V_UNCONNECTED_243,
  SV2V_UNCONNECTED_244,SV2V_UNCONNECTED_245,SV2V_UNCONNECTED_246,
  SV2V_UNCONNECTED_247,SV2V_UNCONNECTED_248,SV2V_UNCONNECTED_249,
  SV2V_UNCONNECTED_250,SV2V_UNCONNECTED_251,SV2V_UNCONNECTED_252,
  SV2V_UNCONNECTED_253,SV2V_UNCONNECTED_254,SV2V_UNCONNECTED_255,
  SV2V_UNCONNECTED_256,SV2V_UNCONNECTED_257,SV2V_UNCONNECTED_258,SV2V_UNCONNECTED_259,
  SV2V_UNCONNECTED_260,SV2V_UNCONNECTED_261,SV2V_UNCONNECTED_262,
  SV2V_UNCONNECTED_263,SV2V_UNCONNECTED_264,SV2V_UNCONNECTED_265,
  SV2V_UNCONNECTED_266,SV2V_UNCONNECTED_267,SV2V_UNCONNECTED_268,
  SV2V_UNCONNECTED_269,SV2V_UNCONNECTED_270,SV2V_UNCONNECTED_271,
  SV2V_UNCONNECTED_272,SV2V_UNCONNECTED_273,SV2V_UNCONNECTED_274,SV2V_UNCONNECTED_275,
  SV2V_UNCONNECTED_276,SV2V_UNCONNECTED_277,SV2V_UNCONNECTED_278,
  SV2V_UNCONNECTED_279,SV2V_UNCONNECTED_280,SV2V_UNCONNECTED_281,
  SV2V_UNCONNECTED_282,SV2V_UNCONNECTED_283,SV2V_UNCONNECTED_284,
  SV2V_UNCONNECTED_285,SV2V_UNCONNECTED_286,SV2V_UNCONNECTED_287,
  SV2V_UNCONNECTED_288,SV2V_UNCONNECTED_289,SV2V_UNCONNECTED_290,SV2V_UNCONNECTED_291,
  SV2V_UNCONNECTED_292,SV2V_UNCONNECTED_293,SV2V_UNCONNECTED_294,
  SV2V_UNCONNECTED_295,SV2V_UNCONNECTED_296,SV2V_UNCONNECTED_297,
  SV2V_UNCONNECTED_298,SV2V_UNCONNECTED_299,SV2V_UNCONNECTED_300,
  SV2V_UNCONNECTED_301,SV2V_UNCONNECTED_302,SV2V_UNCONNECTED_303,
  SV2V_UNCONNECTED_304,SV2V_UNCONNECTED_305,SV2V_UNCONNECTED_306,SV2V_UNCONNECTED_307,
  SV2V_UNCONNECTED_308,SV2V_UNCONNECTED_309,SV2V_UNCONNECTED_310,
  SV2V_UNCONNECTED_311,SV2V_UNCONNECTED_312,SV2V_UNCONNECTED_313,
  SV2V_UNCONNECTED_314,SV2V_UNCONNECTED_315,SV2V_UNCONNECTED_316,
  SV2V_UNCONNECTED_317,SV2V_UNCONNECTED_318,SV2V_UNCONNECTED_319,
  SV2V_UNCONNECTED_320,SV2V_UNCONNECTED_321,SV2V_UNCONNECTED_322,SV2V_UNCONNECTED_323,
  SV2V_UNCONNECTED_324,SV2V_UNCONNECTED_325,SV2V_UNCONNECTED_326,
  SV2V_UNCONNECTED_327,SV2V_UNCONNECTED_328,SV2V_UNCONNECTED_329,
  SV2V_UNCONNECTED_330,SV2V_UNCONNECTED_331,SV2V_UNCONNECTED_332,
  SV2V_UNCONNECTED_333,SV2V_UNCONNECTED_334,SV2V_UNCONNECTED_335,
  SV2V_UNCONNECTED_336,SV2V_UNCONNECTED_337,SV2V_UNCONNECTED_338,SV2V_UNCONNECTED_339,
  SV2V_UNCONNECTED_340,SV2V_UNCONNECTED_341,SV2V_UNCONNECTED_342,
  SV2V_UNCONNECTED_343,SV2V_UNCONNECTED_344,SV2V_UNCONNECTED_345,
  SV2V_UNCONNECTED_346,SV2V_UNCONNECTED_347,SV2V_UNCONNECTED_348,
  SV2V_UNCONNECTED_349,SV2V_UNCONNECTED_350,SV2V_UNCONNECTED_351,
  SV2V_UNCONNECTED_352,SV2V_UNCONNECTED_353,SV2V_UNCONNECTED_354,SV2V_UNCONNECTED_355,
  SV2V_UNCONNECTED_356,SV2V_UNCONNECTED_357,SV2V_UNCONNECTED_358,
  SV2V_UNCONNECTED_359,SV2V_UNCONNECTED_360,SV2V_UNCONNECTED_361,
  SV2V_UNCONNECTED_362,SV2V_UNCONNECTED_363,SV2V_UNCONNECTED_364,
  SV2V_UNCONNECTED_365,SV2V_UNCONNECTED_366,SV2V_UNCONNECTED_367,
  SV2V_UNCONNECTED_368,SV2V_UNCONNECTED_369,SV2V_UNCONNECTED_370,SV2V_UNCONNECTED_371,
  SV2V_UNCONNECTED_372,SV2V_UNCONNECTED_373,SV2V_UNCONNECTED_374,
  SV2V_UNCONNECTED_375,SV2V_UNCONNECTED_376,SV2V_UNCONNECTED_377,
  SV2V_UNCONNECTED_378,SV2V_UNCONNECTED_379,SV2V_UNCONNECTED_380,
  SV2V_UNCONNECTED_381,SV2V_UNCONNECTED_382,SV2V_UNCONNECTED_383,
  SV2V_UNCONNECTED_384,SV2V_UNCONNECTED_385,SV2V_UNCONNECTED_386,SV2V_UNCONNECTED_387,
  SV2V_UNCONNECTED_388,SV2V_UNCONNECTED_389,SV2V_UNCONNECTED_390,
  SV2V_UNCONNECTED_391,SV2V_UNCONNECTED_392,SV2V_UNCONNECTED_393,
  SV2V_UNCONNECTED_394,SV2V_UNCONNECTED_395,SV2V_UNCONNECTED_396,
  SV2V_UNCONNECTED_397,SV2V_UNCONNECTED_398,SV2V_UNCONNECTED_399,
  SV2V_UNCONNECTED_400,SV2V_UNCONNECTED_401,SV2V_UNCONNECTED_402,SV2V_UNCONNECTED_403,
  SV2V_UNCONNECTED_404,SV2V_UNCONNECTED_405,SV2V_UNCONNECTED_406,
  SV2V_UNCONNECTED_407,SV2V_UNCONNECTED_408,SV2V_UNCONNECTED_409,
  SV2V_UNCONNECTED_410,SV2V_UNCONNECTED_411,SV2V_UNCONNECTED_412,
  SV2V_UNCONNECTED_413,SV2V_UNCONNECTED_414,SV2V_UNCONNECTED_415,
  SV2V_UNCONNECTED_416,SV2V_UNCONNECTED_417,SV2V_UNCONNECTED_418,SV2V_UNCONNECTED_419,
  SV2V_UNCONNECTED_420,SV2V_UNCONNECTED_421,SV2V_UNCONNECTED_422,
  SV2V_UNCONNECTED_423,SV2V_UNCONNECTED_424,SV2V_UNCONNECTED_425,
  SV2V_UNCONNECTED_426,SV2V_UNCONNECTED_427,SV2V_UNCONNECTED_428,
  SV2V_UNCONNECTED_429,SV2V_UNCONNECTED_430,SV2V_UNCONNECTED_431,
  SV2V_UNCONNECTED_432,SV2V_UNCONNECTED_433,SV2V_UNCONNECTED_434,SV2V_UNCONNECTED_435,
  SV2V_UNCONNECTED_436,SV2V_UNCONNECTED_437,SV2V_UNCONNECTED_438,
  SV2V_UNCONNECTED_439,SV2V_UNCONNECTED_440,SV2V_UNCONNECTED_441,
  SV2V_UNCONNECTED_442,SV2V_UNCONNECTED_443,SV2V_UNCONNECTED_444,
  SV2V_UNCONNECTED_445,SV2V_UNCONNECTED_446,SV2V_UNCONNECTED_447,
  SV2V_UNCONNECTED_448,SV2V_UNCONNECTED_449,SV2V_UNCONNECTED_450,SV2V_UNCONNECTED_451,
  SV2V_UNCONNECTED_452,SV2V_UNCONNECTED_453,SV2V_UNCONNECTED_454,
  SV2V_UNCONNECTED_455,SV2V_UNCONNECTED_456,SV2V_UNCONNECTED_457,
  SV2V_UNCONNECTED_458,SV2V_UNCONNECTED_459,SV2V_UNCONNECTED_460,
  SV2V_UNCONNECTED_461,SV2V_UNCONNECTED_462,SV2V_UNCONNECTED_463,
  SV2V_UNCONNECTED_464,SV2V_UNCONNECTED_465,SV2V_UNCONNECTED_466,SV2V_UNCONNECTED_467,
  SV2V_UNCONNECTED_468,SV2V_UNCONNECTED_469,SV2V_UNCONNECTED_470,
  SV2V_UNCONNECTED_471,SV2V_UNCONNECTED_472,SV2V_UNCONNECTED_473,
  SV2V_UNCONNECTED_474,SV2V_UNCONNECTED_475,SV2V_UNCONNECTED_476,
  SV2V_UNCONNECTED_477,SV2V_UNCONNECTED_478,SV2V_UNCONNECTED_479,
  SV2V_UNCONNECTED_480,SV2V_UNCONNECTED_481,SV2V_UNCONNECTED_482,SV2V_UNCONNECTED_483,
  SV2V_UNCONNECTED_484,SV2V_UNCONNECTED_485,SV2V_UNCONNECTED_486,
  SV2V_UNCONNECTED_487,SV2V_UNCONNECTED_488,SV2V_UNCONNECTED_489,
  SV2V_UNCONNECTED_490,SV2V_UNCONNECTED_491,SV2V_UNCONNECTED_492,
  SV2V_UNCONNECTED_493,SV2V_UNCONNECTED_494,SV2V_UNCONNECTED_495,
  SV2V_UNCONNECTED_496,SV2V_UNCONNECTED_497,SV2V_UNCONNECTED_498,SV2V_UNCONNECTED_499,
  SV2V_UNCONNECTED_500,SV2V_UNCONNECTED_501,SV2V_UNCONNECTED_502,
  SV2V_UNCONNECTED_503,SV2V_UNCONNECTED_504,SV2V_UNCONNECTED_505,
  SV2V_UNCONNECTED_506,SV2V_UNCONNECTED_507,SV2V_UNCONNECTED_508,
  SV2V_UNCONNECTED_509,SV2V_UNCONNECTED_510,SV2V_UNCONNECTED_511,
  SV2V_UNCONNECTED_512,SV2V_UNCONNECTED_513,SV2V_UNCONNECTED_514,SV2V_UNCONNECTED_515,
  SV2V_UNCONNECTED_516,SV2V_UNCONNECTED_517,SV2V_UNCONNECTED_518,
  SV2V_UNCONNECTED_519,SV2V_UNCONNECTED_520,SV2V_UNCONNECTED_521,
  SV2V_UNCONNECTED_522,SV2V_UNCONNECTED_523,SV2V_UNCONNECTED_524,
  SV2V_UNCONNECTED_525,SV2V_UNCONNECTED_526,SV2V_UNCONNECTED_527,
  SV2V_UNCONNECTED_528,SV2V_UNCONNECTED_529,SV2V_UNCONNECTED_530,SV2V_UNCONNECTED_531,
  SV2V_UNCONNECTED_532,SV2V_UNCONNECTED_533,SV2V_UNCONNECTED_534,
  SV2V_UNCONNECTED_535,SV2V_UNCONNECTED_536,SV2V_UNCONNECTED_537,
  SV2V_UNCONNECTED_538,SV2V_UNCONNECTED_539,SV2V_UNCONNECTED_540,
  SV2V_UNCONNECTED_541,SV2V_UNCONNECTED_542,SV2V_UNCONNECTED_543,
  SV2V_UNCONNECTED_544,SV2V_UNCONNECTED_545,SV2V_UNCONNECTED_546,SV2V_UNCONNECTED_547,
  SV2V_UNCONNECTED_548,SV2V_UNCONNECTED_549,SV2V_UNCONNECTED_550,
  SV2V_UNCONNECTED_551,SV2V_UNCONNECTED_552,SV2V_UNCONNECTED_553,
  SV2V_UNCONNECTED_554,SV2V_UNCONNECTED_555,SV2V_UNCONNECTED_556,
  SV2V_UNCONNECTED_557,SV2V_UNCONNECTED_558,SV2V_UNCONNECTED_559,
  SV2V_UNCONNECTED_560,SV2V_UNCONNECTED_561,SV2V_UNCONNECTED_562,SV2V_UNCONNECTED_563,
  SV2V_UNCONNECTED_564,SV2V_UNCONNECTED_565,SV2V_UNCONNECTED_566,
  SV2V_UNCONNECTED_567,SV2V_UNCONNECTED_568,SV2V_UNCONNECTED_569,
  SV2V_UNCONNECTED_570,SV2V_UNCONNECTED_571,SV2V_UNCONNECTED_572,
  SV2V_UNCONNECTED_573,SV2V_UNCONNECTED_574,SV2V_UNCONNECTED_575,
  SV2V_UNCONNECTED_576,SV2V_UNCONNECTED_577,SV2V_UNCONNECTED_578,SV2V_UNCONNECTED_579,
  SV2V_UNCONNECTED_580,SV2V_UNCONNECTED_581,SV2V_UNCONNECTED_582,
  SV2V_UNCONNECTED_583,SV2V_UNCONNECTED_584,SV2V_UNCONNECTED_585,
  SV2V_UNCONNECTED_586,SV2V_UNCONNECTED_587,SV2V_UNCONNECTED_588,
  SV2V_UNCONNECTED_589,SV2V_UNCONNECTED_590,SV2V_UNCONNECTED_591,
  SV2V_UNCONNECTED_592,SV2V_UNCONNECTED_593,SV2V_UNCONNECTED_594,SV2V_UNCONNECTED_595,
  SV2V_UNCONNECTED_596,SV2V_UNCONNECTED_597,SV2V_UNCONNECTED_598,
  SV2V_UNCONNECTED_599,SV2V_UNCONNECTED_600,SV2V_UNCONNECTED_601,
  SV2V_UNCONNECTED_602,SV2V_UNCONNECTED_603,SV2V_UNCONNECTED_604,
  SV2V_UNCONNECTED_605,SV2V_UNCONNECTED_606,SV2V_UNCONNECTED_607,
  SV2V_UNCONNECTED_608,SV2V_UNCONNECTED_609,SV2V_UNCONNECTED_610,SV2V_UNCONNECTED_611,
  SV2V_UNCONNECTED_612,SV2V_UNCONNECTED_613,SV2V_UNCONNECTED_614,
  SV2V_UNCONNECTED_615,SV2V_UNCONNECTED_616,SV2V_UNCONNECTED_617,
  SV2V_UNCONNECTED_618,SV2V_UNCONNECTED_619,SV2V_UNCONNECTED_620,
  SV2V_UNCONNECTED_621,SV2V_UNCONNECTED_622,SV2V_UNCONNECTED_623,
  SV2V_UNCONNECTED_624,SV2V_UNCONNECTED_625,SV2V_UNCONNECTED_626,SV2V_UNCONNECTED_627,
  SV2V_UNCONNECTED_628,SV2V_UNCONNECTED_629,SV2V_UNCONNECTED_630,
  SV2V_UNCONNECTED_631,SV2V_UNCONNECTED_632,SV2V_UNCONNECTED_633,
  SV2V_UNCONNECTED_634,SV2V_UNCONNECTED_635,SV2V_UNCONNECTED_636,
  SV2V_UNCONNECTED_637,SV2V_UNCONNECTED_638,SV2V_UNCONNECTED_639,
  SV2V_UNCONNECTED_640,SV2V_UNCONNECTED_641,SV2V_UNCONNECTED_642,SV2V_UNCONNECTED_643,
  SV2V_UNCONNECTED_644,SV2V_UNCONNECTED_645,SV2V_UNCONNECTED_646,
  SV2V_UNCONNECTED_647,SV2V_UNCONNECTED_648,SV2V_UNCONNECTED_649,
  SV2V_UNCONNECTED_650,SV2V_UNCONNECTED_651,SV2V_UNCONNECTED_652,
  SV2V_UNCONNECTED_653,SV2V_UNCONNECTED_654,SV2V_UNCONNECTED_655,
  SV2V_UNCONNECTED_656,SV2V_UNCONNECTED_657,SV2V_UNCONNECTED_658,SV2V_UNCONNECTED_659,
  SV2V_UNCONNECTED_660,SV2V_UNCONNECTED_661,SV2V_UNCONNECTED_662,
  SV2V_UNCONNECTED_663,SV2V_UNCONNECTED_664,SV2V_UNCONNECTED_665,
  SV2V_UNCONNECTED_666,SV2V_UNCONNECTED_667,SV2V_UNCONNECTED_668,
  SV2V_UNCONNECTED_669,SV2V_UNCONNECTED_670,SV2V_UNCONNECTED_671,
  SV2V_UNCONNECTED_672,SV2V_UNCONNECTED_673,SV2V_UNCONNECTED_674,SV2V_UNCONNECTED_675,
  SV2V_UNCONNECTED_676,SV2V_UNCONNECTED_677,SV2V_UNCONNECTED_678,
  SV2V_UNCONNECTED_679,SV2V_UNCONNECTED_680,SV2V_UNCONNECTED_681,
  SV2V_UNCONNECTED_682,SV2V_UNCONNECTED_683,SV2V_UNCONNECTED_684,
  SV2V_UNCONNECTED_685,SV2V_UNCONNECTED_686,SV2V_UNCONNECTED_687,
  SV2V_UNCONNECTED_688,SV2V_UNCONNECTED_689,SV2V_UNCONNECTED_690,SV2V_UNCONNECTED_691,
  SV2V_UNCONNECTED_692,SV2V_UNCONNECTED_693,SV2V_UNCONNECTED_694,
  SV2V_UNCONNECTED_695,SV2V_UNCONNECTED_696,SV2V_UNCONNECTED_697,
  SV2V_UNCONNECTED_698,SV2V_UNCONNECTED_699,SV2V_UNCONNECTED_700,
  SV2V_UNCONNECTED_701,SV2V_UNCONNECTED_702,SV2V_UNCONNECTED_703,
  SV2V_UNCONNECTED_704,SV2V_UNCONNECTED_705,SV2V_UNCONNECTED_706,SV2V_UNCONNECTED_707,
  SV2V_UNCONNECTED_708,SV2V_UNCONNECTED_709,SV2V_UNCONNECTED_710,
  SV2V_UNCONNECTED_711,SV2V_UNCONNECTED_712,SV2V_UNCONNECTED_713,
  SV2V_UNCONNECTED_714,SV2V_UNCONNECTED_715,SV2V_UNCONNECTED_716,
  SV2V_UNCONNECTED_717,SV2V_UNCONNECTED_718,SV2V_UNCONNECTED_719,
  SV2V_UNCONNECTED_720,SV2V_UNCONNECTED_721,SV2V_UNCONNECTED_722,SV2V_UNCONNECTED_723,
  SV2V_UNCONNECTED_724,SV2V_UNCONNECTED_725,SV2V_UNCONNECTED_726,
  SV2V_UNCONNECTED_727,SV2V_UNCONNECTED_728,SV2V_UNCONNECTED_729,
  SV2V_UNCONNECTED_730,SV2V_UNCONNECTED_731,SV2V_UNCONNECTED_732,
  SV2V_UNCONNECTED_733,SV2V_UNCONNECTED_734,SV2V_UNCONNECTED_735,
  SV2V_UNCONNECTED_736,SV2V_UNCONNECTED_737,SV2V_UNCONNECTED_738,SV2V_UNCONNECTED_739,
  SV2V_UNCONNECTED_740,SV2V_UNCONNECTED_741,SV2V_UNCONNECTED_742,
  SV2V_UNCONNECTED_743,SV2V_UNCONNECTED_744,SV2V_UNCONNECTED_745,
  SV2V_UNCONNECTED_746,SV2V_UNCONNECTED_747,SV2V_UNCONNECTED_748,
  SV2V_UNCONNECTED_749,SV2V_UNCONNECTED_750,SV2V_UNCONNECTED_751,
  SV2V_UNCONNECTED_752,SV2V_UNCONNECTED_753,SV2V_UNCONNECTED_754,SV2V_UNCONNECTED_755,
  SV2V_UNCONNECTED_756,SV2V_UNCONNECTED_757,SV2V_UNCONNECTED_758,
  SV2V_UNCONNECTED_759,SV2V_UNCONNECTED_760,SV2V_UNCONNECTED_761,
  SV2V_UNCONNECTED_762,SV2V_UNCONNECTED_763,SV2V_UNCONNECTED_764,
  SV2V_UNCONNECTED_765,SV2V_UNCONNECTED_766,SV2V_UNCONNECTED_767,
  SV2V_UNCONNECTED_768,SV2V_UNCONNECTED_769,SV2V_UNCONNECTED_770,SV2V_UNCONNECTED_771,
  SV2V_UNCONNECTED_772,SV2V_UNCONNECTED_773,SV2V_UNCONNECTED_774,
  SV2V_UNCONNECTED_775,SV2V_UNCONNECTED_776,SV2V_UNCONNECTED_777,
  SV2V_UNCONNECTED_778,SV2V_UNCONNECTED_779,SV2V_UNCONNECTED_780,
  SV2V_UNCONNECTED_781,SV2V_UNCONNECTED_782,SV2V_UNCONNECTED_783,
  SV2V_UNCONNECTED_784,SV2V_UNCONNECTED_785,SV2V_UNCONNECTED_786,SV2V_UNCONNECTED_787,
  SV2V_UNCONNECTED_788,SV2V_UNCONNECTED_789,SV2V_UNCONNECTED_790,
  SV2V_UNCONNECTED_791,SV2V_UNCONNECTED_792,SV2V_UNCONNECTED_793,
  SV2V_UNCONNECTED_794,SV2V_UNCONNECTED_795,SV2V_UNCONNECTED_796,
  SV2V_UNCONNECTED_797,SV2V_UNCONNECTED_798,SV2V_UNCONNECTED_799,
  SV2V_UNCONNECTED_800,SV2V_UNCONNECTED_801,SV2V_UNCONNECTED_802,SV2V_UNCONNECTED_803,
  SV2V_UNCONNECTED_804,SV2V_UNCONNECTED_805,SV2V_UNCONNECTED_806,
  SV2V_UNCONNECTED_807,SV2V_UNCONNECTED_808,SV2V_UNCONNECTED_809,
  SV2V_UNCONNECTED_810,SV2V_UNCONNECTED_811,SV2V_UNCONNECTED_812,
  SV2V_UNCONNECTED_813,SV2V_UNCONNECTED_814,SV2V_UNCONNECTED_815,
  SV2V_UNCONNECTED_816,SV2V_UNCONNECTED_817,SV2V_UNCONNECTED_818,SV2V_UNCONNECTED_819,
  SV2V_UNCONNECTED_820,SV2V_UNCONNECTED_821,SV2V_UNCONNECTED_822,
  SV2V_UNCONNECTED_823,SV2V_UNCONNECTED_824,SV2V_UNCONNECTED_825,
  SV2V_UNCONNECTED_826,SV2V_UNCONNECTED_827,SV2V_UNCONNECTED_828,
  SV2V_UNCONNECTED_829,SV2V_UNCONNECTED_830,SV2V_UNCONNECTED_831,
  SV2V_UNCONNECTED_832,SV2V_UNCONNECTED_833,SV2V_UNCONNECTED_834,SV2V_UNCONNECTED_835,
  SV2V_UNCONNECTED_836,SV2V_UNCONNECTED_837,SV2V_UNCONNECTED_838,
  SV2V_UNCONNECTED_839,SV2V_UNCONNECTED_840,SV2V_UNCONNECTED_841,
  SV2V_UNCONNECTED_842,SV2V_UNCONNECTED_843,SV2V_UNCONNECTED_844,
  SV2V_UNCONNECTED_845,SV2V_UNCONNECTED_846,SV2V_UNCONNECTED_847,
  SV2V_UNCONNECTED_848,SV2V_UNCONNECTED_849,SV2V_UNCONNECTED_850,SV2V_UNCONNECTED_851,
  SV2V_UNCONNECTED_852,SV2V_UNCONNECTED_853,SV2V_UNCONNECTED_854,
  SV2V_UNCONNECTED_855,SV2V_UNCONNECTED_856,SV2V_UNCONNECTED_857,
  SV2V_UNCONNECTED_858,SV2V_UNCONNECTED_859,SV2V_UNCONNECTED_860,
  SV2V_UNCONNECTED_861,SV2V_UNCONNECTED_862,SV2V_UNCONNECTED_863,
  SV2V_UNCONNECTED_864,SV2V_UNCONNECTED_865,SV2V_UNCONNECTED_866,SV2V_UNCONNECTED_867,
  SV2V_UNCONNECTED_868,SV2V_UNCONNECTED_869,SV2V_UNCONNECTED_870,
  SV2V_UNCONNECTED_871,SV2V_UNCONNECTED_872,SV2V_UNCONNECTED_873,
  SV2V_UNCONNECTED_874,SV2V_UNCONNECTED_875,SV2V_UNCONNECTED_876,
  SV2V_UNCONNECTED_877,SV2V_UNCONNECTED_878,SV2V_UNCONNECTED_879,
  SV2V_UNCONNECTED_880,SV2V_UNCONNECTED_881,SV2V_UNCONNECTED_882,SV2V_UNCONNECTED_883,
  SV2V_UNCONNECTED_884,SV2V_UNCONNECTED_885,SV2V_UNCONNECTED_886,
  SV2V_UNCONNECTED_887,SV2V_UNCONNECTED_888,SV2V_UNCONNECTED_889,
  SV2V_UNCONNECTED_890,SV2V_UNCONNECTED_891,SV2V_UNCONNECTED_892,
  SV2V_UNCONNECTED_893,SV2V_UNCONNECTED_894,SV2V_UNCONNECTED_895,
  SV2V_UNCONNECTED_896,SV2V_UNCONNECTED_897,SV2V_UNCONNECTED_898,SV2V_UNCONNECTED_899,
  SV2V_UNCONNECTED_900,SV2V_UNCONNECTED_901,SV2V_UNCONNECTED_902,
  SV2V_UNCONNECTED_903,SV2V_UNCONNECTED_904,SV2V_UNCONNECTED_905,
  SV2V_UNCONNECTED_906,SV2V_UNCONNECTED_907,SV2V_UNCONNECTED_908,
  SV2V_UNCONNECTED_909;
  wire [27:0] T4,T212,T216,T218;
  wire [25:0] sigX3,T373,T27,T499,T250,T237,T238,roundUp_sigY3,T239,T242,T272,T251,T273;
  wire [0:0] roundMask,T374,T489,T488,T504;
  wire [26:26] T77;
  wire [26:2] T6,T503;
  wire [24:0] T9;
  wire [7:0] T12,T89;
  wire [15:0] T13,T82,T125,T207,T208;
  wire [9:0] T15,sExpX3_13,T280,T233,T234,T283,T281,T284;
  wire [10:10] sExpX3;
  wire [6:0] T375,CDom_estNormDist,T16,sExpY;
  wire [5:0] T376,T378,T379,T380,T381,T382,T383,T384,T385,T386,T387,T388,T389,T390,T391,T392,
  T393,T394;
  wire [3:0] T411,T412,T413,T414,T415,T416,T417,T418,T88,normTo2ShiftDist;
  wire [2:0] T419,T420,T421,T422,T232;
  wire [1:0] T423,T424,T87,T501,T236;
  wire [49:1] T18;
  wire [50:49] T21;
  wire [74:51] sigSum;
  wire [7:7] T34,T37,T107,T110,T348;
  wire [6:6] T35,T108,T341,T345;
  wire [7:6] T38,T41,T111,T114;
  wire [5:4] T39,T112;
  wire [15:15] T53,T56,T148;
  wire [14:14] T54;
  wire [15:14] T57,T60;
  wire [13:12] T58;
  wire [15:12] T61,T64;
  wire [11:8] T62;
  wire [15:8] absSigSumExtraMask;
  wire [42:16] cFirstNormAbsSigSum;
  wire [42:0] T192,notCDom_neg_cFirstNormAbsSigSum,T200,T193;
  wire [41:0] T487,CDom_firstNormAbsSigSum,notCDom_pos_firstNormAbsSigSum,T146,T127,T162,T154,
  T172,T163,T182,T173;
  wire [31:31] T128;
  wire [17:0] T141;
  wire [74:18] notSigSum;
  wire [41:41] T491,T492,T493,T494;
  wire [26:0] T498;
  wire [23:0] sigY3;
  wire [22:0] T318,T322,fractY;
  wire [22:22] T313,T319;
  wire [8:0] T333,T338,T340,T343,T346,T344,T349,T347,T352,T350,T353;
  wire [8:8] T332,T334,T339,T351,T354;
  assign io_exceptionFlags[3] = 1'b0;
  assign { SV2V_UNCONNECTED_1, SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, sigX3_27, T374[0:0], sigX3[25:1] } = { cFirstNormAbsSigSum, T125[15:1] } >> normTo2ShiftDist;
  assign T228 = sExpX3_13 <= { 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T501 };
  assign sigX3Shift1 = { sigX3_27, T374[0:0] } == 1'b0;
  assign isZeroY = { sigX3_27, T374[0:0], sigX3[25:25] } == 1'b0;
  assign T328 = { T232[1:0], sExpY } < { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 };
  assign N197 = io_fromPreMul_highExpB[1] | io_fromPreMul_highExpB[2];
  assign N198 = io_fromPreMul_highExpB[0] | N197;
  assign N199 = ~N198;
  assign N200 = io_fromPreMul_highExpA[1] | io_fromPreMul_highExpA[2];
  assign N201 = io_fromPreMul_highExpA[0] | N200;
  assign N202 = ~N201;
  assign N203 = ~T232[1];
  assign N204 = ~T232[0];
  assign N205 = N203 | T232[2];
  assign N206 = N204 | N205;
  assign N207 = ~N206;
  assign N208 = io_fromPreMul_highExpC[1] & io_fromPreMul_highExpC[2];
  assign N209 = io_fromPreMul_highExpA[1] & io_fromPreMul_highExpA[2];
  assign N210 = io_fromPreMul_highExpB[1] & io_fromPreMul_highExpB[2];
  assign N211 = T236[0] | T236[1];
  assign N212 = ~N211;
  assign N213 = T216[26] | T216[27];
  assign N214 = T216[25] | N213;
  assign N215 = T216[24] | N214;
  assign N216 = T216[23] | N215;
  assign N217 = T216[22] | N216;
  assign N218 = T216[21] | N217;
  assign N219 = T216[20] | N218;
  assign N220 = T216[19] | N219;
  assign N221 = T216[18] | N220;
  assign N222 = T216[17] | N221;
  assign N223 = T216[16] | N222;
  assign N224 = T216[15] | N223;
  assign N225 = T216[14] | N224;
  assign N226 = T216[13] | N225;
  assign N227 = T216[12] | N226;
  assign N228 = T216[11] | N227;
  assign N229 = T216[10] | N228;
  assign N230 = T216[9] | N229;
  assign N231 = T216[8] | N230;
  assign N232 = T216[7] | N231;
  assign N233 = T216[6] | N232;
  assign N234 = T216[5] | N233;
  assign N235 = T216[4] | N234;
  assign N236 = T216[3] | N235;
  assign N237 = T216[2] | N236;
  assign N238 = T216[1] | N237;
  assign N239 = T216[0] | N238;
  assign N240 = ~N239;
  assign N241 = T212[26] | T212[27];
  assign N242 = T212[25] | N241;
  assign N243 = T212[24] | N242;
  assign N244 = T212[23] | N243;
  assign N245 = T212[22] | N244;
  assign N246 = T212[21] | N245;
  assign N247 = T212[20] | N246;
  assign N248 = T212[19] | N247;
  assign N249 = T212[18] | N248;
  assign N250 = T212[17] | N249;
  assign N251 = T212[16] | N250;
  assign N252 = T212[15] | N251;
  assign N253 = T212[14] | N252;
  assign N254 = T212[13] | N253;
  assign N255 = T212[12] | N254;
  assign N256 = T212[11] | N255;
  assign N257 = T212[10] | N256;
  assign N258 = T212[9] | N257;
  assign N259 = T212[8] | N258;
  assign N260 = T212[7] | N259;
  assign N261 = T212[6] | N260;
  assign N262 = T212[5] | N261;
  assign N263 = T212[4] | N262;
  assign N264 = T212[3] | N263;
  assign N265 = T212[2] | N264;
  assign N266 = T212[1] | N265;
  assign N267 = T212[0] | N266;
  assign N268 = T4[26] | T4[27];
  assign N269 = T4[25] | N268;
  assign N270 = T4[24] | N269;
  assign N271 = T4[23] | N270;
  assign N272 = T4[22] | N271;
  assign N273 = T4[21] | N272;
  assign N274 = T4[20] | N273;
  assign N275 = T4[19] | N274;
  assign N276 = T4[18] | N275;
  assign N277 = T4[17] | N276;
  assign N278 = T4[16] | N277;
  assign N279 = T4[15] | N278;
  assign N280 = T4[14] | N279;
  assign N281 = T4[13] | N280;
  assign N282 = T4[12] | N281;
  assign N283 = T4[11] | N282;
  assign N284 = T4[10] | N283;
  assign N285 = T4[9] | N284;
  assign N286 = T4[8] | N285;
  assign N287 = T4[7] | N286;
  assign N288 = T4[6] | N287;
  assign N289 = T4[5] | N288;
  assign N290 = T4[4] | N289;
  assign N291 = T4[3] | N290;
  assign N292 = T4[2] | N291;
  assign N293 = T4[1] | N292;
  assign N294 = T4[0] | N293;
  assign N295 = io_fromPreMul_roundingMode[0] | io_fromPreMul_roundingMode[1];
  assign N296 = ~N295;
  assign N297 = io_fromPreMul_roundingMode[0] & io_fromPreMul_roundingMode[1];
  assign N298 = T207[14] | T207[15];
  assign N299 = T207[13] | N298;
  assign N300 = T207[12] | N299;
  assign N301 = T207[11] | N300;
  assign N302 = T207[10] | N301;
  assign N303 = T207[9] | N302;
  assign N304 = T207[8] | N303;
  assign N305 = T207[7] | N304;
  assign N306 = T207[6] | N305;
  assign N307 = T207[5] | N306;
  assign N308 = T207[4] | N307;
  assign N309 = T207[3] | N308;
  assign N310 = T207[2] | N309;
  assign N311 = T207[1] | N310;
  assign N312 = T207[0] | N311;
  assign N313 = ~N312;
  assign N314 = T82[14] | T82[15];
  assign N315 = T82[13] | N314;
  assign N316 = T82[12] | N315;
  assign N317 = T82[11] | N316;
  assign N318 = T82[10] | N317;
  assign N319 = T82[9] | N318;
  assign N320 = T82[8] | N319;
  assign N321 = T82[7] | N320;
  assign N322 = T82[6] | N321;
  assign N323 = T82[5] | N322;
  assign N324 = T82[4] | N323;
  assign N325 = T82[3] | N324;
  assign N326 = T82[2] | N325;
  assign N327 = T82[1] | N326;
  assign N328 = T82[0] | N327;
  assign N329 = ~io_fromPreMul_roundingMode[1];
  assign N330 = io_fromPreMul_roundingMode[0] | N329;
  assign N331 = ~N330;
  assign N332 = io_fromPreMul_highExpC[1] | io_fromPreMul_highExpC[2];
  assign N333 = io_fromPreMul_highExpC[0] | N332;
  assign N334 = ~N333;
  assign { SV2V_UNCONNECTED_16, absSigSumExtraMask_1, T87, T88, T89 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> normTo2ShiftDist;
  assign { SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, SV2V_UNCONNECTED_32, SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, SV2V_UNCONNECTED_49, SV2V_UNCONNECTED_50, SV2V_UNCONNECTED_51, SV2V_UNCONNECTED_52, SV2V_UNCONNECTED_53, SV2V_UNCONNECTED_54, SV2V_UNCONNECTED_55, SV2V_UNCONNECTED_56, SV2V_UNCONNECTED_57, SV2V_UNCONNECTED_58, SV2V_UNCONNECTED_59, SV2V_UNCONNECTED_60, SV2V_UNCONNECTED_61, SV2V_UNCONNECTED_62, SV2V_UNCONNECTED_63, SV2V_UNCONNECTED_64, SV2V_UNCONNECTED_65, SV2V_UNCONNECTED_66, SV2V_UNCONNECTED_67, SV2V_UNCONNECTED_68, SV2V_UNCONNECTED_69, SV2V_UNCONNECTED_70, SV2V_UNCONNECTED_71, SV2V_UNCONNECTED_72, SV2V_UNCONNECTED_73, SV2V_UNCONNECTED_74, SV2V_UNCONNECTED_75, SV2V_UNCONNECTED_76, SV2V_UNCONNECTED_77, SV2V_UNCONNECTED_78, SV2V_UNCONNECTED_79, SV2V_UNCONNECTED_80, SV2V_UNCONNECTED_81, SV2V_UNCONNECTED_82, SV2V_UNCONNECTED_83, SV2V_UNCONNECTED_84, SV2V_UNCONNECTED_85, SV2V_UNCONNECTED_86, SV2V_UNCONNECTED_87, SV2V_UNCONNECTED_88, SV2V_UNCONNECTED_89, SV2V_UNCONNECTED_90, SV2V_UNCONNECTED_91, SV2V_UNCONNECTED_92, SV2V_UNCONNECTED_93, SV2V_UNCONNECTED_94, SV2V_UNCONNECTED_95, SV2V_UNCONNECTED_96, SV2V_UNCONNECTED_97, SV2V_UNCONNECTED_98, SV2V_UNCONNECTED_99, SV2V_UNCONNECTED_100, SV2V_UNCONNECTED_101, SV2V_UNCONNECTED_102, SV2V_UNCONNECTED_103, SV2V_UNCONNECTED_104, SV2V_UNCONNECTED_105, SV2V_UNCONNECTED_106, SV2V_UNCONNECTED_107, SV2V_UNCONNECTED_108, SV2V_UNCONNECTED_109, SV2V_UNCONNECTED_110, SV2V_UNCONNECTED_111, SV2V_UNCONNECTED_112, SV2V_UNCONNECTED_113, SV2V_UNCONNECTED_114, SV2V_UNCONNECTED_115, SV2V_UNCONNECTED_116, SV2V_UNCONNECTED_117, SV2V_UNCONNECTED_118, SV2V_UNCONNECTED_119, SV2V_UNCONNECTED_120, SV2V_UNCONNECTED_121, SV2V_UNCONNECTED_122, SV2V_UNCONNECTED_123, SV2V_UNCONNECTED_124, SV2V_UNCONNECTED_125, SV2V_UNCONNECTED_126, SV2V_UNCONNECTED_127, SV2V_UNCONNECTED_128, SV2V_UNCONNECTED_129, SV2V_UNCONNECTED_130, SV2V_UNCONNECTED_131, SV2V_UNCONNECTED_132, SV2V_UNCONNECTED_133, SV2V_UNCONNECTED_134, SV2V_UNCONNECTED_135, SV2V_UNCONNECTED_136, SV2V_UNCONNECTED_137, SV2V_UNCONNECTED_138, SV2V_UNCONNECTED_139, SV2V_UNCONNECTED_140, SV2V_UNCONNECTED_141, SV2V_UNCONNECTED_142, SV2V_UNCONNECTED_143, SV2V_UNCONNECTED_144, SV2V_UNCONNECTED_145, SV2V_UNCONNECTED_146, SV2V_UNCONNECTED_147, SV2V_UNCONNECTED_148, SV2V_UNCONNECTED_149, SV2V_UNCONNECTED_150, SV2V_UNCONNECTED_151, SV2V_UNCONNECTED_152, SV2V_UNCONNECTED_153, SV2V_UNCONNECTED_154, SV2V_UNCONNECTED_155, SV2V_UNCONNECTED_156, SV2V_UNCONNECTED_157, SV2V_UNCONNECTED_158, SV2V_UNCONNECTED_159, SV2V_UNCONNECTED_160, SV2V_UNCONNECTED_161, SV2V_UNCONNECTED_162, SV2V_UNCONNECTED_163, SV2V_UNCONNECTED_164, SV2V_UNCONNECTED_165, SV2V_UNCONNECTED_166, SV2V_UNCONNECTED_167, SV2V_UNCONNECTED_168, SV2V_UNCONNECTED_169, SV2V_UNCONNECTED_170, SV2V_UNCONNECTED_171, SV2V_UNCONNECTED_172, SV2V_UNCONNECTED_173, SV2V_UNCONNECTED_174, SV2V_UNCONNECTED_175, SV2V_UNCONNECTED_176, SV2V_UNCONNECTED_177, SV2V_UNCONNECTED_178, SV2V_UNCONNECTED_179, SV2V_UNCONNECTED_180, SV2V_UNCONNECTED_181, SV2V_UNCONNECTED_182, SV2V_UNCONNECTED_183, SV2V_UNCONNECTED_184, SV2V_UNCONNECTED_185, SV2V_UNCONNECTED_186, SV2V_UNCONNECTED_187, SV2V_UNCONNECTED_188, SV2V_UNCONNECTED_189, SV2V_UNCONNECTED_190, SV2V_UNCONNECTED_191, SV2V_UNCONNECTED_192, SV2V_UNCONNECTED_193, SV2V_UNCONNECTED_194, SV2V_UNCONNECTED_195, SV2V_UNCONNECTED_196, SV2V_UNCONNECTED_197, SV2V_UNCONNECTED_198, SV2V_UNCONNECTED_199, SV2V_UNCONNECTED_200, SV2V_UNCONNECTED_201, SV2V_UNCONNECTED_202, SV2V_UNCONNECTED_203, SV2V_UNCONNECTED_204, SV2V_UNCONNECTED_205, SV2V_UNCONNECTED_206, SV2V_UNCONNECTED_207, SV2V_UNCONNECTED_208, SV2V_UNCONNECTED_209, SV2V_UNCONNECTED_210, SV2V_UNCONNECTED_211, SV2V_UNCONNECTED_212, SV2V_UNCONNECTED_213, SV2V_UNCONNECTED_214, SV2V_UNCONNECTED_215, SV2V_UNCONNECTED_216, SV2V_UNCONNECTED_217, SV2V_UNCONNECTED_218, SV2V_UNCONNECTED_219, SV2V_UNCONNECTED_220, SV2V_UNCONNECTED_221, SV2V_UNCONNECTED_222, SV2V_UNCONNECTED_223, SV2V_UNCONNECTED_224, SV2V_UNCONNECTED_225, SV2V_UNCONNECTED_226, SV2V_UNCONNECTED_227, SV2V_UNCONNECTED_228, SV2V_UNCONNECTED_229, SV2V_UNCONNECTED_230, SV2V_UNCONNECTED_231, SV2V_UNCONNECTED_232, SV2V_UNCONNECTED_233, SV2V_UNCONNECTED_234, SV2V_UNCONNECTED_235, SV2V_UNCONNECTED_236, SV2V_UNCONNECTED_237, SV2V_UNCONNECTED_238, SV2V_UNCONNECTED_239, SV2V_UNCONNECTED_240, SV2V_UNCONNECTED_241, SV2V_UNCONNECTED_242, SV2V_UNCONNECTED_243, SV2V_UNCONNECTED_244, SV2V_UNCONNECTED_245, SV2V_UNCONNECTED_246, SV2V_UNCONNECTED_247, SV2V_UNCONNECTED_248, SV2V_UNCONNECTED_249, SV2V_UNCONNECTED_250, SV2V_UNCONNECTED_251, SV2V_UNCONNECTED_252, SV2V_UNCONNECTED_253, SV2V_UNCONNECTED_254, SV2V_UNCONNECTED_255, SV2V_UNCONNECTED_256, SV2V_UNCONNECTED_257, SV2V_UNCONNECTED_258, SV2V_UNCONNECTED_259, SV2V_UNCONNECTED_260, SV2V_UNCONNECTED_261, SV2V_UNCONNECTED_262, SV2V_UNCONNECTED_263, SV2V_UNCONNECTED_264, SV2V_UNCONNECTED_265, SV2V_UNCONNECTED_266, SV2V_UNCONNECTED_267, SV2V_UNCONNECTED_268, SV2V_UNCONNECTED_269, SV2V_UNCONNECTED_270, SV2V_UNCONNECTED_271, SV2V_UNCONNECTED_272, SV2V_UNCONNECTED_273, SV2V_UNCONNECTED_274, SV2V_UNCONNECTED_275, SV2V_UNCONNECTED_276, SV2V_UNCONNECTED_277, SV2V_UNCONNECTED_278, SV2V_UNCONNECTED_279, SV2V_UNCONNECTED_280, SV2V_UNCONNECTED_281, SV2V_UNCONNECTED_282, SV2V_UNCONNECTED_283, SV2V_UNCONNECTED_284, SV2V_UNCONNECTED_285, SV2V_UNCONNECTED_286, SV2V_UNCONNECTED_287, SV2V_UNCONNECTED_288, SV2V_UNCONNECTED_289, SV2V_UNCONNECTED_290, SV2V_UNCONNECTED_291, SV2V_UNCONNECTED_292, SV2V_UNCONNECTED_293, SV2V_UNCONNECTED_294, SV2V_UNCONNECTED_295, SV2V_UNCONNECTED_296, SV2V_UNCONNECTED_297, SV2V_UNCONNECTED_298, SV2V_UNCONNECTED_299, SV2V_UNCONNECTED_300, SV2V_UNCONNECTED_301, SV2V_UNCONNECTED_302, SV2V_UNCONNECTED_303, SV2V_UNCONNECTED_304, SV2V_UNCONNECTED_305, SV2V_UNCONNECTED_306, SV2V_UNCONNECTED_307, SV2V_UNCONNECTED_308, SV2V_UNCONNECTED_309, SV2V_UNCONNECTED_310, SV2V_UNCONNECTED_311, SV2V_UNCONNECTED_312, SV2V_UNCONNECTED_313, SV2V_UNCONNECTED_314, SV2V_UNCONNECTED_315, SV2V_UNCONNECTED_316, SV2V_UNCONNECTED_317, SV2V_UNCONNECTED_318, SV2V_UNCONNECTED_319, SV2V_UNCONNECTED_320, SV2V_UNCONNECTED_321, SV2V_UNCONNECTED_322, SV2V_UNCONNECTED_323, SV2V_UNCONNECTED_324, SV2V_UNCONNECTED_325, SV2V_UNCONNECTED_326, SV2V_UNCONNECTED_327, SV2V_UNCONNECTED_328, SV2V_UNCONNECTED_329, SV2V_UNCONNECTED_330, SV2V_UNCONNECTED_331, SV2V_UNCONNECTED_332, SV2V_UNCONNECTED_333, SV2V_UNCONNECTED_334, SV2V_UNCONNECTED_335, SV2V_UNCONNECTED_336, SV2V_UNCONNECTED_337, SV2V_UNCONNECTED_338, SV2V_UNCONNECTED_339, SV2V_UNCONNECTED_340, SV2V_UNCONNECTED_341, SV2V_UNCONNECTED_342, SV2V_UNCONNECTED_343, SV2V_UNCONNECTED_344, SV2V_UNCONNECTED_345, SV2V_UNCONNECTED_346, SV2V_UNCONNECTED_347, SV2V_UNCONNECTED_348, SV2V_UNCONNECTED_349, SV2V_UNCONNECTED_350, SV2V_UNCONNECTED_351, SV2V_UNCONNECTED_352, SV2V_UNCONNECTED_353, SV2V_UNCONNECTED_354, SV2V_UNCONNECTED_355, SV2V_UNCONNECTED_356, SV2V_UNCONNECTED_357, SV2V_UNCONNECTED_358, SV2V_UNCONNECTED_359, SV2V_UNCONNECTED_360, SV2V_UNCONNECTED_361, SV2V_UNCONNECTED_362, SV2V_UNCONNECTED_363, SV2V_UNCONNECTED_364, SV2V_UNCONNECTED_365, SV2V_UNCONNECTED_366, SV2V_UNCONNECTED_367, SV2V_UNCONNECTED_368, SV2V_UNCONNECTED_369, SV2V_UNCONNECTED_370, SV2V_UNCONNECTED_371, SV2V_UNCONNECTED_372, SV2V_UNCONNECTED_373, SV2V_UNCONNECTED_374, SV2V_UNCONNECTED_375, SV2V_UNCONNECTED_376, SV2V_UNCONNECTED_377, SV2V_UNCONNECTED_378, SV2V_UNCONNECTED_379, SV2V_UNCONNECTED_380, SV2V_UNCONNECTED_381, SV2V_UNCONNECTED_382, SV2V_UNCONNECTED_383, SV2V_UNCONNECTED_384, SV2V_UNCONNECTED_385, SV2V_UNCONNECTED_386, SV2V_UNCONNECTED_387, SV2V_UNCONNECTED_388, SV2V_UNCONNECTED_389, SV2V_UNCONNECTED_390, SV2V_UNCONNECTED_391, SV2V_UNCONNECTED_392, SV2V_UNCONNECTED_393, SV2V_UNCONNECTED_394, SV2V_UNCONNECTED_395, SV2V_UNCONNECTED_396, SV2V_UNCONNECTED_397, SV2V_UNCONNECTED_398, SV2V_UNCONNECTED_399, SV2V_UNCONNECTED_400, SV2V_UNCONNECTED_401, SV2V_UNCONNECTED_402, SV2V_UNCONNECTED_403, SV2V_UNCONNECTED_404, SV2V_UNCONNECTED_405, SV2V_UNCONNECTED_406, SV2V_UNCONNECTED_407, SV2V_UNCONNECTED_408, SV2V_UNCONNECTED_409, SV2V_UNCONNECTED_410, SV2V_UNCONNECTED_411, SV2V_UNCONNECTED_412, SV2V_UNCONNECTED_413, SV2V_UNCONNECTED_414, SV2V_UNCONNECTED_415, SV2V_UNCONNECTED_416, SV2V_UNCONNECTED_417, SV2V_UNCONNECTED_418, SV2V_UNCONNECTED_419, SV2V_UNCONNECTED_420, SV2V_UNCONNECTED_421, SV2V_UNCONNECTED_422, SV2V_UNCONNECTED_423, SV2V_UNCONNECTED_424, SV2V_UNCONNECTED_425, SV2V_UNCONNECTED_426, SV2V_UNCONNECTED_427, SV2V_UNCONNECTED_428, SV2V_UNCONNECTED_429, SV2V_UNCONNECTED_430, SV2V_UNCONNECTED_431, SV2V_UNCONNECTED_432, SV2V_UNCONNECTED_433, SV2V_UNCONNECTED_434, SV2V_UNCONNECTED_435, SV2V_UNCONNECTED_436, SV2V_UNCONNECTED_437, SV2V_UNCONNECTED_438, SV2V_UNCONNECTED_439, SV2V_UNCONNECTED_440, SV2V_UNCONNECTED_441, SV2V_UNCONNECTED_442, SV2V_UNCONNECTED_443, SV2V_UNCONNECTED_444, SV2V_UNCONNECTED_445, SV2V_UNCONNECTED_446, SV2V_UNCONNECTED_447, SV2V_UNCONNECTED_448, SV2V_UNCONNECTED_449, SV2V_UNCONNECTED_450, SV2V_UNCONNECTED_451, SV2V_UNCONNECTED_452, SV2V_UNCONNECTED_453, SV2V_UNCONNECTED_454, SV2V_UNCONNECTED_455, SV2V_UNCONNECTED_456, SV2V_UNCONNECTED_457, SV2V_UNCONNECTED_458, SV2V_UNCONNECTED_459, SV2V_UNCONNECTED_460, SV2V_UNCONNECTED_461, SV2V_UNCONNECTED_462, SV2V_UNCONNECTED_463, SV2V_UNCONNECTED_464, SV2V_UNCONNECTED_465, SV2V_UNCONNECTED_466, SV2V_UNCONNECTED_467, SV2V_UNCONNECTED_468, SV2V_UNCONNECTED_469, SV2V_UNCONNECTED_470, SV2V_UNCONNECTED_471, SV2V_UNCONNECTED_472, SV2V_UNCONNECTED_473, SV2V_UNCONNECTED_474, SV2V_UNCONNECTED_475, SV2V_UNCONNECTED_476, SV2V_UNCONNECTED_477, SV2V_UNCONNECTED_478, SV2V_UNCONNECTED_479, SV2V_UNCONNECTED_480, SV2V_UNCONNECTED_481, SV2V_UNCONNECTED_482, SV2V_UNCONNECTED_483, SV2V_UNCONNECTED_484, SV2V_UNCONNECTED_485, SV2V_UNCONNECTED_486, SV2V_UNCONNECTED_487, SV2V_UNCONNECTED_488, SV2V_UNCONNECTED_489, SV2V_UNCONNECTED_490, SV2V_UNCONNECTED_491, SV2V_UNCONNECTED_492, SV2V_UNCONNECTED_493, SV2V_UNCONNECTED_494, SV2V_UNCONNECTED_495, SV2V_UNCONNECTED_496, SV2V_UNCONNECTED_497, SV2V_UNCONNECTED_498, SV2V_UNCONNECTED_499, SV2V_UNCONNECTED_500, SV2V_UNCONNECTED_501, SV2V_UNCONNECTED_502, SV2V_UNCONNECTED_503, SV2V_UNCONNECTED_504, SV2V_UNCONNECTED_505, SV2V_UNCONNECTED_506, SV2V_UNCONNECTED_507, SV2V_UNCONNECTED_508, SV2V_UNCONNECTED_509, SV2V_UNCONNECTED_510, SV2V_UNCONNECTED_511, SV2V_UNCONNECTED_512, SV2V_UNCONNECTED_513, SV2V_UNCONNECTED_514, SV2V_UNCONNECTED_515, SV2V_UNCONNECTED_516, SV2V_UNCONNECTED_517, SV2V_UNCONNECTED_518, SV2V_UNCONNECTED_519, SV2V_UNCONNECTED_520, SV2V_UNCONNECTED_521, SV2V_UNCONNECTED_522, SV2V_UNCONNECTED_523, SV2V_UNCONNECTED_524, SV2V_UNCONNECTED_525, SV2V_UNCONNECTED_526, SV2V_UNCONNECTED_527, SV2V_UNCONNECTED_528, SV2V_UNCONNECTED_529, SV2V_UNCONNECTED_530, SV2V_UNCONNECTED_531, SV2V_UNCONNECTED_532, SV2V_UNCONNECTED_533, SV2V_UNCONNECTED_534, SV2V_UNCONNECTED_535, SV2V_UNCONNECTED_536, SV2V_UNCONNECTED_537, SV2V_UNCONNECTED_538, SV2V_UNCONNECTED_539, SV2V_UNCONNECTED_540, SV2V_UNCONNECTED_541, SV2V_UNCONNECTED_542, SV2V_UNCONNECTED_543, SV2V_UNCONNECTED_544, SV2V_UNCONNECTED_545, SV2V_UNCONNECTED_546, SV2V_UNCONNECTED_547, SV2V_UNCONNECTED_548, SV2V_UNCONNECTED_549, SV2V_UNCONNECTED_550, SV2V_UNCONNECTED_551, SV2V_UNCONNECTED_552, SV2V_UNCONNECTED_553, SV2V_UNCONNECTED_554, SV2V_UNCONNECTED_555, SV2V_UNCONNECTED_556, SV2V_UNCONNECTED_557, SV2V_UNCONNECTED_558, SV2V_UNCONNECTED_559, SV2V_UNCONNECTED_560, SV2V_UNCONNECTED_561, SV2V_UNCONNECTED_562, SV2V_UNCONNECTED_563, SV2V_UNCONNECTED_564, SV2V_UNCONNECTED_565, SV2V_UNCONNECTED_566, SV2V_UNCONNECTED_567, SV2V_UNCONNECTED_568, SV2V_UNCONNECTED_569, SV2V_UNCONNECTED_570, SV2V_UNCONNECTED_571, SV2V_UNCONNECTED_572, SV2V_UNCONNECTED_573, SV2V_UNCONNECTED_574, SV2V_UNCONNECTED_575, SV2V_UNCONNECTED_576, SV2V_UNCONNECTED_577, SV2V_UNCONNECTED_578, SV2V_UNCONNECTED_579, SV2V_UNCONNECTED_580, SV2V_UNCONNECTED_581, SV2V_UNCONNECTED_582, SV2V_UNCONNECTED_583, SV2V_UNCONNECTED_584, SV2V_UNCONNECTED_585, SV2V_UNCONNECTED_586, SV2V_UNCONNECTED_587, SV2V_UNCONNECTED_588, SV2V_UNCONNECTED_589, SV2V_UNCONNECTED_590, SV2V_UNCONNECTED_591, SV2V_UNCONNECTED_592, SV2V_UNCONNECTED_593, SV2V_UNCONNECTED_594, SV2V_UNCONNECTED_595, SV2V_UNCONNECTED_596, SV2V_UNCONNECTED_597, SV2V_UNCONNECTED_598, SV2V_UNCONNECTED_599, SV2V_UNCONNECTED_600, SV2V_UNCONNECTED_601, SV2V_UNCONNECTED_602, SV2V_UNCONNECTED_603, SV2V_UNCONNECTED_604, SV2V_UNCONNECTED_605, SV2V_UNCONNECTED_606, SV2V_UNCONNECTED_607, SV2V_UNCONNECTED_608, SV2V_UNCONNECTED_609, SV2V_UNCONNECTED_610, SV2V_UNCONNECTED_611, SV2V_UNCONNECTED_612, SV2V_UNCONNECTED_613, SV2V_UNCONNECTED_614, SV2V_UNCONNECTED_615, SV2V_UNCONNECTED_616, SV2V_UNCONNECTED_617, SV2V_UNCONNECTED_618, SV2V_UNCONNECTED_619, SV2V_UNCONNECTED_620, SV2V_UNCONNECTED_621, SV2V_UNCONNECTED_622, SV2V_UNCONNECTED_623, SV2V_UNCONNECTED_624, SV2V_UNCONNECTED_625, SV2V_UNCONNECTED_626, SV2V_UNCONNECTED_627, SV2V_UNCONNECTED_628, SV2V_UNCONNECTED_629, SV2V_UNCONNECTED_630, SV2V_UNCONNECTED_631, SV2V_UNCONNECTED_632, SV2V_UNCONNECTED_633, SV2V_UNCONNECTED_634, SV2V_UNCONNECTED_635, SV2V_UNCONNECTED_636, SV2V_UNCONNECTED_637, SV2V_UNCONNECTED_638, SV2V_UNCONNECTED_639, SV2V_UNCONNECTED_640, SV2V_UNCONNECTED_641, SV2V_UNCONNECTED_642, SV2V_UNCONNECTED_643, SV2V_UNCONNECTED_644, SV2V_UNCONNECTED_645, SV2V_UNCONNECTED_646, SV2V_UNCONNECTED_647, SV2V_UNCONNECTED_648, SV2V_UNCONNECTED_649, SV2V_UNCONNECTED_650, SV2V_UNCONNECTED_651, SV2V_UNCONNECTED_652, SV2V_UNCONNECTED_653, SV2V_UNCONNECTED_654, SV2V_UNCONNECTED_655, SV2V_UNCONNECTED_656, SV2V_UNCONNECTED_657, SV2V_UNCONNECTED_658, SV2V_UNCONNECTED_659, SV2V_UNCONNECTED_660, SV2V_UNCONNECTED_661, SV2V_UNCONNECTED_662, SV2V_UNCONNECTED_663, SV2V_UNCONNECTED_664, SV2V_UNCONNECTED_665, SV2V_UNCONNECTED_666, SV2V_UNCONNECTED_667, SV2V_UNCONNECTED_668, SV2V_UNCONNECTED_669, SV2V_UNCONNECTED_670, SV2V_UNCONNECTED_671, SV2V_UNCONNECTED_672, SV2V_UNCONNECTED_673, SV2V_UNCONNECTED_674, SV2V_UNCONNECTED_675, SV2V_UNCONNECTED_676, SV2V_UNCONNECTED_677, SV2V_UNCONNECTED_678, SV2V_UNCONNECTED_679, SV2V_UNCONNECTED_680, SV2V_UNCONNECTED_681, SV2V_UNCONNECTED_682, SV2V_UNCONNECTED_683, SV2V_UNCONNECTED_684, SV2V_UNCONNECTED_685, SV2V_UNCONNECTED_686, SV2V_UNCONNECTED_687, SV2V_UNCONNECTED_688, SV2V_UNCONNECTED_689, SV2V_UNCONNECTED_690, SV2V_UNCONNECTED_691, SV2V_UNCONNECTED_692, SV2V_UNCONNECTED_693, SV2V_UNCONNECTED_694, SV2V_UNCONNECTED_695, SV2V_UNCONNECTED_696, SV2V_UNCONNECTED_697, SV2V_UNCONNECTED_698, SV2V_UNCONNECTED_699, SV2V_UNCONNECTED_700, SV2V_UNCONNECTED_701, SV2V_UNCONNECTED_702, SV2V_UNCONNECTED_703, SV2V_UNCONNECTED_704, SV2V_UNCONNECTED_705, SV2V_UNCONNECTED_706, SV2V_UNCONNECTED_707, SV2V_UNCONNECTED_708, SV2V_UNCONNECTED_709, SV2V_UNCONNECTED_710, SV2V_UNCONNECTED_711, SV2V_UNCONNECTED_712, SV2V_UNCONNECTED_713, SV2V_UNCONNECTED_714, SV2V_UNCONNECTED_715, SV2V_UNCONNECTED_716, SV2V_UNCONNECTED_717, SV2V_UNCONNECTED_718, SV2V_UNCONNECTED_719, SV2V_UNCONNECTED_720, SV2V_UNCONNECTED_721, SV2V_UNCONNECTED_722, SV2V_UNCONNECTED_723, SV2V_UNCONNECTED_724, SV2V_UNCONNECTED_725, SV2V_UNCONNECTED_726, SV2V_UNCONNECTED_727, SV2V_UNCONNECTED_728, SV2V_UNCONNECTED_729, SV2V_UNCONNECTED_730, SV2V_UNCONNECTED_731, SV2V_UNCONNECTED_732, SV2V_UNCONNECTED_733, SV2V_UNCONNECTED_734, SV2V_UNCONNECTED_735, SV2V_UNCONNECTED_736, SV2V_UNCONNECTED_737, SV2V_UNCONNECTED_738, SV2V_UNCONNECTED_739, SV2V_UNCONNECTED_740, SV2V_UNCONNECTED_741, SV2V_UNCONNECTED_742, SV2V_UNCONNECTED_743, SV2V_UNCONNECTED_744, SV2V_UNCONNECTED_745, SV2V_UNCONNECTED_746, SV2V_UNCONNECTED_747, SV2V_UNCONNECTED_748, SV2V_UNCONNECTED_749, SV2V_UNCONNECTED_750, SV2V_UNCONNECTED_751, SV2V_UNCONNECTED_752, SV2V_UNCONNECTED_753, SV2V_UNCONNECTED_754, SV2V_UNCONNECTED_755, SV2V_UNCONNECTED_756, SV2V_UNCONNECTED_757, SV2V_UNCONNECTED_758, SV2V_UNCONNECTED_759, SV2V_UNCONNECTED_760, SV2V_UNCONNECTED_761, SV2V_UNCONNECTED_762, SV2V_UNCONNECTED_763, SV2V_UNCONNECTED_764, SV2V_UNCONNECTED_765, SV2V_UNCONNECTED_766, SV2V_UNCONNECTED_767, SV2V_UNCONNECTED_768, SV2V_UNCONNECTED_769, SV2V_UNCONNECTED_770, SV2V_UNCONNECTED_771, SV2V_UNCONNECTED_772, SV2V_UNCONNECTED_773, SV2V_UNCONNECTED_774, SV2V_UNCONNECTED_775, SV2V_UNCONNECTED_776, SV2V_UNCONNECTED_777, SV2V_UNCONNECTED_778, SV2V_UNCONNECTED_779, SV2V_UNCONNECTED_780, SV2V_UNCONNECTED_781, SV2V_UNCONNECTED_782, SV2V_UNCONNECTED_783, SV2V_UNCONNECTED_784, SV2V_UNCONNECTED_785, SV2V_UNCONNECTED_786, SV2V_UNCONNECTED_787, SV2V_UNCONNECTED_788, SV2V_UNCONNECTED_789, SV2V_UNCONNECTED_790, SV2V_UNCONNECTED_791, SV2V_UNCONNECTED_792, SV2V_UNCONNECTED_793, SV2V_UNCONNECTED_794, SV2V_UNCONNECTED_795, SV2V_UNCONNECTED_796, SV2V_UNCONNECTED_797, SV2V_UNCONNECTED_798, SV2V_UNCONNECTED_799, SV2V_UNCONNECTED_800, SV2V_UNCONNECTED_801, SV2V_UNCONNECTED_802, SV2V_UNCONNECTED_803, SV2V_UNCONNECTED_804, SV2V_UNCONNECTED_805, SV2V_UNCONNECTED_806, SV2V_UNCONNECTED_807, SV2V_UNCONNECTED_808, SV2V_UNCONNECTED_809, SV2V_UNCONNECTED_810, SV2V_UNCONNECTED_811, SV2V_UNCONNECTED_812, SV2V_UNCONNECTED_813, SV2V_UNCONNECTED_814, SV2V_UNCONNECTED_815, SV2V_UNCONNECTED_816, SV2V_UNCONNECTED_817, SV2V_UNCONNECTED_818, SV2V_UNCONNECTED_819, SV2V_UNCONNECTED_820, SV2V_UNCONNECTED_821, SV2V_UNCONNECTED_822, SV2V_UNCONNECTED_823, SV2V_UNCONNECTED_824, SV2V_UNCONNECTED_825, SV2V_UNCONNECTED_826, SV2V_UNCONNECTED_827, SV2V_UNCONNECTED_828, SV2V_UNCONNECTED_829, SV2V_UNCONNECTED_830, SV2V_UNCONNECTED_831, SV2V_UNCONNECTED_832, SV2V_UNCONNECTED_833, SV2V_UNCONNECTED_834, SV2V_UNCONNECTED_835, SV2V_UNCONNECTED_836, SV2V_UNCONNECTED_837, SV2V_UNCONNECTED_838, SV2V_UNCONNECTED_839, SV2V_UNCONNECTED_840, SV2V_UNCONNECTED_841, SV2V_UNCONNECTED_842, SV2V_UNCONNECTED_843, SV2V_UNCONNECTED_844, SV2V_UNCONNECTED_845, SV2V_UNCONNECTED_846, SV2V_UNCONNECTED_847, SV2V_UNCONNECTED_848, SV2V_UNCONNECTED_849, SV2V_UNCONNECTED_850, SV2V_UNCONNECTED_851, SV2V_UNCONNECTED_852, SV2V_UNCONNECTED_853, SV2V_UNCONNECTED_854, SV2V_UNCONNECTED_855, SV2V_UNCONNECTED_856, SV2V_UNCONNECTED_857, SV2V_UNCONNECTED_858, SV2V_UNCONNECTED_859, SV2V_UNCONNECTED_860, SV2V_UNCONNECTED_861, SV2V_UNCONNECTED_862, SV2V_UNCONNECTED_863, SV2V_UNCONNECTED_864, SV2V_UNCONNECTED_865, SV2V_UNCONNECTED_866, SV2V_UNCONNECTED_867, SV2V_UNCONNECTED_868, SV2V_UNCONNECTED_869, SV2V_UNCONNECTED_870, SV2V_UNCONNECTED_871, SV2V_UNCONNECTED_872, SV2V_UNCONNECTED_873, SV2V_UNCONNECTED_874, SV2V_UNCONNECTED_875, SV2V_UNCONNECTED_876, SV2V_UNCONNECTED_877, SV2V_UNCONNECTED_878, SV2V_UNCONNECTED_879, SV2V_UNCONNECTED_880, SV2V_UNCONNECTED_881, SV2V_UNCONNECTED_882, SV2V_UNCONNECTED_883, SV2V_UNCONNECTED_884, SV2V_UNCONNECTED_885, SV2V_UNCONNECTED_886, SV2V_UNCONNECTED_887, SV2V_UNCONNECTED_888, SV2V_UNCONNECTED_889, SV2V_UNCONNECTED_890, SV2V_UNCONNECTED_891, SV2V_UNCONNECTED_892, SV2V_UNCONNECTED_893, SV2V_UNCONNECTED_894, SV2V_UNCONNECTED_895, SV2V_UNCONNECTED_896, SV2V_UNCONNECTED_897, SV2V_UNCONNECTED_898, SV2V_UNCONNECTED_899, SV2V_UNCONNECTED_900, SV2V_UNCONNECTED_901, SV2V_UNCONNECTED_902, SV2V_UNCONNECTED_903, SV2V_UNCONNECTED_904, SV2V_UNCONNECTED_905, SV2V_UNCONNECTED_906, SV2V_UNCONNECTED_907, SV2V_UNCONNECTED_908, SV2V_UNCONNECTED_909, T9[0:0], T12, T13 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> T15;
  assign N335 = N368 | N351;
  assign N336 = N385 | N400;
  assign N337 = notSigSum[32] | notSigSum[33];
  assign N338 = notSigSum[31] | N337;
  assign N339 = notSigSum[30] | N338;
  assign N340 = notSigSum[29] | N339;
  assign N341 = notSigSum[28] | N340;
  assign N342 = notSigSum[27] | N341;
  assign N343 = notSigSum[26] | N342;
  assign N344 = notSigSum[25] | N343;
  assign N345 = notSigSum[24] | N344;
  assign N346 = notSigSum[23] | N345;
  assign N347 = notSigSum[22] | N346;
  assign N348 = notSigSum[21] | N347;
  assign N349 = notSigSum[20] | N348;
  assign N350 = notSigSum[19] | N349;
  assign N351 = notSigSum[18] | N350;
  assign N352 = T141[16] | T141[17];
  assign N353 = T141[15] | N352;
  assign N354 = T141[14] | N353;
  assign N355 = T141[13] | N354;
  assign N356 = T141[12] | N355;
  assign N357 = T141[11] | N356;
  assign N358 = T141[10] | N357;
  assign N359 = T141[9] | N358;
  assign N360 = T141[8] | N359;
  assign N361 = T141[7] | N360;
  assign N362 = T141[6] | N361;
  assign N363 = T141[5] | N362;
  assign N364 = T141[4] | N363;
  assign N365 = T141[3] | N364;
  assign N366 = T141[2] | N365;
  assign N367 = T141[1] | N366;
  assign N368 = T141[0] | N367;
  assign N369 = io_mulAddResult[15] | io_mulAddResult[16];
  assign N370 = io_mulAddResult[14] | N369;
  assign N371 = io_mulAddResult[13] | N370;
  assign N372 = io_mulAddResult[12] | N371;
  assign N373 = io_mulAddResult[11] | N372;
  assign N374 = io_mulAddResult[10] | N373;
  assign N375 = io_mulAddResult[9] | N374;
  assign N376 = io_mulAddResult[8] | N375;
  assign N377 = io_mulAddResult[7] | N376;
  assign N378 = io_mulAddResult[6] | N377;
  assign N379 = io_mulAddResult[5] | N378;
  assign N380 = io_mulAddResult[4] | N379;
  assign N381 = io_mulAddResult[3] | N380;
  assign N382 = io_mulAddResult[2] | N381;
  assign N383 = io_mulAddResult[1] | N382;
  assign N384 = io_mulAddResult[0] | N383;
  assign N385 = io_fromPreMul_bit0AlignedNegSigC | N384;
  assign N386 = io_mulAddResult[31] | io_mulAddResult[32];
  assign N387 = io_mulAddResult[30] | N386;
  assign N388 = io_mulAddResult[29] | N387;
  assign N389 = io_mulAddResult[28] | N388;
  assign N390 = io_mulAddResult[27] | N389;
  assign N391 = io_mulAddResult[26] | N390;
  assign N392 = io_mulAddResult[25] | N391;
  assign N393 = io_mulAddResult[24] | N392;
  assign N394 = io_mulAddResult[23] | N393;
  assign N395 = io_mulAddResult[22] | N394;
  assign N396 = io_mulAddResult[21] | N395;
  assign N397 = io_mulAddResult[20] | N396;
  assign N398 = io_mulAddResult[19] | N397;
  assign N399 = io_mulAddResult[18] | N398;
  assign N400 = io_mulAddResult[17] | N399;
  assign T27 = io_fromPreMul_highAlignedNegSigC + 1'b1;
  assign T475 = io_fromPreMul_CAlignDist[4:0] - 1'b1;
  assign { T128[31:31], T128_0 } = 1'b0 - T488[0];
  assign { T148[15:15], T148_0 } = 1'b0 - T488[0];
  assign T16 = { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } - T376;
  assign { sExpX3[10:10], sExpX3_13 } = io_fromPreMul_sExpSum - T375;
  assign T234 = sExpX3_13 - 1'b1;
  assign T284 = sExpX3_13 + 1'b1;
  assign { T77[26:26], T77_0 } = 1'b0 - sExpX3[10];
  assign roundUp_sigY3 = T242 + 1'b1;
  assign { T313[22:22], T313_0 } = 1'b0 - T504[0];
  assign inexactY = (N0)? T215 : 
                    (N1)? anyRound : 1'b0;
  assign N0 = doIncrSig;
  assign N1 = N132;
  assign T375 = (N2)? CDom_estNormDist : 
                (N3)? T16 : 1'b0;
  assign N2 = io_fromPreMul_isCDominant;
  assign N3 = N192;
  assign T376 = (N4)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N5)? T378 : 1'b0;
  assign N4 = T18[49];
  assign N5 = N133;
  assign T378 = (N6)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N7)? T379 : 1'b0;
  assign N6 = T18[48];
  assign N7 = N134;
  assign T379 = (N8)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N9)? T380 : 1'b0;
  assign N8 = T18[47];
  assign N9 = N135;
  assign T380 = (N10)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N11)? T381 : 1'b0;
  assign N10 = T18[46];
  assign N11 = N136;
  assign T381 = (N12)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N13)? T382 : 1'b0;
  assign N12 = T18[45];
  assign N13 = N137;
  assign T382 = (N14)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N15)? T383 : 1'b0;
  assign N14 = T18[44];
  assign N15 = N138;
  assign T383 = (N16)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N17)? T384 : 1'b0;
  assign N16 = T18[43];
  assign N17 = N139;
  assign T384 = (N18)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N19)? T385 : 1'b0;
  assign N18 = T18[42];
  assign N19 = N140;
  assign T385 = (N20)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N21)? T386 : 1'b0;
  assign N20 = T18[41];
  assign N21 = N141;
  assign T386 = (N22)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N23)? T387 : 1'b0;
  assign N22 = T18[40];
  assign N23 = N142;
  assign T387 = (N24)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N25)? T388 : 1'b0;
  assign N24 = T18[39];
  assign N25 = N143;
  assign T388 = (N26)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N27)? T389 : 1'b0;
  assign N26 = T18[38];
  assign N27 = N144;
  assign T389 = (N28)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N29)? T390 : 1'b0;
  assign N28 = T18[37];
  assign N29 = N145;
  assign T390 = (N30)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N31)? T391 : 1'b0;
  assign N30 = T18[36];
  assign N31 = N146;
  assign T391 = (N32)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N33)? T392 : 1'b0;
  assign N32 = T18[35];
  assign N33 = N147;
  assign T392 = (N34)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N35)? T393 : 1'b0;
  assign N34 = T18[34];
  assign N35 = N148;
  assign T393 = (N36)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N37)? T394 : 1'b0;
  assign N36 = T18[33];
  assign N37 = N149;
  assign T394[4:0] = (N38)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N39)? T395 : 1'b0;
  assign N38 = T394[5];
  assign N39 = N150;
  assign T395 = (N40)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N41)? T396 : 1'b0;
  assign N40 = T18[31];
  assign N41 = N151;
  assign T396 = (N42)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N43)? T397 : 1'b0;
  assign N42 = T18[30];
  assign N43 = N152;
  assign T397 = (N44)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N45)? T398 : 1'b0;
  assign N44 = T18[29];
  assign N45 = N153;
  assign T398 = (N46)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N47)? T399 : 1'b0;
  assign N46 = T18[28];
  assign N47 = N154;
  assign T399 = (N48)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N49)? T400 : 1'b0;
  assign N48 = T18[27];
  assign N49 = N155;
  assign T400 = (N50)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N51)? T401 : 1'b0;
  assign N50 = T18[26];
  assign N51 = N156;
  assign T401 = (N52)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N53)? T402 : 1'b0;
  assign N52 = T18[25];
  assign N53 = N157;
  assign T402 = (N54)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N55)? T403 : 1'b0;
  assign N54 = T18[24];
  assign N55 = N158;
  assign T403 = (N56)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N57)? T404 : 1'b0;
  assign N56 = T18[23];
  assign N57 = N159;
  assign T404 = (N58)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N59)? T405 : 1'b0;
  assign N58 = T18[22];
  assign N59 = N160;
  assign T405 = (N60)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N61)? T406 : 1'b0;
  assign N60 = T18[21];
  assign N61 = N161;
  assign T406 = (N62)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N63)? T407 : 1'b0;
  assign N62 = T18[20];
  assign N63 = N162;
  assign T407 = (N64)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N65)? T408 : 1'b0;
  assign N64 = T18[19];
  assign N65 = N163;
  assign T408 = (N66)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N67)? T409 : 1'b0;
  assign N66 = T18[18];
  assign N67 = N164;
  assign T409 = (N68)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N69)? T410 : 1'b0;
  assign N68 = T18[17];
  assign N69 = N165;
  assign T410[3:0] = (N70)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N71)? T411 : 1'b0;
  assign N70 = T410[4];
  assign N71 = N166;
  assign T411 = (N72)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N73)? T412 : 1'b0;
  assign N72 = T18[15];
  assign N73 = N167;
  assign T412 = (N74)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N75)? T413 : 1'b0;
  assign N74 = T18[14];
  assign N75 = N168;
  assign T413 = (N76)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N77)? T414 : 1'b0;
  assign N76 = T18[13];
  assign N77 = N169;
  assign T414 = (N78)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N79)? T415 : 1'b0;
  assign N78 = T18[12];
  assign N79 = N170;
  assign T415 = (N80)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N81)? T416 : 1'b0;
  assign N80 = T18[11];
  assign N81 = N171;
  assign T416 = (N82)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N83)? T417 : 1'b0;
  assign N82 = T18[10];
  assign N83 = N172;
  assign T417 = (N84)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N85)? T418 : 1'b0;
  assign N84 = T18[9];
  assign N85 = N173;
  assign T418[2:0] = (N86)? { 1'b0, 1'b0, 1'b0 } : 
                     (N87)? T419 : 1'b0;
  assign N86 = T418[3];
  assign N87 = N174;
  assign T419 = (N88)? { 1'b1, 1'b1, 1'b1 } : 
                (N89)? T420 : 1'b0;
  assign N88 = T18[7];
  assign N89 = N175;
  assign T420 = (N90)? { 1'b1, 1'b1, 1'b0 } : 
                (N91)? T421 : 1'b0;
  assign N90 = T18[6];
  assign N91 = N176;
  assign T421 = (N92)? { 1'b1, 1'b0, 1'b1 } : 
                (N93)? T422 : 1'b0;
  assign N92 = T18[5];
  assign N93 = N177;
  assign T422[1:0] = (N94)? { 1'b0, 1'b0 } : 
                     (N95)? T423 : 1'b0;
  assign N94 = T422[2];
  assign N95 = N178;
  assign T423 = (N96)? { 1'b1, 1'b1 } : 
                (N97)? T424 : 1'b0;
  assign N96 = T18[3];
  assign N97 = N179;
  assign T424[0] = (N98)? 1'b0 : 
                   (N99)? T18[1] : 1'b0;
  assign N98 = T424[1];
  assign N99 = N180;
  assign { sigSum, T21 } = (N100)? T27 : 
                           (N101)? io_fromPreMul_highAlignedNegSigC : 1'b0;
  assign N100 = io_mulAddResult[48];
  assign N101 = N181;
  assign CDom_estNormDist = (N102)? io_fromPreMul_CAlignDist : 
                            (N103)? { 1'b0, 1'b0, T475 } : 1'b0;
  assign N102 = T32;
  assign N103 = N182;
  assign sigX3[0] = (N0)? N313 : 
                    (N1)? N328 : 1'b0;
  assign { cFirstNormAbsSigSum, T125 } = (N104)? T192 : 
                                         (N105)? { 1'b0, T487 } : 1'b0;
  assign N104 = sigSum[51];
  assign N105 = N183;
  assign T487 = (N2)? CDom_firstNormAbsSigSum : 
                (N3)? notCDom_pos_firstNormAbsSigSum : 1'b0;
  assign notCDom_pos_firstNormAbsSigSum = (N106)? T146 : 
                                          (N107)? T127 : 1'b0;
  assign N106 = T16[5];
  assign N107 = N184;
  assign T127 = (N108)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T21, io_mulAddResult[47:17], T489[0:0] } : 
                (N109)? { io_mulAddResult[9:0], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128[31:31], T128_0 } : 1'b0;
  assign N108 = T16[4];
  assign N109 = N185;
  assign T489[0] = (N110)? T138 : 
                   (N111)? N385 : 1'b0;
  assign N110 = T488[0];
  assign N111 = N186;
  assign T146 = (N108)? { io_mulAddResult[25:0], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148[15:15], T148_0 } : 
                (N109)? io_mulAddResult[41:0] : 1'b0;
  assign T192 = (N2)? { 1'b0, CDom_firstNormAbsSigSum } : 
                (N3)? notCDom_neg_cFirstNormAbsSigSum : 1'b0;
  assign notCDom_neg_cFirstNormAbsSigSum = (N106)? T200 : 
                                           (N107)? T193 : 1'b0;
  assign T193 = (N108)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, notSigSum[49:18], N368 } : 
                (N109)? { T141[11:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T200 = (N108)? { notSigSum[27:18], T141[17:1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N109)? { 1'b0, notSigSum[42:18], T141[17:1] } : 1'b0;
  assign T233 = (N112)? T234 : 
                (N113)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N112 = N212;
  assign N113 = N211;
  assign T237 = (N114)? T238 : 
                (N115)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N114 = roundEven;
  assign N115 = N188;
  assign roundEven = (N0)? T247 : 
                     (N1)? T244 : 1'b0;
  assign T251 = (N116)? roundUp_sigY3 : 
                (N117)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N116 = T252;
  assign N117 = N189;
  assign roundDirectUp = (N118)? N331 : 
                         (N119)? N297 : 1'b0;
  assign N118 = signY;
  assign N119 = N190;
  assign signY = (N120)? N331 : 
                 (N121)? T255 : 1'b0;
  assign N120 = isZeroY;
  assign N121 = N191;
  assign doNegSignSum = (N2)? T256 : 
                        (N3)? sigSum[51] : 1'b0;
  assign T272 = (N122)? T273 : 
                (N123)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N122 = T276;
  assign N123 = N193;
  assign T281 = (N124)? sExpX3_13 : 
                (N125)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N124 = T236[0];
  assign N125 = N194;
  assign T283 = (N126)? T284 : 
                (N127)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N126 = T236[1];
  assign N127 = N195;
  assign T322 = (N128)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N129)? fractY : 1'b0;
  assign N128 = T325;
  assign N129 = N196;
  assign fractY = (N130)? sigY3[22:0] : 
                  (N131)? sigY3[23:1] : 1'b0;
  assign N130 = sigX3Shift1;
  assign N131 = N187;
  assign io_exceptionFlags[0] = io_exceptionFlags[2] | T3;
  assign T3 = commonCase & inexactY;
  assign N132 = ~doIncrSig;
  assign anyRound = N267 | N294;
  assign T4[27] = sigX3_27 & 1'b0;
  assign T4[26] = T374[0] & 1'b0;
  assign T4[25] = sigX3[25] & T373[25];
  assign T4[24] = sigX3[24] & T373[24];
  assign T4[23] = sigX3[23] & T373[23];
  assign T4[22] = sigX3[22] & T373[22];
  assign T4[21] = sigX3[21] & T373[21];
  assign T4[20] = sigX3[20] & T373[20];
  assign T4[19] = sigX3[19] & T373[19];
  assign T4[18] = sigX3[18] & T373[18];
  assign T4[17] = sigX3[17] & T373[17];
  assign T4[16] = sigX3[16] & T373[16];
  assign T4[15] = sigX3[15] & T373[15];
  assign T4[14] = sigX3[14] & T373[14];
  assign T4[13] = sigX3[13] & T373[13];
  assign T4[12] = sigX3[12] & T373[12];
  assign T4[11] = sigX3[11] & T373[11];
  assign T4[10] = sigX3[10] & T373[10];
  assign T4[9] = sigX3[9] & T373[9];
  assign T4[8] = sigX3[8] & T373[8];
  assign T4[7] = sigX3[7] & T373[7];
  assign T4[6] = sigX3[6] & T373[6];
  assign T4[5] = sigX3[5] & T373[5];
  assign T4[4] = sigX3[4] & T373[4];
  assign T4[3] = sigX3[3] & T373[3];
  assign T4[2] = sigX3[2] & T373[2];
  assign T4[1] = sigX3[1] & T373[1];
  assign T4[0] = sigX3[0] & T373[0];
  assign T373[25] = T77[26] | T6[26];
  assign T373[24] = T77[26] | T6[25];
  assign T373[23] = T77[26] | T6[24];
  assign T373[22] = T77[26] | T6[23];
  assign T373[21] = T77[26] | T6[22];
  assign T373[20] = T77[26] | T6[21];
  assign T373[19] = T77[26] | T6[20];
  assign T373[18] = T77[26] | T6[19];
  assign T373[17] = T77[26] | T6[18];
  assign T373[16] = T77[26] | T6[17];
  assign T373[15] = T77[26] | T6[16];
  assign T373[14] = T77[26] | T6[15];
  assign T373[13] = T77[26] | T6[14];
  assign T373[12] = T77[26] | T6[13];
  assign T373[11] = T77[26] | T6[12];
  assign T373[10] = T77[26] | T6[11];
  assign T373[9] = T77[26] | T6[10];
  assign T373[8] = T77[26] | T6[9];
  assign T373[7] = T77[26] | T6[8];
  assign T373[6] = T77[26] | T6[7];
  assign T373[5] = T77[26] | T6[6];
  assign T373[4] = T77[26] | T6[5];
  assign T373[3] = T77[26] | T6[4];
  assign T373[2] = T77[26] | T6[3];
  assign T373[1] = T77[26] | T6[2];
  assign T373[0] = T77[26] | 1'b1;
  assign roundMask[0] = T77_0 | 1'b1;
  assign T6[26] = T9[24] | 1'b0;
  assign T6[25] = T9[23] | 1'b0;
  assign T6[24] = T9[22] | 1'b0;
  assign T6[23] = T9[21] | 1'b0;
  assign T6[22] = T9[20] | 1'b0;
  assign T6[21] = T9[19] | 1'b0;
  assign T6[20] = T9[18] | 1'b0;
  assign T6[19] = T9[17] | 1'b0;
  assign T6[18] = T9[16] | 1'b0;
  assign T6[17] = T9[15] | 1'b0;
  assign T6[16] = T9[14] | 1'b0;
  assign T6[15] = T9[13] | 1'b0;
  assign T6[14] = T9[12] | 1'b0;
  assign T6[13] = T9[11] | 1'b0;
  assign T6[12] = T9[10] | 1'b0;
  assign T6[11] = T9[9] | 1'b0;
  assign T6[10] = T9[8] | 1'b0;
  assign T6[9] = T9[7] | 1'b0;
  assign T6[8] = T9[6] | 1'b0;
  assign T6[7] = T9[5] | 1'b0;
  assign T6[6] = T9[4] | 1'b0;
  assign T6[5] = T9[3] | 1'b0;
  assign T6[4] = T9[2] | 1'b0;
  assign T6[3] = T9[1] | 1'b0;
  assign T6[2] = T9[0] | T374[0];
  assign T15[9] = ~sExpX3_13[9];
  assign T15[8] = ~sExpX3_13[8];
  assign T15[7] = ~sExpX3_13[7];
  assign T15[6] = ~sExpX3_13[6];
  assign T15[5] = ~sExpX3_13[5];
  assign T15[4] = ~sExpX3_13[4];
  assign T15[3] = ~sExpX3_13[3];
  assign T15[2] = ~sExpX3_13[2];
  assign T15[1] = ~sExpX3_13[1];
  assign T15[0] = ~sExpX3_13[0];
  assign N133 = ~T18[49];
  assign N134 = ~T18[48];
  assign N135 = ~T18[47];
  assign N136 = ~T18[46];
  assign N137 = ~T18[45];
  assign N138 = ~T18[44];
  assign N139 = ~T18[43];
  assign N140 = ~T18[42];
  assign N141 = ~T18[41];
  assign N142 = ~T18[40];
  assign N143 = ~T18[39];
  assign N144 = ~T18[38];
  assign N145 = ~T18[37];
  assign N146 = ~T18[36];
  assign N147 = ~T18[35];
  assign N148 = ~T18[34];
  assign N149 = ~T18[33];
  assign N150 = ~T18[32];
  assign T394[5] = T18[32];
  assign N151 = ~T18[31];
  assign N152 = ~T18[30];
  assign N153 = ~T18[29];
  assign N154 = ~T18[28];
  assign N155 = ~T18[27];
  assign N156 = ~T18[26];
  assign N157 = ~T18[25];
  assign N158 = ~T18[24];
  assign N159 = ~T18[23];
  assign N160 = ~T18[22];
  assign N161 = ~T18[21];
  assign N162 = ~T18[20];
  assign N163 = ~T18[19];
  assign N164 = ~T18[18];
  assign N165 = ~T18[17];
  assign N166 = ~T18[16];
  assign T410[4] = T18[16];
  assign N167 = ~T18[15];
  assign N168 = ~T18[14];
  assign N169 = ~T18[13];
  assign N170 = ~T18[12];
  assign N171 = ~T18[11];
  assign N172 = ~T18[10];
  assign N173 = ~T18[9];
  assign N174 = ~T18[8];
  assign T418[3] = T18[8];
  assign N175 = ~T18[7];
  assign N176 = ~T18[6];
  assign N177 = ~T18[5];
  assign N178 = ~T18[4];
  assign T422[2] = T18[4];
  assign N179 = ~T18[3];
  assign N180 = ~T18[2];
  assign T424[1] = T18[2];
  assign T18[49] = T21[50] ^ T21[49];
  assign T18[48] = T21[49] ^ io_mulAddResult[47];
  assign T18[47] = io_mulAddResult[47] ^ io_mulAddResult[46];
  assign T18[46] = io_mulAddResult[46] ^ io_mulAddResult[45];
  assign T18[45] = io_mulAddResult[45] ^ io_mulAddResult[44];
  assign T18[44] = io_mulAddResult[44] ^ io_mulAddResult[43];
  assign T18[43] = io_mulAddResult[43] ^ io_mulAddResult[42];
  assign T18[42] = io_mulAddResult[42] ^ io_mulAddResult[41];
  assign T18[41] = io_mulAddResult[41] ^ io_mulAddResult[40];
  assign T18[40] = io_mulAddResult[40] ^ io_mulAddResult[39];
  assign T18[39] = io_mulAddResult[39] ^ io_mulAddResult[38];
  assign T18[38] = io_mulAddResult[38] ^ io_mulAddResult[37];
  assign T18[37] = io_mulAddResult[37] ^ io_mulAddResult[36];
  assign T18[36] = io_mulAddResult[36] ^ io_mulAddResult[35];
  assign T18[35] = io_mulAddResult[35] ^ io_mulAddResult[34];
  assign T18[34] = io_mulAddResult[34] ^ io_mulAddResult[33];
  assign T18[33] = io_mulAddResult[33] ^ io_mulAddResult[32];
  assign T18[32] = io_mulAddResult[32] ^ io_mulAddResult[31];
  assign T18[31] = io_mulAddResult[31] ^ io_mulAddResult[30];
  assign T18[30] = io_mulAddResult[30] ^ io_mulAddResult[29];
  assign T18[29] = io_mulAddResult[29] ^ io_mulAddResult[28];
  assign T18[28] = io_mulAddResult[28] ^ io_mulAddResult[27];
  assign T18[27] = io_mulAddResult[27] ^ io_mulAddResult[26];
  assign T18[26] = io_mulAddResult[26] ^ io_mulAddResult[25];
  assign T18[25] = io_mulAddResult[25] ^ io_mulAddResult[24];
  assign T18[24] = io_mulAddResult[24] ^ io_mulAddResult[23];
  assign T18[23] = io_mulAddResult[23] ^ io_mulAddResult[22];
  assign T18[22] = io_mulAddResult[22] ^ io_mulAddResult[21];
  assign T18[21] = io_mulAddResult[21] ^ io_mulAddResult[20];
  assign T18[20] = io_mulAddResult[20] ^ io_mulAddResult[19];
  assign T18[19] = io_mulAddResult[19] ^ io_mulAddResult[18];
  assign T18[18] = io_mulAddResult[18] ^ io_mulAddResult[17];
  assign T18[17] = io_mulAddResult[17] ^ io_mulAddResult[16];
  assign T18[16] = io_mulAddResult[16] ^ io_mulAddResult[15];
  assign T18[15] = io_mulAddResult[15] ^ io_mulAddResult[14];
  assign T18[14] = io_mulAddResult[14] ^ io_mulAddResult[13];
  assign T18[13] = io_mulAddResult[13] ^ io_mulAddResult[12];
  assign T18[12] = io_mulAddResult[12] ^ io_mulAddResult[11];
  assign T18[11] = io_mulAddResult[11] ^ io_mulAddResult[10];
  assign T18[10] = io_mulAddResult[10] ^ io_mulAddResult[9];
  assign T18[9] = io_mulAddResult[9] ^ io_mulAddResult[8];
  assign T18[8] = io_mulAddResult[8] ^ io_mulAddResult[7];
  assign T18[7] = io_mulAddResult[7] ^ io_mulAddResult[6];
  assign T18[6] = io_mulAddResult[6] ^ io_mulAddResult[5];
  assign T18[5] = io_mulAddResult[5] ^ io_mulAddResult[4];
  assign T18[4] = io_mulAddResult[4] ^ io_mulAddResult[3];
  assign T18[3] = io_mulAddResult[3] ^ io_mulAddResult[2];
  assign T18[2] = io_mulAddResult[2] ^ io_mulAddResult[1];
  assign T18[1] = io_mulAddResult[1] ^ io_mulAddResult[0];
  assign N181 = ~io_mulAddResult[48];
  assign N182 = ~T32;
  assign T32 = io_fromPreMul_CAlignDist_0 | T488[0];
  assign T488[0] = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T9[8] = 1'b0 | T34[7];
  assign T9[7] = T37[7] | 1'b0;
  assign T9[6] = 1'b0 | T34_5;
  assign T9[5] = T35[6] | 1'b0;
  assign T9[4] = 1'b0 | T34_3;
  assign T9[3] = T35_4 | 1'b0;
  assign T9[2] = 1'b0 | T34_1;
  assign T9[1] = T35_2 | 1'b0;
  assign T37[7] = 1'b0 | T38[7];
  assign T34[7] = 1'b0 | T38[6];
  assign T35[6] = T41[7] | 1'b0;
  assign T34_5 = T41[6] | 1'b0;
  assign T35_4 = 1'b0 | T38_3;
  assign T34_3 = 1'b0 | T38_2;
  assign T35_2 = T39[5] | 1'b0;
  assign T34_1 = T39[4] | 1'b0;
  assign T41[7] = 1'b0 | T12[3];
  assign T41[6] = 1'b0 | T12[2];
  assign T38[7] = 1'b0 | T12[1];
  assign T38[6] = 1'b0 | T12[0];
  assign T39[5] = T12[7] | 1'b0;
  assign T39[4] = T12[6] | 1'b0;
  assign T38_3 = T12[5] | 1'b0;
  assign T38_2 = T12[4] | 1'b0;
  assign T9[24] = 1'b0 | T53[15];
  assign T9[23] = T56[15] | 1'b0;
  assign T9[22] = 1'b0 | T53_13;
  assign T9[21] = T54[14] | 1'b0;
  assign T9[20] = 1'b0 | T53_11;
  assign T9[19] = T54_12 | 1'b0;
  assign T9[18] = 1'b0 | T53_9;
  assign T9[17] = T54_10 | 1'b0;
  assign T9[16] = 1'b0 | T53_7;
  assign T9[15] = T54_8 | 1'b0;
  assign T9[14] = 1'b0 | T53_5;
  assign T9[13] = T54_6 | 1'b0;
  assign T9[12] = 1'b0 | T53_3;
  assign T9[11] = T54_4 | 1'b0;
  assign T9[10] = 1'b0 | T53_1;
  assign T9[9] = T54_2 | 1'b0;
  assign T56[15] = 1'b0 | T57[15];
  assign T53[15] = 1'b0 | T57[14];
  assign T54[14] = T60[15] | 1'b0;
  assign T53_13 = T60[14] | 1'b0;
  assign T54_12 = 1'b0 | T57_11;
  assign T53_11 = 1'b0 | T57_10;
  assign T54_10 = T58[13] | 1'b0;
  assign T53_9 = T58[12] | 1'b0;
  assign T54_8 = 1'b0 | T57_7;
  assign T53_7 = 1'b0 | T57_6;
  assign T54_6 = T58_9 | 1'b0;
  assign T53_5 = T58_8 | 1'b0;
  assign T54_4 = 1'b0 | T57_3;
  assign T53_3 = 1'b0 | T57_2;
  assign T54_2 = T58_5 | 1'b0;
  assign T53_1 = T58_4 | 1'b0;
  assign T60[15] = 1'b0 | T61[15];
  assign T60[14] = 1'b0 | T61[14];
  assign T57[15] = 1'b0 | T61[13];
  assign T57[14] = 1'b0 | T61[12];
  assign T58[13] = T64[15] | 1'b0;
  assign T58[12] = T64[14] | 1'b0;
  assign T57_11 = T64[13] | 1'b0;
  assign T57_10 = T64[12] | 1'b0;
  assign T58_9 = 1'b0 | T61_7;
  assign T58_8 = 1'b0 | T61_6;
  assign T57_7 = 1'b0 | T61_5;
  assign T57_6 = 1'b0 | T61_4;
  assign T58_5 = T62[11] | 1'b0;
  assign T58_4 = T62[10] | 1'b0;
  assign T57_3 = T62[9] | 1'b0;
  assign T57_2 = T62[8] | 1'b0;
  assign T64[15] = 1'b0 | T13[7];
  assign T64[14] = 1'b0 | T13[6];
  assign T64[13] = 1'b0 | T13[5];
  assign T64[12] = 1'b0 | T13[4];
  assign T61[15] = 1'b0 | T13[3];
  assign T61[14] = 1'b0 | T13[2];
  assign T61[13] = 1'b0 | T13[1];
  assign T61[12] = 1'b0 | T13[0];
  assign T62[11] = T13[15] | 1'b0;
  assign T62[10] = T13[14] | 1'b0;
  assign T62[9] = T13[13] | 1'b0;
  assign T62[8] = T13[12] | 1'b0;
  assign T61_7 = T13[11] | 1'b0;
  assign T61_6 = T13[10] | 1'b0;
  assign T61_5 = T13[9] | 1'b0;
  assign T61_4 = T13[8] | 1'b0;
  assign T82[15] = T125[15] & absSigSumExtraMask[15];
  assign T82[14] = T125[14] & absSigSumExtraMask[14];
  assign T82[13] = T125[13] & absSigSumExtraMask[13];
  assign T82[12] = T125[12] & absSigSumExtraMask[12];
  assign T82[11] = T125[11] & absSigSumExtraMask[11];
  assign T82[10] = T125[10] & absSigSumExtraMask[10];
  assign T82[9] = T125[9] & absSigSumExtraMask[9];
  assign T82[8] = T125[8] & absSigSumExtraMask[8];
  assign T82[7] = T125[7] & T88[0];
  assign T82[6] = T125[6] & T88[1];
  assign T82[5] = T125[5] & T88[2];
  assign T82[4] = T125[4] & T88[3];
  assign T82[3] = T125[3] & T87[0];
  assign T82[2] = T125[2] & T87[1];
  assign T82[1] = T125[1] & absSigSumExtraMask_1;
  assign T82[0] = T125[0] & 1'b1;
  assign normTo2ShiftDist[3] = ~T375[3];
  assign normTo2ShiftDist[2] = ~T375[2];
  assign normTo2ShiftDist[1] = ~T375[1];
  assign normTo2ShiftDist[0] = ~T375[0];
  assign absSigSumExtraMask[15] = 1'b0 | T107[7];
  assign absSigSumExtraMask[14] = T110[7] | 1'b0;
  assign absSigSumExtraMask[13] = 1'b0 | T107_5;
  assign absSigSumExtraMask[12] = T108[6] | 1'b0;
  assign absSigSumExtraMask[11] = 1'b0 | T107_3;
  assign absSigSumExtraMask[10] = T108_4 | 1'b0;
  assign absSigSumExtraMask[9] = 1'b0 | T107_1;
  assign absSigSumExtraMask[8] = T108_2 | 1'b0;
  assign T110[7] = 1'b0 | T111[7];
  assign T107[7] = 1'b0 | T111[6];
  assign T108[6] = T114[7] | 1'b0;
  assign T107_5 = T114[6] | 1'b0;
  assign T108_4 = 1'b0 | T111_3;
  assign T107_3 = 1'b0 | T111_2;
  assign T108_2 = T112[5] | 1'b0;
  assign T107_1 = T112[4] | 1'b0;
  assign T114[7] = 1'b0 | T89[3];
  assign T114[6] = 1'b0 | T89[2];
  assign T111[7] = 1'b0 | T89[1];
  assign T111[6] = 1'b0 | T89[0];
  assign T112[5] = T89[7] | 1'b0;
  assign T112[4] = T89[6] | 1'b0;
  assign T111_3 = T89[5] | 1'b0;
  assign T111_2 = T89[4] | 1'b0;
  assign N183 = ~sigSum[51];
  assign N184 = ~T16[5];
  assign N185 = ~T16[4];
  assign N186 = ~T488[0];
  assign T138 = ~N368;
  assign notSigSum[74] = ~sigSum[74];
  assign notSigSum[73] = ~sigSum[73];
  assign notSigSum[72] = ~sigSum[72];
  assign notSigSum[71] = ~sigSum[71];
  assign notSigSum[70] = ~sigSum[70];
  assign notSigSum[69] = ~sigSum[69];
  assign notSigSum[68] = ~sigSum[68];
  assign notSigSum[67] = ~sigSum[67];
  assign notSigSum[66] = ~sigSum[66];
  assign notSigSum[65] = ~sigSum[65];
  assign notSigSum[64] = ~sigSum[64];
  assign notSigSum[63] = ~sigSum[63];
  assign notSigSum[62] = ~sigSum[62];
  assign notSigSum[61] = ~sigSum[61];
  assign notSigSum[60] = ~sigSum[60];
  assign notSigSum[59] = ~sigSum[59];
  assign notSigSum[58] = ~sigSum[58];
  assign notSigSum[57] = ~sigSum[57];
  assign notSigSum[56] = ~sigSum[56];
  assign notSigSum[55] = ~sigSum[55];
  assign notSigSum[54] = ~sigSum[54];
  assign notSigSum[53] = ~sigSum[53];
  assign notSigSum[52] = ~sigSum[52];
  assign notSigSum[51] = ~sigSum[51];
  assign notSigSum[50] = ~T21[50];
  assign notSigSum[49] = ~T21[49];
  assign notSigSum[48] = ~io_mulAddResult[47];
  assign notSigSum[47] = ~io_mulAddResult[46];
  assign notSigSum[46] = ~io_mulAddResult[45];
  assign notSigSum[45] = ~io_mulAddResult[44];
  assign notSigSum[44] = ~io_mulAddResult[43];
  assign notSigSum[43] = ~io_mulAddResult[42];
  assign notSigSum[42] = ~io_mulAddResult[41];
  assign notSigSum[41] = ~io_mulAddResult[40];
  assign notSigSum[40] = ~io_mulAddResult[39];
  assign notSigSum[39] = ~io_mulAddResult[38];
  assign notSigSum[38] = ~io_mulAddResult[37];
  assign notSigSum[37] = ~io_mulAddResult[36];
  assign notSigSum[36] = ~io_mulAddResult[35];
  assign notSigSum[35] = ~io_mulAddResult[34];
  assign notSigSum[34] = ~io_mulAddResult[33];
  assign notSigSum[33] = ~io_mulAddResult[32];
  assign notSigSum[32] = ~io_mulAddResult[31];
  assign notSigSum[31] = ~io_mulAddResult[30];
  assign notSigSum[30] = ~io_mulAddResult[29];
  assign notSigSum[29] = ~io_mulAddResult[28];
  assign notSigSum[28] = ~io_mulAddResult[27];
  assign notSigSum[27] = ~io_mulAddResult[26];
  assign notSigSum[26] = ~io_mulAddResult[25];
  assign notSigSum[25] = ~io_mulAddResult[24];
  assign notSigSum[24] = ~io_mulAddResult[23];
  assign notSigSum[23] = ~io_mulAddResult[22];
  assign notSigSum[22] = ~io_mulAddResult[21];
  assign notSigSum[21] = ~io_mulAddResult[20];
  assign notSigSum[20] = ~io_mulAddResult[19];
  assign notSigSum[19] = ~io_mulAddResult[18];
  assign notSigSum[18] = ~io_mulAddResult[17];
  assign T141[17] = ~io_mulAddResult[16];
  assign T141[16] = ~io_mulAddResult[15];
  assign T141[15] = ~io_mulAddResult[14];
  assign T141[14] = ~io_mulAddResult[13];
  assign T141[13] = ~io_mulAddResult[12];
  assign T141[12] = ~io_mulAddResult[11];
  assign T141[11] = ~io_mulAddResult[10];
  assign T141[10] = ~io_mulAddResult[9];
  assign T141[9] = ~io_mulAddResult[8];
  assign T141[8] = ~io_mulAddResult[7];
  assign T141[7] = ~io_mulAddResult[6];
  assign T141[6] = ~io_mulAddResult[5];
  assign T141[5] = ~io_mulAddResult[4];
  assign T141[4] = ~io_mulAddResult[3];
  assign T141[3] = ~io_mulAddResult[2];
  assign T141[2] = ~io_mulAddResult[1];
  assign T141[1] = ~io_mulAddResult[0];
  assign T141[0] = ~io_fromPreMul_bit0AlignedNegSigC;
  assign CDom_firstNormAbsSigSum[41] = T162[41] | T154[41];
  assign CDom_firstNormAbsSigSum[40] = T162[40] | T154[40];
  assign CDom_firstNormAbsSigSum[39] = T162[39] | T154[39];
  assign CDom_firstNormAbsSigSum[38] = T162[38] | T154[38];
  assign CDom_firstNormAbsSigSum[37] = T162[37] | T154[37];
  assign CDom_firstNormAbsSigSum[36] = T162[36] | T154[36];
  assign CDom_firstNormAbsSigSum[35] = T162[35] | T154[35];
  assign CDom_firstNormAbsSigSum[34] = T162[34] | T154[34];
  assign CDom_firstNormAbsSigSum[33] = T162[33] | T154[33];
  assign CDom_firstNormAbsSigSum[32] = T162[32] | T154[32];
  assign CDom_firstNormAbsSigSum[31] = T162[31] | T154[31];
  assign CDom_firstNormAbsSigSum[30] = T162[30] | T154[30];
  assign CDom_firstNormAbsSigSum[29] = T162[29] | T154[29];
  assign CDom_firstNormAbsSigSum[28] = T162[28] | T154[28];
  assign CDom_firstNormAbsSigSum[27] = T162[27] | T154[27];
  assign CDom_firstNormAbsSigSum[26] = T162[26] | T154[26];
  assign CDom_firstNormAbsSigSum[25] = T162[25] | T154[25];
  assign CDom_firstNormAbsSigSum[24] = T162[24] | T154[24];
  assign CDom_firstNormAbsSigSum[23] = T162[23] | T154[23];
  assign CDom_firstNormAbsSigSum[22] = T162[22] | T154[22];
  assign CDom_firstNormAbsSigSum[21] = T162[21] | T154[21];
  assign CDom_firstNormAbsSigSum[20] = T162[20] | T154[20];
  assign CDom_firstNormAbsSigSum[19] = T162[19] | T154[19];
  assign CDom_firstNormAbsSigSum[18] = T162[18] | T154[18];
  assign CDom_firstNormAbsSigSum[17] = T162[17] | T154[17];
  assign CDom_firstNormAbsSigSum[16] = T162[16] | T154[16];
  assign CDom_firstNormAbsSigSum[15] = T162[15] | T154[15];
  assign CDom_firstNormAbsSigSum[14] = T162[14] | T154[14];
  assign CDom_firstNormAbsSigSum[13] = T162[13] | T154[13];
  assign CDom_firstNormAbsSigSum[12] = T162[12] | T154[12];
  assign CDom_firstNormAbsSigSum[11] = T162[11] | T154[11];
  assign CDom_firstNormAbsSigSum[10] = T162[10] | T154[10];
  assign CDom_firstNormAbsSigSum[9] = T162[9] | T154[9];
  assign CDom_firstNormAbsSigSum[8] = T162[8] | T154[8];
  assign CDom_firstNormAbsSigSum[7] = T162[7] | T154[7];
  assign CDom_firstNormAbsSigSum[6] = T162[6] | T154[6];
  assign CDom_firstNormAbsSigSum[5] = T162[5] | T154[5];
  assign CDom_firstNormAbsSigSum[4] = T162[4] | T154[4];
  assign CDom_firstNormAbsSigSum[3] = T162[3] | T154[3];
  assign CDom_firstNormAbsSigSum[2] = T162[2] | T154[2];
  assign CDom_firstNormAbsSigSum[1] = T162[1] | T154[1];
  assign CDom_firstNormAbsSigSum[0] = T162[0] | T154[0];
  assign T154[41] = T491[41] & notSigSum[58];
  assign T154[40] = T491[41] & notSigSum[57];
  assign T154[39] = T491[41] & notSigSum[56];
  assign T154[38] = T491[41] & notSigSum[55];
  assign T154[37] = T491[41] & notSigSum[54];
  assign T154[36] = T491[41] & notSigSum[53];
  assign T154[35] = T491[41] & notSigSum[52];
  assign T154[34] = T491[41] & notSigSum[51];
  assign T154[33] = T491[41] & notSigSum[50];
  assign T154[32] = T491[41] & notSigSum[49];
  assign T154[31] = T491[41] & notSigSum[48];
  assign T154[30] = T491[41] & notSigSum[47];
  assign T154[29] = T491[41] & notSigSum[46];
  assign T154[28] = T491[41] & notSigSum[45];
  assign T154[27] = T491[41] & notSigSum[44];
  assign T154[26] = T491[41] & notSigSum[43];
  assign T154[25] = T491[41] & notSigSum[42];
  assign T154[24] = T491[41] & notSigSum[41];
  assign T154[23] = T491[41] & notSigSum[40];
  assign T154[22] = T491[41] & notSigSum[39];
  assign T154[21] = T491[41] & notSigSum[38];
  assign T154[20] = T491[41] & notSigSum[37];
  assign T154[19] = T491[41] & notSigSum[36];
  assign T154[18] = T491[41] & notSigSum[35];
  assign T154[17] = T491[41] & notSigSum[34];
  assign T154[16] = T491[41] & notSigSum[33];
  assign T154[15] = T491[41] & notSigSum[32];
  assign T154[14] = T491[41] & notSigSum[31];
  assign T154[13] = T491[41] & notSigSum[30];
  assign T154[12] = T491[41] & notSigSum[29];
  assign T154[11] = T491[41] & notSigSum[28];
  assign T154[10] = T491[41] & notSigSum[27];
  assign T154[9] = T491[41] & notSigSum[26];
  assign T154[8] = T491[41] & notSigSum[25];
  assign T154[7] = T491[41] & notSigSum[24];
  assign T154[6] = T491[41] & notSigSum[23];
  assign T154[5] = T491[41] & notSigSum[22];
  assign T154[4] = T491[41] & notSigSum[21];
  assign T154[3] = T491[41] & notSigSum[20];
  assign T154[2] = T491[41] & notSigSum[19];
  assign T154[1] = T491[41] & notSigSum[18];
  assign T154[0] = T491[41] & N368;
  assign T491[41] = T159;
  assign T159 = T488[0] & CDom_estNormDist[4];
  assign T162[41] = T172[41] | T163[41];
  assign T162[40] = T172[40] | T163[40];
  assign T162[39] = T172[39] | T163[39];
  assign T162[38] = T172[38] | T163[38];
  assign T162[37] = T172[37] | T163[37];
  assign T162[36] = T172[36] | T163[36];
  assign T162[35] = T172[35] | T163[35];
  assign T162[34] = T172[34] | T163[34];
  assign T162[33] = T172[33] | T163[33];
  assign T162[32] = T172[32] | T163[32];
  assign T162[31] = T172[31] | T163[31];
  assign T162[30] = T172[30] | T163[30];
  assign T162[29] = T172[29] | T163[29];
  assign T162[28] = T172[28] | T163[28];
  assign T162[27] = T172[27] | T163[27];
  assign T162[26] = T172[26] | T163[26];
  assign T162[25] = T172[25] | T163[25];
  assign T162[24] = T172[24] | T163[24];
  assign T162[23] = T172[23] | T163[23];
  assign T162[22] = T172[22] | T163[22];
  assign T162[21] = T172[21] | T163[21];
  assign T162[20] = T172[20] | T163[20];
  assign T162[19] = T172[19] | T163[19];
  assign T162[18] = T172[18] | T163[18];
  assign T162[17] = T172[17] | T163[17];
  assign T162[16] = T172[16] | T163[16];
  assign T162[15] = T172[15] | T163[15];
  assign T162[14] = T172[14] | T163[14];
  assign T162[13] = T172[13] | T163[13];
  assign T162[12] = T172[12] | T163[12];
  assign T162[11] = T172[11] | T163[11];
  assign T162[10] = T172[10] | T163[10];
  assign T162[9] = T172[9] | T163[9];
  assign T162[8] = T172[8] | T163[8];
  assign T162[7] = T172[7] | T163[7];
  assign T162[6] = T172[6] | T163[6];
  assign T162[5] = T172[5] | T163[5];
  assign T162[4] = T172[4] | T163[4];
  assign T162[3] = T172[3] | T163[3];
  assign T162[2] = T172[2] | T163[2];
  assign T162[1] = T172[1] | T163[1];
  assign T162[0] = T172[0] | T163[0];
  assign T163[41] = T492[41] & notSigSum[74];
  assign T163[40] = T492[41] & notSigSum[73];
  assign T163[39] = T492[41] & notSigSum[72];
  assign T163[38] = T492[41] & notSigSum[71];
  assign T163[37] = T492[41] & notSigSum[70];
  assign T163[36] = T492[41] & notSigSum[69];
  assign T163[35] = T492[41] & notSigSum[68];
  assign T163[34] = T492[41] & notSigSum[67];
  assign T163[33] = T492[41] & notSigSum[66];
  assign T163[32] = T492[41] & notSigSum[65];
  assign T163[31] = T492[41] & notSigSum[64];
  assign T163[30] = T492[41] & notSigSum[63];
  assign T163[29] = T492[41] & notSigSum[62];
  assign T163[28] = T492[41] & notSigSum[61];
  assign T163[27] = T492[41] & notSigSum[60];
  assign T163[26] = T492[41] & notSigSum[59];
  assign T163[25] = T492[41] & notSigSum[58];
  assign T163[24] = T492[41] & notSigSum[57];
  assign T163[23] = T492[41] & notSigSum[56];
  assign T163[22] = T492[41] & notSigSum[55];
  assign T163[21] = T492[41] & notSigSum[54];
  assign T163[20] = T492[41] & notSigSum[53];
  assign T163[19] = T492[41] & notSigSum[52];
  assign T163[18] = T492[41] & notSigSum[51];
  assign T163[17] = T492[41] & notSigSum[50];
  assign T163[16] = T492[41] & notSigSum[49];
  assign T163[15] = T492[41] & notSigSum[48];
  assign T163[14] = T492[41] & notSigSum[47];
  assign T163[13] = T492[41] & notSigSum[46];
  assign T163[12] = T492[41] & notSigSum[45];
  assign T163[11] = T492[41] & notSigSum[44];
  assign T163[10] = T492[41] & notSigSum[43];
  assign T163[9] = T492[41] & notSigSum[42];
  assign T163[8] = T492[41] & notSigSum[41];
  assign T163[7] = T492[41] & notSigSum[40];
  assign T163[6] = T492[41] & notSigSum[39];
  assign T163[5] = T492[41] & notSigSum[38];
  assign T163[4] = T492[41] & notSigSum[37];
  assign T163[3] = T492[41] & notSigSum[36];
  assign T163[2] = T492[41] & notSigSum[35];
  assign T163[1] = T492[41] & notSigSum[34];
  assign T163[0] = T492[41] & N335;
  assign T492[41] = T168;
  assign T168 = T488[0] & T170;
  assign T170 = ~CDom_estNormDist[4];
  assign T172[41] = T182[41] | T173[41];
  assign T172[40] = T182[40] | T173[40];
  assign T172[39] = T182[39] | T173[39];
  assign T172[38] = T182[38] | T173[38];
  assign T172[37] = T182[37] | T173[37];
  assign T172[36] = T182[36] | T173[36];
  assign T172[35] = T182[35] | T173[35];
  assign T172[34] = T182[34] | T173[34];
  assign T172[33] = T182[33] | T173[33];
  assign T172[32] = T182[32] | T173[32];
  assign T172[31] = T182[31] | T173[31];
  assign T172[30] = T182[30] | T173[30];
  assign T172[29] = T182[29] | T173[29];
  assign T172[28] = T182[28] | T173[28];
  assign T172[27] = T182[27] | T173[27];
  assign T172[26] = T182[26] | T173[26];
  assign T172[25] = T182[25] | T173[25];
  assign T172[24] = T182[24] | T173[24];
  assign T172[23] = T182[23] | T173[23];
  assign T172[22] = T182[22] | T173[22];
  assign T172[21] = T182[21] | T173[21];
  assign T172[20] = T182[20] | T173[20];
  assign T172[19] = T182[19] | T173[19];
  assign T172[18] = T182[18] | T173[18];
  assign T172[17] = T182[17] | T173[17];
  assign T172[16] = T182[16] | T173[16];
  assign T172[15] = T182[15] | T173[15];
  assign T172[14] = T182[14] | T173[14];
  assign T172[13] = T182[13] | T173[13];
  assign T172[12] = T182[12] | T173[12];
  assign T172[11] = T182[11] | T173[11];
  assign T172[10] = T182[10] | T173[10];
  assign T172[9] = T182[9] | T173[9];
  assign T172[8] = T182[8] | T173[8];
  assign T172[7] = T182[7] | T173[7];
  assign T172[6] = T182[6] | T173[6];
  assign T172[5] = T182[5] | T173[5];
  assign T172[4] = T182[4] | T173[4];
  assign T172[3] = T182[3] | T173[3];
  assign T172[2] = T182[2] | T173[2];
  assign T172[1] = T182[1] | T173[1];
  assign T172[0] = T182[0] | T173[0];
  assign T173[41] = T493[41] & sigSum[58];
  assign T173[40] = T493[41] & sigSum[57];
  assign T173[39] = T493[41] & sigSum[56];
  assign T173[38] = T493[41] & sigSum[55];
  assign T173[37] = T493[41] & sigSum[54];
  assign T173[36] = T493[41] & sigSum[53];
  assign T173[35] = T493[41] & sigSum[52];
  assign T173[34] = T493[41] & sigSum[51];
  assign T173[33] = T493[41] & T21[50];
  assign T173[32] = T493[41] & T21[49];
  assign T173[31] = T493[41] & io_mulAddResult[47];
  assign T173[30] = T493[41] & io_mulAddResult[46];
  assign T173[29] = T493[41] & io_mulAddResult[45];
  assign T173[28] = T493[41] & io_mulAddResult[44];
  assign T173[27] = T493[41] & io_mulAddResult[43];
  assign T173[26] = T493[41] & io_mulAddResult[42];
  assign T173[25] = T493[41] & io_mulAddResult[41];
  assign T173[24] = T493[41] & io_mulAddResult[40];
  assign T173[23] = T493[41] & io_mulAddResult[39];
  assign T173[22] = T493[41] & io_mulAddResult[38];
  assign T173[21] = T493[41] & io_mulAddResult[37];
  assign T173[20] = T493[41] & io_mulAddResult[36];
  assign T173[19] = T493[41] & io_mulAddResult[35];
  assign T173[18] = T493[41] & io_mulAddResult[34];
  assign T173[17] = T493[41] & io_mulAddResult[33];
  assign T173[16] = T493[41] & io_mulAddResult[32];
  assign T173[15] = T493[41] & io_mulAddResult[31];
  assign T173[14] = T493[41] & io_mulAddResult[30];
  assign T173[13] = T493[41] & io_mulAddResult[29];
  assign T173[12] = T493[41] & io_mulAddResult[28];
  assign T173[11] = T493[41] & io_mulAddResult[27];
  assign T173[10] = T493[41] & io_mulAddResult[26];
  assign T173[9] = T493[41] & io_mulAddResult[25];
  assign T173[8] = T493[41] & io_mulAddResult[24];
  assign T173[7] = T493[41] & io_mulAddResult[23];
  assign T173[6] = T493[41] & io_mulAddResult[22];
  assign T173[5] = T493[41] & io_mulAddResult[21];
  assign T173[4] = T493[41] & io_mulAddResult[20];
  assign T173[3] = T493[41] & io_mulAddResult[19];
  assign T173[2] = T493[41] & io_mulAddResult[18];
  assign T173[1] = T493[41] & io_mulAddResult[17];
  assign T173[0] = T493[41] & N385;
  assign T493[41] = T178;
  assign T178 = T181 & CDom_estNormDist[4];
  assign T181 = ~T488[0];
  assign T182[41] = T494[41] & sigSum[74];
  assign T182[40] = T494[41] & sigSum[73];
  assign T182[39] = T494[41] & sigSum[72];
  assign T182[38] = T494[41] & sigSum[71];
  assign T182[37] = T494[41] & sigSum[70];
  assign T182[36] = T494[41] & sigSum[69];
  assign T182[35] = T494[41] & sigSum[68];
  assign T182[34] = T494[41] & sigSum[67];
  assign T182[33] = T494[41] & sigSum[66];
  assign T182[32] = T494[41] & sigSum[65];
  assign T182[31] = T494[41] & sigSum[64];
  assign T182[30] = T494[41] & sigSum[63];
  assign T182[29] = T494[41] & sigSum[62];
  assign T182[28] = T494[41] & sigSum[61];
  assign T182[27] = T494[41] & sigSum[60];
  assign T182[26] = T494[41] & sigSum[59];
  assign T182[25] = T494[41] & sigSum[58];
  assign T182[24] = T494[41] & sigSum[57];
  assign T182[23] = T494[41] & sigSum[56];
  assign T182[22] = T494[41] & sigSum[55];
  assign T182[21] = T494[41] & sigSum[54];
  assign T182[20] = T494[41] & sigSum[53];
  assign T182[19] = T494[41] & sigSum[52];
  assign T182[18] = T494[41] & sigSum[51];
  assign T182[17] = T494[41] & T21[50];
  assign T182[16] = T494[41] & T21[49];
  assign T182[15] = T494[41] & io_mulAddResult[47];
  assign T182[14] = T494[41] & io_mulAddResult[46];
  assign T182[13] = T494[41] & io_mulAddResult[45];
  assign T182[12] = T494[41] & io_mulAddResult[44];
  assign T182[11] = T494[41] & io_mulAddResult[43];
  assign T182[10] = T494[41] & io_mulAddResult[42];
  assign T182[9] = T494[41] & io_mulAddResult[41];
  assign T182[8] = T494[41] & io_mulAddResult[40];
  assign T182[7] = T494[41] & io_mulAddResult[39];
  assign T182[6] = T494[41] & io_mulAddResult[38];
  assign T182[5] = T494[41] & io_mulAddResult[37];
  assign T182[4] = T494[41] & io_mulAddResult[36];
  assign T182[3] = T494[41] & io_mulAddResult[35];
  assign T182[2] = T494[41] & io_mulAddResult[34];
  assign T182[1] = T494[41] & io_mulAddResult[33];
  assign T182[0] = T494[41] & N336;
  assign T494[41] = T187;
  assign T187 = T191 & T189;
  assign T189 = ~CDom_estNormDist[4];
  assign T191 = ~T488[0];
  assign T207[15] = T208[15] & absSigSumExtraMask[15];
  assign T207[14] = T208[14] & absSigSumExtraMask[14];
  assign T207[13] = T208[13] & absSigSumExtraMask[13];
  assign T207[12] = T208[12] & absSigSumExtraMask[12];
  assign T207[11] = T208[11] & absSigSumExtraMask[11];
  assign T207[10] = T208[10] & absSigSumExtraMask[10];
  assign T207[9] = T208[9] & absSigSumExtraMask[9];
  assign T207[8] = T208[8] & absSigSumExtraMask[8];
  assign T207[7] = T208[7] & T88[0];
  assign T207[6] = T208[6] & T88[1];
  assign T207[5] = T208[5] & T88[2];
  assign T207[4] = T208[4] & T88[3];
  assign T207[3] = T208[3] & T87[0];
  assign T207[2] = T208[2] & T87[1];
  assign T207[1] = T208[1] & absSigSumExtraMask_1;
  assign T207[0] = T208[0] & 1'b1;
  assign T208[15] = ~T125[15];
  assign T208[14] = ~T125[14];
  assign T208[13] = ~T125[13];
  assign T208[12] = ~T125[12];
  assign T208[11] = ~T125[11];
  assign T208[10] = ~T125[10];
  assign T208[9] = ~T125[9];
  assign T208[8] = ~T125[8];
  assign T208[7] = ~T125[7];
  assign T208[6] = ~T125[6];
  assign T208[5] = ~T125[5];
  assign T208[4] = ~T125[4];
  assign T208[3] = ~T125[3];
  assign T208[2] = ~T125[2];
  assign T208[1] = ~T125[1];
  assign T208[0] = ~T125[0];
  assign T212[27] = sigX3_27 & 1'b0;
  assign T212[26] = T374[0] & T498[26];
  assign T212[25] = sigX3[25] & T498[25];
  assign T212[24] = sigX3[24] & T498[24];
  assign T212[23] = sigX3[23] & T498[23];
  assign T212[22] = sigX3[22] & T498[22];
  assign T212[21] = sigX3[21] & T498[21];
  assign T212[20] = sigX3[20] & T498[20];
  assign T212[19] = sigX3[19] & T498[19];
  assign T212[18] = sigX3[18] & T498[18];
  assign T212[17] = sigX3[17] & T498[17];
  assign T212[16] = sigX3[16] & T498[16];
  assign T212[15] = sigX3[15] & T498[15];
  assign T212[14] = sigX3[14] & T498[14];
  assign T212[13] = sigX3[13] & T498[13];
  assign T212[12] = sigX3[12] & T498[12];
  assign T212[11] = sigX3[11] & T498[11];
  assign T212[10] = sigX3[10] & T498[10];
  assign T212[9] = sigX3[9] & T498[9];
  assign T212[8] = sigX3[8] & T498[8];
  assign T212[7] = sigX3[7] & T498[7];
  assign T212[6] = sigX3[6] & T498[6];
  assign T212[5] = sigX3[5] & T498[5];
  assign T212[4] = sigX3[4] & T498[4];
  assign T212[3] = sigX3[3] & T498[3];
  assign T212[2] = sigX3[2] & T498[2];
  assign T212[1] = sigX3[1] & T498[1];
  assign T212[0] = sigX3[0] & T498[0];
  assign T498[26] = 1'b0 & T373[25];
  assign T498[25] = T499[25] & T373[24];
  assign T498[24] = T499[24] & T373[23];
  assign T498[23] = T499[23] & T373[22];
  assign T498[22] = T499[22] & T373[21];
  assign T498[21] = T499[21] & T373[20];
  assign T498[20] = T499[20] & T373[19];
  assign T498[19] = T499[19] & T373[18];
  assign T498[18] = T499[18] & T373[17];
  assign T498[17] = T499[17] & T373[16];
  assign T498[16] = T499[16] & T373[15];
  assign T498[15] = T499[15] & T373[14];
  assign T498[14] = T499[14] & T373[13];
  assign T498[13] = T499[13] & T373[12];
  assign T498[12] = T499[12] & T373[11];
  assign T498[11] = T499[11] & T373[10];
  assign T498[10] = T499[10] & T373[9];
  assign T498[9] = T499[9] & T373[8];
  assign T498[8] = T499[8] & T373[7];
  assign T498[7] = T499[7] & T373[6];
  assign T498[6] = T499[6] & T373[5];
  assign T498[5] = T499[5] & T373[4];
  assign T498[4] = T499[4] & T373[3];
  assign T498[3] = T499[3] & T373[2];
  assign T498[2] = T499[2] & T373[1];
  assign T498[1] = T499[1] & T373[0];
  assign T498[0] = T499[0] & roundMask[0];
  assign T499[25] = ~T373[25];
  assign T499[24] = ~T373[24];
  assign T499[23] = ~T373[23];
  assign T499[22] = ~T373[22];
  assign T499[21] = ~T373[21];
  assign T499[20] = ~T373[20];
  assign T499[19] = ~T373[19];
  assign T499[18] = ~T373[18];
  assign T499[17] = ~T373[17];
  assign T499[16] = ~T373[16];
  assign T499[15] = ~T373[15];
  assign T499[14] = ~T373[14];
  assign T499[13] = ~T373[13];
  assign T499[12] = ~T373[12];
  assign T499[11] = ~T373[11];
  assign T499[10] = ~T373[10];
  assign T499[9] = ~T373[9];
  assign T499[8] = ~T373[8];
  assign T499[7] = ~T373[7];
  assign T499[6] = ~T373[6];
  assign T499[5] = ~T373[5];
  assign T499[4] = ~T373[4];
  assign T499[3] = ~T373[3];
  assign T499[2] = ~T373[2];
  assign T499[1] = ~T373[1];
  assign T499[0] = ~T373[0];
  assign T215 = ~allRound;
  assign allRound = N267 & N240;
  assign T216[27] = T218[27] & 1'b0;
  assign T216[26] = T218[26] & 1'b0;
  assign T216[25] = T218[25] & T373[25];
  assign T216[24] = T218[24] & T373[24];
  assign T216[23] = T218[23] & T373[23];
  assign T216[22] = T218[22] & T373[22];
  assign T216[21] = T218[21] & T373[21];
  assign T216[20] = T218[20] & T373[20];
  assign T216[19] = T218[19] & T373[19];
  assign T216[18] = T218[18] & T373[18];
  assign T216[17] = T218[17] & T373[17];
  assign T216[16] = T218[16] & T373[16];
  assign T216[15] = T218[15] & T373[15];
  assign T216[14] = T218[14] & T373[14];
  assign T216[13] = T218[13] & T373[13];
  assign T216[12] = T218[12] & T373[12];
  assign T216[11] = T218[11] & T373[11];
  assign T216[10] = T218[10] & T373[10];
  assign T216[9] = T218[9] & T373[9];
  assign T216[8] = T218[8] & T373[8];
  assign T216[7] = T218[7] & T373[7];
  assign T216[6] = T218[6] & T373[6];
  assign T216[5] = T218[5] & T373[5];
  assign T216[4] = T218[4] & T373[4];
  assign T216[3] = T218[3] & T373[3];
  assign T216[2] = T218[2] & T373[2];
  assign T216[1] = T218[1] & T373[1];
  assign T216[0] = T218[0] & T373[0];
  assign T218[27] = ~sigX3_27;
  assign T218[26] = ~T374[0];
  assign T218[25] = ~sigX3[25];
  assign T218[24] = ~sigX3[24];
  assign T218[23] = ~sigX3[23];
  assign T218[22] = ~sigX3[22];
  assign T218[21] = ~sigX3[21];
  assign T218[20] = ~sigX3[20];
  assign T218[19] = ~sigX3[19];
  assign T218[18] = ~sigX3[18];
  assign T218[17] = ~sigX3[17];
  assign T218[16] = ~sigX3[16];
  assign T218[15] = ~sigX3[15];
  assign T218[14] = ~sigX3[14];
  assign T218[13] = ~sigX3[13];
  assign T218[12] = ~sigX3[12];
  assign T218[11] = ~sigX3[11];
  assign T218[10] = ~sigX3[10];
  assign T218[9] = ~sigX3[9];
  assign T218[8] = ~sigX3[8];
  assign T218[7] = ~sigX3[7];
  assign T218[6] = ~sigX3[6];
  assign T218[5] = ~sigX3[5];
  assign T218[4] = ~sigX3[4];
  assign T218[3] = ~sigX3[3];
  assign T218[2] = ~sigX3[2];
  assign T218[1] = ~sigX3[1];
  assign T218[0] = ~sigX3[0];
  assign doIncrSig = T219 & T488[0];
  assign T219 = T221 & T220;
  assign T220 = ~sigSum[51];
  assign T221 = ~io_fromPreMul_isCDominant;
  assign commonCase = T223 & T222;
  assign T222 = ~notSpecial_addZeros;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & N334;
  assign T223 = ~addSpecial;
  assign addSpecial = mulSpecial | N208;
  assign mulSpecial = N209 | N210;
  assign io_exceptionFlags[1] = commonCase & underflowY;
  assign underflowY = inexactY & T227;
  assign T227 = sExpX3[10] | T228;
  assign N187 = ~sigX3Shift1;
  assign T501[1] = sigX3Shift1;
  assign T501[0] = N187;
  assign io_exceptionFlags[2] = commonCase & N207;
  assign T232[2] = T280[9] | T233[9];
  assign T232[1] = T280[8] | T233[8];
  assign T232[0] = T280[7] | T233[7];
  assign sExpY[6] = T280[6] | T233[6];
  assign sExpY[5] = T280[5] | T233[5];
  assign sExpY[4] = T280[4] | T233[4];
  assign sExpY[3] = T280[3] | T233[3];
  assign sExpY[2] = T280[2] | T233[2];
  assign sExpY[1] = T280[1] | T233[1];
  assign sExpY[0] = T280[0] | T233[0];
  assign T236[1] = T250[25] | T237[25];
  assign T236[0] = T250[24] | T237[24];
  assign sigY3[23] = T250[23] | T237[23];
  assign sigY3[22] = T250[22] | T237[22];
  assign sigY3[21] = T250[21] | T237[21];
  assign sigY3[20] = T250[20] | T237[20];
  assign sigY3[19] = T250[19] | T237[19];
  assign sigY3[18] = T250[18] | T237[18];
  assign sigY3[17] = T250[17] | T237[17];
  assign sigY3[16] = T250[16] | T237[16];
  assign sigY3[15] = T250[15] | T237[15];
  assign sigY3[14] = T250[14] | T237[14];
  assign sigY3[13] = T250[13] | T237[13];
  assign sigY3[12] = T250[12] | T237[12];
  assign sigY3[11] = T250[11] | T237[11];
  assign sigY3[10] = T250[10] | T237[10];
  assign sigY3[9] = T250[9] | T237[9];
  assign sigY3[8] = T250[8] | T237[8];
  assign sigY3[7] = T250[7] | T237[7];
  assign sigY3[6] = T250[6] | T237[6];
  assign sigY3[5] = T250[5] | T237[5];
  assign sigY3[4] = T250[4] | T237[4];
  assign sigY3[3] = T250[3] | T237[3];
  assign sigY3[2] = T250[2] | T237[2];
  assign sigY3[1] = T250[1] | T237[1];
  assign sigY3[0] = T250[0] | T237[0];
  assign N188 = ~roundEven;
  assign T238[25] = roundUp_sigY3[25] & T239[25];
  assign T238[24] = roundUp_sigY3[24] & T239[24];
  assign T238[23] = roundUp_sigY3[23] & T239[23];
  assign T238[22] = roundUp_sigY3[22] & T239[22];
  assign T238[21] = roundUp_sigY3[21] & T239[21];
  assign T238[20] = roundUp_sigY3[20] & T239[20];
  assign T238[19] = roundUp_sigY3[19] & T239[19];
  assign T238[18] = roundUp_sigY3[18] & T239[18];
  assign T238[17] = roundUp_sigY3[17] & T239[17];
  assign T238[16] = roundUp_sigY3[16] & T239[16];
  assign T238[15] = roundUp_sigY3[15] & T239[15];
  assign T238[14] = roundUp_sigY3[14] & T239[14];
  assign T238[13] = roundUp_sigY3[13] & T239[13];
  assign T238[12] = roundUp_sigY3[12] & T239[12];
  assign T238[11] = roundUp_sigY3[11] & T239[11];
  assign T238[10] = roundUp_sigY3[10] & T239[10];
  assign T238[9] = roundUp_sigY3[9] & T239[9];
  assign T238[8] = roundUp_sigY3[8] & T239[8];
  assign T238[7] = roundUp_sigY3[7] & T239[7];
  assign T238[6] = roundUp_sigY3[6] & T239[6];
  assign T238[5] = roundUp_sigY3[5] & T239[5];
  assign T238[4] = roundUp_sigY3[4] & T239[4];
  assign T238[3] = roundUp_sigY3[3] & T239[3];
  assign T238[2] = roundUp_sigY3[2] & T239[2];
  assign T238[1] = roundUp_sigY3[1] & T239[1];
  assign T238[0] = roundUp_sigY3[0] & T239[0];
  assign T239[25] = ~T373[25];
  assign T239[24] = ~T373[24];
  assign T239[23] = ~T373[23];
  assign T239[22] = ~T373[22];
  assign T239[21] = ~T373[21];
  assign T239[20] = ~T373[20];
  assign T239[19] = ~T373[19];
  assign T239[18] = ~T373[18];
  assign T239[17] = ~T373[17];
  assign T239[16] = ~T373[16];
  assign T239[15] = ~T373[15];
  assign T239[14] = ~T373[14];
  assign T239[13] = ~T373[13];
  assign T239[12] = ~T373[12];
  assign T239[11] = ~T373[11];
  assign T239[10] = ~T373[10];
  assign T239[9] = ~T373[9];
  assign T239[8] = ~T373[8];
  assign T239[7] = ~T373[7];
  assign T239[6] = ~T373[6];
  assign T239[5] = ~T373[5];
  assign T239[4] = ~T373[4];
  assign T239[3] = ~T373[3];
  assign T239[2] = ~T373[2];
  assign T239[1] = ~T373[1];
  assign T239[0] = ~T373[0];
  assign T242[25] = sigX3_27 | 1'b0;
  assign T242[24] = T374[0] | T373[25];
  assign T242[23] = sigX3[25] | T373[24];
  assign T242[22] = sigX3[24] | T373[23];
  assign T242[21] = sigX3[23] | T373[22];
  assign T242[20] = sigX3[22] | T373[21];
  assign T242[19] = sigX3[21] | T373[20];
  assign T242[18] = sigX3[20] | T373[19];
  assign T242[17] = sigX3[19] | T373[18];
  assign T242[16] = sigX3[18] | T373[17];
  assign T242[15] = sigX3[17] | T373[16];
  assign T242[14] = sigX3[16] | T373[15];
  assign T242[13] = sigX3[15] | T373[14];
  assign T242[12] = sigX3[14] | T373[13];
  assign T242[11] = sigX3[13] | T373[12];
  assign T242[10] = sigX3[12] | T373[11];
  assign T242[9] = sigX3[11] | T373[10];
  assign T242[8] = sigX3[10] | T373[9];
  assign T242[7] = sigX3[9] | T373[8];
  assign T242[6] = sigX3[8] | T373[7];
  assign T242[5] = sigX3[7] | T373[6];
  assign T242[4] = sigX3[6] | T373[5];
  assign T242[3] = sigX3[5] | T373[4];
  assign T242[2] = sigX3[4] | T373[3];
  assign T242[1] = sigX3[3] | T373[2];
  assign T242[0] = sigX3[2] | T373[1];
  assign T244 = T246 & T245;
  assign T245 = ~N294;
  assign T246 = N296 & N267;
  assign T247 = T248 & N240;
  assign T248 = N296 & T249;
  assign T249 = ~N267;
  assign T250[25] = T272[25] | T251[25];
  assign T250[24] = T272[24] | T251[24];
  assign T250[23] = T272[23] | T251[23];
  assign T250[22] = T272[22] | T251[22];
  assign T250[21] = T272[21] | T251[21];
  assign T250[20] = T272[20] | T251[20];
  assign T250[19] = T272[19] | T251[19];
  assign T250[18] = T272[18] | T251[18];
  assign T250[17] = T272[17] | T251[17];
  assign T250[16] = T272[16] | T251[16];
  assign T250[15] = T272[15] | T251[15];
  assign T250[14] = T272[14] | T251[14];
  assign T250[13] = T272[13] | T251[13];
  assign T250[12] = T272[12] | T251[12];
  assign T250[11] = T272[11] | T251[11];
  assign T250[10] = T272[10] | T251[10];
  assign T250[9] = T272[9] | T251[9];
  assign T250[8] = T272[8] | T251[8];
  assign T250[7] = T272[7] | T251[7];
  assign T250[6] = T272[6] | T251[6];
  assign T250[5] = T272[5] | T251[5];
  assign T250[4] = T272[4] | T251[4];
  assign T250[3] = T272[3] | T251[3];
  assign T250[2] = T272[2] | T251[2];
  assign T250[1] = T272[1] | T251[1];
  assign T250[0] = T272[0] | T251[0];
  assign N189 = ~T252;
  assign T252 = T259 | T253;
  assign T253 = doIncrSig & roundDirectUp;
  assign N190 = ~signY;
  assign N191 = ~isZeroY;
  assign T255 = io_fromPreMul_signProd ^ doNegSignSum;
  assign N192 = ~io_fromPreMul_isCDominant;
  assign T256 = T488[0] & T257;
  assign T257 = ~N334;
  assign T259 = T262 | T260;
  assign T260 = T261 & N267;
  assign T261 = doIncrSig & N296;
  assign T262 = T264 | T263;
  assign T263 = doIncrSig & allRound;
  assign T264 = T268 | T265;
  assign T265 = T266 & anyRound;
  assign T266 = T267 & roundDirectUp;
  assign T267 = ~doIncrSig;
  assign T268 = T269 & N294;
  assign T269 = T270 & N267;
  assign T270 = T271 & N296;
  assign T271 = ~doIncrSig;
  assign N193 = ~T276;
  assign T273[25] = sigX3_27 & 1'b0;
  assign T273[24] = T374[0] & T503[26];
  assign T273[23] = sigX3[25] & T503[25];
  assign T273[22] = sigX3[24] & T503[24];
  assign T273[21] = sigX3[23] & T503[23];
  assign T273[20] = sigX3[22] & T503[22];
  assign T273[19] = sigX3[21] & T503[21];
  assign T273[18] = sigX3[20] & T503[20];
  assign T273[17] = sigX3[19] & T503[19];
  assign T273[16] = sigX3[18] & T503[18];
  assign T273[15] = sigX3[17] & T503[17];
  assign T273[14] = sigX3[16] & T503[16];
  assign T273[13] = sigX3[15] & T503[15];
  assign T273[12] = sigX3[14] & T503[14];
  assign T273[11] = sigX3[13] & T503[13];
  assign T273[10] = sigX3[12] & T503[12];
  assign T273[9] = sigX3[11] & T503[11];
  assign T273[8] = sigX3[10] & T503[10];
  assign T273[7] = sigX3[9] & T503[9];
  assign T273[6] = sigX3[8] & T503[8];
  assign T273[5] = sigX3[7] & T503[7];
  assign T273[4] = sigX3[6] & T503[6];
  assign T273[3] = sigX3[5] & T503[5];
  assign T273[2] = sigX3[4] & T503[4];
  assign T273[1] = sigX3[3] & T503[3];
  assign T273[0] = sigX3[2] & T503[2];
  assign T503[26] = ~T373[25];
  assign T503[25] = ~T373[24];
  assign T503[24] = ~T373[23];
  assign T503[23] = ~T373[22];
  assign T503[22] = ~T373[21];
  assign T503[21] = ~T373[20];
  assign T503[20] = ~T373[19];
  assign T503[19] = ~T373[18];
  assign T503[18] = ~T373[17];
  assign T503[17] = ~T373[16];
  assign T503[16] = ~T373[15];
  assign T503[15] = ~T373[14];
  assign T503[14] = ~T373[13];
  assign T503[13] = ~T373[12];
  assign T503[12] = ~T373[11];
  assign T503[11] = ~T373[10];
  assign T503[10] = ~T373[9];
  assign T503[9] = ~T373[8];
  assign T503[8] = ~T373[7];
  assign T503[7] = ~T373[6];
  assign T503[6] = ~T373[5];
  assign T503[5] = ~T373[4];
  assign T503[4] = ~T373[3];
  assign T503[3] = ~T373[2];
  assign T503[2] = ~T373[1];
  assign T276 = T279 & T278;
  assign T278 = ~roundEven;
  assign T279 = ~T252;
  assign T280[9] = T283[9] | T281[9];
  assign T280[8] = T283[8] | T281[8];
  assign T280[7] = T283[7] | T281[7];
  assign T280[6] = T283[6] | T281[6];
  assign T280[5] = T283[5] | T281[5];
  assign T280[4] = T283[4] | T281[4];
  assign T280[3] = T283[3] | T281[3];
  assign T280[2] = T283[2] | T281[2];
  assign T280[1] = T283[1] | T281[1];
  assign T280[0] = T283[0] | T281[0];
  assign N194 = ~T236[0];
  assign N195 = ~T236[1];
  assign io_exceptionFlags[4] = T305 | notSigNaN_invalid;
  assign notSigNaN_invalid = T302 | T287;
  assign T287 = T288 & T488[0];
  assign T288 = T291 & isInfC;
  assign isInfC = N208 & T289;
  assign T289 = ~io_fromPreMul_highExpC[0];
  assign T291 = T297 & T292;
  assign T292 = isInfA | isInfB;
  assign isInfB = N210 & T293;
  assign T293 = ~io_fromPreMul_highExpB[0];
  assign isInfA = N209 & T295;
  assign T295 = ~io_fromPreMul_highExpA[0];
  assign T297 = T300 & T298;
  assign T298 = ~isNaNB;
  assign isNaNB = N210 & io_fromPreMul_highExpB[0];
  assign T300 = ~isNaNA;
  assign isNaNA = N209 & io_fromPreMul_highExpA[0];
  assign T302 = T304 | T303;
  assign T303 = N202 & isInfB;
  assign T304 = isInfA & N199;
  assign T305 = T308 | isSigNaNC;
  assign isSigNaNC = isNaNC & T306;
  assign T306 = ~io_fromPreMul_isNaN_isQuietNaNC;
  assign isNaNC = N208 & io_fromPreMul_highExpC[0];
  assign T308 = isSigNaNA | isSigNaNB;
  assign isSigNaNB = isNaNB & T309;
  assign T309 = ~io_fromPreMul_isNaN_isQuietNaNB;
  assign isSigNaNA = isNaNA & T310;
  assign T310 = ~io_fromPreMul_isNaN_isQuietNaNA;
  assign io_out[22] = T318[22] | T313[22];
  assign io_out[21] = T318[21] | T313[22];
  assign io_out[20] = T318[20] | T313[22];
  assign io_out[19] = T318[19] | T313[22];
  assign io_out[18] = T318[18] | T313[22];
  assign io_out[17] = T318[17] | T313[22];
  assign io_out[16] = T318[16] | T313[22];
  assign io_out[15] = T318[15] | T313[22];
  assign io_out[14] = T318[14] | T313[22];
  assign io_out[13] = T318[13] | T313[22];
  assign io_out[12] = T318[12] | T313[22];
  assign io_out[11] = T318[11] | T313[22];
  assign io_out[10] = T318[10] | T313[22];
  assign io_out[9] = T318[9] | T313[22];
  assign io_out[8] = T318[8] | T313[22];
  assign io_out[7] = T318[7] | T313[22];
  assign io_out[6] = T318[6] | T313[22];
  assign io_out[5] = T318[5] | T313[22];
  assign io_out[4] = T318[4] | T313[22];
  assign io_out[3] = T318[3] | T313[22];
  assign io_out[2] = T318[2] | T313[22];
  assign io_out[1] = T318[1] | T313[22];
  assign io_out[0] = T318[0] | T313_0;
  assign T504[0] = io_exceptionFlags[2] & T314;
  assign T314 = ~overflowY_roundMagUp;
  assign overflowY_roundMagUp = N296 | roundMagUp;
  assign roundMagUp = T317 | T315;
  assign T315 = N297 & T316;
  assign T316 = ~signY;
  assign T317 = N331 & signY;
  assign T318[22] = T322[22] | T319[22];
  assign T318[21] = T322[21] | 1'b0;
  assign T318[20] = T322[20] | 1'b0;
  assign T318[19] = T322[19] | 1'b0;
  assign T318[18] = T322[18] | 1'b0;
  assign T318[17] = T322[17] | 1'b0;
  assign T318[16] = T322[16] | 1'b0;
  assign T318[15] = T322[15] | 1'b0;
  assign T318[14] = T322[14] | 1'b0;
  assign T318[13] = T322[13] | 1'b0;
  assign T318[12] = T322[12] | 1'b0;
  assign T318[11] = T322[11] | 1'b0;
  assign T318[10] = T322[10] | 1'b0;
  assign T318[9] = T322[9] | 1'b0;
  assign T318[8] = T322[8] | 1'b0;
  assign T318[7] = T322[7] | 1'b0;
  assign T318[6] = T322[6] | 1'b0;
  assign T318[5] = T322[5] | 1'b0;
  assign T318[4] = T322[4] | 1'b0;
  assign T318[3] = T322[3] | 1'b0;
  assign T318[2] = T322[2] | 1'b0;
  assign T318[1] = T322[1] | 1'b0;
  assign T318[0] = T322[0] | 1'b0;
  assign T319[22] = T320 | notSigNaN_invalid;
  assign T320 = T321 | isNaNC;
  assign T321 = isNaNA | isNaNB;
  assign N196 = ~T325;
  assign T325 = T326 | T319[22];
  assign T326 = totalUnderflowY & roundMagUp;
  assign totalUnderflowY = T331 & T327;
  assign T327 = T232[2] | T328;
  assign T331 = ~isZeroY;
  assign io_out[31] = T333[8] | T332[8];
  assign io_out[30] = T333[7] | T332[8];
  assign io_out[29] = T333[6] | T332[8];
  assign io_out[28] = T333[5] | 1'b0;
  assign io_out[27] = T333[4] | 1'b0;
  assign io_out[26] = T333[3] | 1'b0;
  assign io_out[25] = T333[2] | 1'b0;
  assign io_out[24] = T333[1] | 1'b0;
  assign io_out[23] = T333[0] | 1'b0;
  assign T332[8] = T319[22];
  assign T333[8] = T338[8] | T334[8];
  assign T333[7] = T338[7] | T334[8];
  assign T333[6] = T338[6] | 1'b0;
  assign T333[5] = T338[5] | 1'b0;
  assign T333[4] = T338[4] | 1'b0;
  assign T333[3] = T338[3] | 1'b0;
  assign T333[2] = T338[2] | 1'b0;
  assign T333[1] = T338[1] | 1'b0;
  assign T333[0] = T338[0] | 1'b0;
  assign T334[8] = notNaN_isInfOut;
  assign notNaN_isInfOut = T336 | T335;
  assign T335 = io_exceptionFlags[2] & overflowY_roundMagUp;
  assign T336 = T337 | isInfC;
  assign T337 = isInfA | isInfB;
  assign T338[8] = T340[8] | T339[8];
  assign T338[7] = T340[7] | 1'b0;
  assign T338[6] = T340[6] | T339[8];
  assign T338[5] = T340[5] | T339[8];
  assign T338[4] = T340[4] | T339[8];
  assign T338[3] = T340[3] | T339[8];
  assign T338[2] = T340[2] | T339[8];
  assign T338[1] = T340[1] | T339[8];
  assign T338[0] = T340[0] | T339[8];
  assign T339[8] = T504[0];
  assign T340[8] = T343[8] | 1'b0;
  assign T340[7] = T343[7] | 1'b0;
  assign T340[6] = T343[6] | T341[6];
  assign T340[5] = T343[5] | T341[6];
  assign T340[4] = T343[4] | 1'b0;
  assign T340[3] = T343[3] | T341[6];
  assign T340[2] = T343[2] | 1'b0;
  assign T340[1] = T343[1] | T341[6];
  assign T340[0] = T343[0] | T341[6];
  assign T341[6] = pegMinFiniteMagOut;
  assign pegMinFiniteMagOut = T342 & roundMagUp;
  assign T342 = commonCase & totalUnderflowY;
  assign T343[8] = T346[8] & T344[8];
  assign T343[7] = T346[7] & T344[7];
  assign T343[6] = T346[6] & T344[6];
  assign T343[5] = T346[5] & T344[5];
  assign T343[4] = T346[4] & T344[4];
  assign T343[3] = T346[3] & T344[3];
  assign T343[2] = T346[2] & T344[2];
  assign T343[1] = T346[1] & T344[1];
  assign T343[0] = T346[0] & T344[0];
  assign T344[8] = ~1'b0;
  assign T344[7] = ~1'b0;
  assign T344[6] = ~T345[6];
  assign T344[5] = ~1'b0;
  assign T344[4] = ~1'b0;
  assign T344[3] = ~1'b0;
  assign T344[2] = ~1'b0;
  assign T344[1] = ~1'b0;
  assign T344[0] = ~1'b0;
  assign T345[6] = notNaN_isInfOut;
  assign T346[8] = T349[8] & T347[8];
  assign T346[7] = T349[7] & T347[7];
  assign T346[6] = T349[6] & T347[6];
  assign T346[5] = T349[5] & T347[5];
  assign T346[4] = T349[4] & T347[4];
  assign T346[3] = T349[3] & T347[3];
  assign T346[2] = T349[2] & T347[2];
  assign T346[1] = T349[1] & T347[1];
  assign T346[0] = T349[0] & T347[0];
  assign T347[8] = ~1'b0;
  assign T347[7] = ~T348[7];
  assign T347[6] = ~1'b0;
  assign T347[5] = ~1'b0;
  assign T347[4] = ~1'b0;
  assign T347[3] = ~1'b0;
  assign T347[2] = ~1'b0;
  assign T347[1] = ~1'b0;
  assign T347[0] = ~1'b0;
  assign T348[7] = T504[0];
  assign T349[8] = T352[8] & T350[8];
  assign T349[7] = T352[7] & T350[7];
  assign T349[6] = T352[6] & T350[6];
  assign T349[5] = T352[5] & T350[5];
  assign T349[4] = T352[4] & T350[4];
  assign T349[3] = T352[3] & T350[3];
  assign T349[2] = T352[2] & T350[2];
  assign T349[1] = T352[1] & T350[1];
  assign T349[0] = T352[0] & T350[0];
  assign T350[8] = ~T351[8];
  assign T350[7] = ~T351[8];
  assign T350[6] = ~1'b0;
  assign T350[5] = ~1'b0;
  assign T350[4] = ~T351[8];
  assign T350[3] = ~1'b0;
  assign T350[2] = ~T351[8];
  assign T350[1] = ~1'b0;
  assign T350[0] = ~1'b0;
  assign T351[8] = pegMinFiniteMagOut;
  assign T352[8] = T232[1] & T353[8];
  assign T352[7] = T232[0] & T353[7];
  assign T352[6] = sExpY[6] & T353[6];
  assign T352[5] = sExpY[5] & T353[5];
  assign T352[4] = sExpY[4] & T353[4];
  assign T352[3] = sExpY[3] & T353[3];
  assign T352[2] = sExpY[2] & T353[2];
  assign T352[1] = sExpY[1] & T353[1];
  assign T352[0] = sExpY[0] & T353[0];
  assign T353[8] = ~T354[8];
  assign T353[7] = ~T354[8];
  assign T353[6] = ~T354[8];
  assign T353[5] = ~1'b0;
  assign T353[4] = ~1'b0;
  assign T353[3] = ~1'b0;
  assign T353[2] = ~1'b0;
  assign T353[1] = ~1'b0;
  assign T353[0] = ~1'b0;
  assign T354[8] = notSpecial_isZeroOut;
  assign notSpecial_isZeroOut = T355 | totalUnderflowY;
  assign T355 = notSpecial_addZeros | isZeroY;
  assign io_out[32] = T357 | T356;
  assign T356 = commonCase & signY;
  assign T357 = T372 & uncommonCaseSignOut;
  assign uncommonCaseSignOut = T362 | T358;
  assign T358 = T359 & N331;
  assign T359 = T360 & T488[0];
  assign T360 = T361 & notSpecial_addZeros;
  assign T361 = ~mulSpecial;
  assign T362 = T366 | T363;
  assign T363 = T364 & io_fromPreMul_opSignC;
  assign T364 = T365 & N208;
  assign T365 = ~mulSpecial;
  assign T366 = T370 | T367;
  assign T367 = T368 & io_fromPreMul_signProd;
  assign T368 = mulSpecial & T369;
  assign T369 = ~N208;
  assign T370 = T371 & io_fromPreMul_opSignC;
  assign T371 = ~T488[0];
  assign T372 = ~T319[22];

endmodule