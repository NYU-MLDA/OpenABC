module bp_fe_bht_bht_idx_width_p9
(
  clk_i,
  reset_i,
  w_v_i,
  idx_w_i,
  correct_i,
  r_v_i,
  idx_r_i,
  predict_o
);

  input [8:0] idx_w_i;
  input [8:0] idx_r_i;
  input clk_i;
  input reset_i;
  input w_v_i;
  input correct_i;
  input r_v_i;
  output predict_o;
  wire predict_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,
  N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,
  N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,
  N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,
  N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,
  N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,
  N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,
  N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,
  N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,
  N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,
  N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,
  N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,
  N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,
  N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,
  N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,
  N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,
  N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,
  N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
  N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,
  N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,
  N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,
  N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,
  N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,
  N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,
  N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,
  N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,
  N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,
  N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,
  N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,
  N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,
  N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,
  N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,
  N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,
  N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,
  N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,
  N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,
  N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,
  N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,
  N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,
  N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,
  N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,
  N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,
  N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,
  N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,
  N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,
  N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,
  N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
  N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,
  N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,
  N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,
  N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,
  N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,
  N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,
  N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,
  N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,
  N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,
  N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,
  N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,
  N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,
  N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,
  N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,
  N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,
  N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,
  N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,
  N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,
  N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,
  N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,
  N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,
  N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,
  N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,
  N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,
  N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,
  N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,
  N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,
  N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,
  N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,
  N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,
  N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,
  N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,
  N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,
  N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,
  N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,
  N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,
  N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,
  N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,
  N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,
  N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,
  N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,
  N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,
  N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,
  N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,
  N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,
  N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,
  N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,
  N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,
  N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,
  N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,
  N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,
  N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,
  N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,
  N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,
  N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,
  N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,
  N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,
  N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,
  N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,
  N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,
  N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,
  N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,
  N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,
  N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,
  N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,
  N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,
  N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,
  N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,
  N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,
  N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,
  N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,
  N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,
  N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,
  N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,
  N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,
  N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,
  N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,
  N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,
  N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,
  N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,
  N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,
  N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,
  N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,
  N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,
  N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,
  N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,
  N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,
  N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,
  N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,
  N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,
  N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,
  N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
  N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,
  N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,
  N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,
  N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,
  N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,
  N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,
  N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,
  N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,
  N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,
  N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,
  N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,
  N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,
  N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
  N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,
  N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,
  N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
  N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,
  N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,
  N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
  N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,
  N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,
  N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,
  N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,
  N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,
  N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,
  N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,
  N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,
  N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,
  N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,
  N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,
  N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,
  N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,
  N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,
  N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,
  N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,
  N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,
  N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,
  N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,
  N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,
  N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,
  N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,
  N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,
  N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,
  N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,
  N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,
  N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,
  N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,
  N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,
  N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,
  N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,
  N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,
  N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,
  N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,
  N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,
  N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,
  N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,
  N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,
  N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,
  N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,
  N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,
  N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,
  N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,
  N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,
  N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,
  N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,
  N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,
  N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,
  N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,
  N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,
  N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,
  N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,
  N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,
  N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,
  N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,
  N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,
  N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,
  N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,
  N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,
  N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,
  N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,
  N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,
  N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,
  N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,
  N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,
  N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,
  N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,
  N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,
  N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,
  N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,
  N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,
  N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,
  N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,
  N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,
  N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,
  N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,
  N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,
  N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,
  N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,
  N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,
  N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,
  N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,
  N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,
  N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,
  N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,
  N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,
  N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,
  N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,
  N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,
  N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,
  N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,
  N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,
  N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,
  N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,
  N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,
  N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,
  N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,
  N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,
  N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,
  N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,
  N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,
  N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,
  N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,
  N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,
  N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,
  N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,
  N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,
  N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,
  N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,
  N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,
  N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,
  N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,
  N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,
  N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,
  N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,
  N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,
  N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,
  N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,
  N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,
  N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,
  N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,
  N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,
  N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,
  N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,
  N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,
  N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,
  N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,
  N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,
  N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,
  N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,
  N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,
  N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,
  N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,
  N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,
  N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,
  N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,
  N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,
  N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,
  N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,
  N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,
  N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,
  N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,
  N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,
  N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,
  N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,
  N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,
  N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,
  N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,
  N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,
  N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,
  N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,
  N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,
  N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,
  N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,
  N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,
  N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,
  N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,
  N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,
  N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,
  N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,
  N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,
  N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,
  N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,
  N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,
  N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,
  N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,
  N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,
  N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,
  N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,
  N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,
  N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,
  N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,
  N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,
  N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,
  N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,
  N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,
  N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,
  N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,
  N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,
  N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,
  N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,
  N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,
  N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,
  N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,
  N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,
  N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,
  N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,
  N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,
  N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,
  N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,
  N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,
  N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,
  N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,
  N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,
  N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,
  N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,
  N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,
  N5956,N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,
  N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,
  N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,
  N5996,N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,
  N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,
  N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,
  N6036,N6037,N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,
  N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,
  N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,
  N6076,N6077,N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,
  N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,
  N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,
  N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,
  N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,
  N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,
  N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,
  N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,
  N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,
  N6196,N6197,N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,
  N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,
  N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6235,
  N6236,N6237,N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,
  N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,
  N6263,N6264,N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,N6274,N6275,
  N6276,N6277,N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,
  N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,
  N6303,N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,N6314,N6315,
  N6316,N6317,N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,
  N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,
  N6343,N6344,N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354,N6355,
  N6356,N6357,N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,
  N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,
  N6383,N6384,N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394,N6395,
  N6396,N6397,N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,
  N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,
  N6423,N6424,N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,N6434,N6435,
  N6436,N6437,N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,
  N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,
  N6463,N6464,N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,N6474,N6475,
  N6476,N6477,N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,
  N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,
  N6503,N6504,N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514,N6515,
  N6516,N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,
  N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,
  N6543,N6544,N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,N6554,N6555,
  N6556,N6557,N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,
  N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,
  N6583,N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,N6594,N6595,
  N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,
  N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,
  N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,N6634,N6635,
  N6636,N6637,N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,
  N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,
  N6663,N6664,N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,N6674,N6675,
  N6676,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,
  N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,
  N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,
  N6716,N6717,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,
  N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,
  N6743,N6744,N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,N6754,N6755,
  N6756,N6757,N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,
  N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,
  N6783,N6784,N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,
  N6796,N6797,N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,
  N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,
  N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,N6834,N6835,
  N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,
  N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,
  N6863,N6864,N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,N6874,N6875,
  N6876,N6877,N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,
  N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,
  N6903,N6904,N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,N6914,N6915,
  N6916,N6917,N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,
  N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,
  N6943,N6944,N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,N6954,N6955,
  N6956,N6957,N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,
  N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,
  N6983,N6984,N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,N6994,N6995,
  N6996,N6997,N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,
  N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,
  N7023,N7024,N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,N7034,N7035,
  N7036,N7037,N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,
  N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,
  N7063,N7064,N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,N7074,N7075,
  N7076,N7077,N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,
  N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,
  N7103,N7104,N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,N7114,N7115,
  N7116,N7117,N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,
  N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,
  N7143,N7144,N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,N7154,N7155,
  N7156,N7157,N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,
  N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,
  N7183,N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,N7193,N7194,N7195,
  N7196,N7197,N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,
  N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,
  N7223,N7224,N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,N7233,N7234,N7235,
  N7236,N7237,N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,
  N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,
  N7263,N7264,N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,N7273,N7274,N7275,
  N7276,N7277,N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,
  N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,
  N7303,N7304,N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,N7313,N7314,N7315,
  N7316,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,
  N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,
  N7343,N7344,N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,N7353,N7354,N7355,
  N7356,N7357,N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,
  N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,
  N7383,N7384,N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,N7393,N7394,N7395,
  N7396,N7397,N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,
  N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,
  N7423,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7433,N7434,N7435,
  N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7449,
  N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,
  N7463,N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,N7473,N7474,N7475,
  N7476,N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,
  N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,N7500,N7501,N7502,
  N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,N7513,N7514,N7515,
  N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,N7529,
  N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,N7540,N7541,N7542,
  N7543,N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,N7553,N7554,N7555,
  N7556,N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7569,
  N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580,N7581,N7582,
  N7583,N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,N7593,N7594,N7595,
  N7596,N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,N7609,
  N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,N7620,N7621,N7622,
  N7623,N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633,N7634,N7635,
  N7636,N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,N7649,
  N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661,N7662,
  N7663,N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,
  N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,
  N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7702,
  N7703,N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,N7713,N7714,N7715,
  N7716,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,N7729,
  N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,
  N7743,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,N7753,N7754,N7755,
  N7756,N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,N7769,
  N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,N7780,N7781,N7782,
  N7783,N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,N7793,N7794,N7795,
  N7796,N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,N7809,
  N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,N7820,N7821,N7822,
  N7823,N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,N7833,N7834,N7835,
  N7836,N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,N7849,
  N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,N7860,N7861,N7862,
  N7863,N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,N7873,N7874,N7875,
  N7876,N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889,
  N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,N7900,N7901,N7902,
  N7903,N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,N7913,N7914,N7915,
  N7916,N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,N7929,
  N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,N7939,N7940,N7941,N7942,
  N7943,N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,N7952,N7953,N7954,N7955,
  N7956,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,N7965,N7966,N7967,N7968,N7969,
  N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,N7979,N7980,N7981,N7982,
  N7983,N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,N7992,N7993,N7994,N7995,
  N7996,N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,N8005,N8006,N8007,N8008,N8009,
  N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,N8019,N8020,N8021,N8022,
  N8023,N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,N8032,N8033,N8034,N8035,
  N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,N8045,N8046,N8047,N8048,N8049,
  N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,N8059,N8060,N8061,N8062,
  N8063,N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,N8072,N8073,N8074,N8075,
  N8076,N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,N8085,N8086,N8087,N8088,N8089,
  N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,N8099,N8100,N8101,N8102,
  N8103,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,N8112,N8113,N8114,N8115,
  N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,N8125,N8126,N8127,N8128,N8129,
  N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,N8139,N8140,N8141,N8142,
  N8143,N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,N8152,N8153,N8154,N8155,
  N8156,N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,N8165,N8166,N8167,N8168,N8169,
  N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,N8179,N8180,N8181,N8182,
  N8183,N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,N8192,N8193,N8194,N8195,
  N8196,N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,N8205,N8206,N8207,N8208,N8209,
  N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,N8219,N8220,N8221,N8222,
  N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,N8232,N8233,N8234,N8235,
  N8236,N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,N8245,N8246,N8247,N8248,N8249,
  N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,N8259,N8260,N8261,N8262,
  N8263,N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,N8272,N8273,N8274,N8275,
  N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,N8285,N8286,N8287,N8288,N8289,
  N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,N8299,N8300,N8301,N8302,
  N8303,N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,N8312,N8313,N8314,N8315,
  N8316,N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324,N8325,N8326,N8327,N8328,N8329,
  N8330,N8331,N8332,N8333,N8334,N8335,N8336,N8337,N8338,N8339,N8340,N8341,N8342,
  N8343,N8344,N8345,N8346,N8347,N8348,N8349,N8350,N8351,N8352,N8353,N8354,N8355,
  N8356,N8357,N8358,N8359,N8360,N8361,N8362,N8363,N8364,N8365,N8366,N8367,N8368,N8369,
  N8370,N8371,N8372,N8373,N8374,N8375,N8376,N8377,N8378,N8379,N8380,N8381,N8382,
  N8383,N8384,N8385,N8386,N8387,N8388,N8389,N8390,N8391,N8392,N8393,N8394,N8395,
  N8396,N8397,N8398,N8399,N8400,N8401,N8402,N8403,N8404,N8405,N8406,N8407,N8408,N8409,
  N8410,N8411,N8412,N8413,N8414,N8415,N8416,N8417,N8418,N8419,N8420,N8421,N8422,
  N8423,N8424,N8425,N8426,N8427,N8428,N8429,N8430,N8431,N8432,N8433,N8434,N8435,
  N8436,N8437,N8438,N8439,N8440,N8441,N8442,N8443,N8444,N8445,N8446,N8447,N8448,N8449,
  N8450,N8451,N8452,N8453,N8454,N8455,N8456,N8457,N8458,N8459,N8460,N8461,N8462,
  N8463,N8464,N8465,N8466,N8467,N8468,N8469,N8470,N8471,N8472,N8473,N8474,N8475,
  N8476,N8477,N8478,N8479,N8480,N8481,N8482,N8483,N8484,N8485,N8486,N8487,N8488,N8489,
  N8490,N8491,N8492,N8493,N8494,N8495,N8496,N8497,N8498,N8499,N8500,N8501,N8502,
  N8503,N8504,N8505,N8506,N8507,N8508,N8509,N8510,N8511,N8512,N8513,N8514,N8515,
  N8516,N8517,N8518,N8519,N8520,N8521,N8522,N8523,N8524,N8525,N8526,N8527,N8528,N8529,
  N8530,N8531,N8532,N8533,N8534,N8535,N8536,N8537,N8538,N8539,N8540,N8541,N8542,
  N8543,N8544,N8545,N8546,N8547,N8548,N8549,N8550,N8551,N8552,N8553,N8554,N8555,
  N8556,N8557,N8558,N8559,N8560,N8561,N8562,N8563,N8564,N8565,N8566,N8567,N8568,N8569,
  N8570,N8571,N8572,N8573,N8574,N8575,N8576,N8577,N8578,N8579,N8580,N8581,N8582,
  N8583,N8584,N8585,N8586,N8587,N8588,N8589,N8590,N8591,N8592,N8593,N8594,N8595,
  N8596,N8597,N8598,N8599,N8600,N8601,N8602,N8603,N8604,N8605,N8606,N8607,N8608,N8609,
  N8610,N8611,N8612,N8613,N8614,N8615,N8616,N8617,N8618,N8619,N8620,N8621,N8622,
  N8623,N8624,N8625,N8626,N8627,N8628,N8629,N8630,N8631,N8632,N8633,N8634,N8635,
  N8636,N8637,N8638,N8639,N8640,N8641,N8642,N8643,N8644,N8645,N8646,N8647,N8648,N8649,
  N8650,N8651,N8652,N8653,N8654,N8655,N8656,N8657,N8658,N8659,N8660,N8661,N8662,
  N8663,N8664,N8665,N8666,N8667,N8668,N8669,N8670,N8671,N8672,N8673,N8674,N8675,
  N8676,N8677,N8678,N8679,N8680,N8681,N8682,N8683,N8684,N8685,N8686,N8687,N8688,N8689,
  N8690,N8691,N8692,N8693,N8694,N8695,N8696,N8697,N8698,N8699,N8700,N8701,N8702,
  N8703,N8704,N8705,N8706,N8707,N8708,N8709,N8710,N8711,N8712,N8713,N8714,N8715,
  N8716,N8717,N8718,N8719,N8720,N8721,N8722,N8723,N8724,N8725,N8726,N8727,N8728,N8729,
  N8730,N8731,N8732,N8733,N8734,N8735,N8736,N8737,N8738,N8739,N8740,N8741,N8742,
  N8743,N8744,N8745,N8746,N8747,N8748,N8749,N8750,N8751,N8752,N8753,N8754,N8755,
  N8756,N8757,N8758,N8759,N8760,N8761,N8762,N8763,N8764,N8765,N8766,N8767,N8768,N8769,
  N8770,N8771,N8772,N8773,N8774,N8775,N8776,N8777,N8778,N8779,N8780,N8781,N8782,
  N8783,N8784,N8785,N8786,N8787,N8788,N8789,N8790,N8791,N8792,N8793,N8794,N8795,
  N8796,N8797,N8798,N8799,N8800,N8801,N8802,N8803,N8804,N8805,N8806,N8807,N8808,N8809,
  N8810,N8811,N8812,N8813,N8814,N8815,N8816,N8817,N8818,N8819,N8820,N8821,N8822,
  N8823,N8824,N8825,N8826,N8827,N8828,N8829,N8830,N8831,N8832,N8833,N8834,N8835,
  N8836,N8837,N8838,N8839,N8840,N8841,N8842,N8843,N8844,N8845,N8846,N8847,N8848,N8849,
  N8850,N8851,N8852,N8853,N8854,N8855,N8856,N8857,N8858,N8859,N8860,N8861,N8862,
  N8863,N8864,N8865,N8866,N8867,N8868,N8869,N8870,N8871,N8872,N8873,N8874,N8875,
  N8876,N8877,N8878,N8879,N8880,N8881,N8882,N8883,N8884,N8885,N8886,N8887,N8888,N8889,
  N8890,N8891,N8892,N8893,N8894,N8895,N8896,N8897,N8898,N8899,N8900,N8901,N8902,
  N8903,N8904,N8905,N8906,N8907,N8908,N8909,N8910,N8911,N8912,N8913,N8914,N8915,
  N8916,N8917,N8918,N8919,N8920,N8921,N8922,N8923,N8924,N8925,N8926,N8927,N8928,N8929,
  N8930,N8931,N8932,N8933,N8934,N8935,N8936,N8937,N8938,N8939,N8940,N8941,N8942,
  N8943,N8944,N8945,N8946,N8947,N8948,N8949,N8950,N8951,N8952,N8953,N8954,N8955,
  N8956,N8957,N8958,N8959,N8960,N8961,N8962,N8963,N8964,N8965,N8966,N8967,N8968,N8969,
  N8970,N8971,N8972,N8973,N8974,N8975,N8976,N8977,N8978,N8979,N8980,N8981,N8982,
  N8983,N8984,N8985,N8986,N8987,N8988,N8989,N8990,N8991,N8992,N8993,N8994,N8995,
  N8996,N8997,N8998,N8999,N9000,N9001,N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009,
  N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017,N9018,N9019,N9020,N9021,N9022,
  N9023,N9024,N9025,N9026,N9027,N9028,N9029,N9030,N9031,N9032,N9033,N9034,N9035,
  N9036,N9037,N9038,N9039,N9040,N9041,N9042,N9043,N9044,N9045,N9046,N9047,N9048,N9049,
  N9050,N9051,N9052,N9053,N9054,N9055,N9056,N9057,N9058,N9059,N9060,N9061,N9062,
  N9063,N9064,N9065,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073,N9074,N9075,
  N9076,N9077,N9078,N9079,N9080,N9081,N9082,N9083,N9084,N9085,N9086,N9087,N9088,N9089,
  N9090,N9091,N9092,N9093,N9094,N9095,N9096,N9097,N9098,N9099,N9100,N9101,N9102,
  N9103,N9104,N9105,N9106,N9107,N9108,N9109,N9110,N9111,N9112,N9113,N9114,N9115,
  N9116,N9117,N9118,N9119,N9120,N9121,N9122,N9123,N9124,N9125,N9126,N9127,N9128,N9129,
  N9130,N9131,N9132,N9133,N9134,N9135,N9136,N9137,N9138,N9139,N9140,N9141,N9142,
  N9143,N9144,N9145,N9146,N9147,N9148,N9149,N9150,N9151,N9152,N9153,N9154,N9155,
  N9156,N9157,N9158,N9159,N9160,N9161,N9162,N9163,N9164,N9165,N9166,N9167,N9168,N9169,
  N9170,N9171,N9172,N9173,N9174,N9175,N9176,N9177,N9178,N9179,N9180,N9181,N9182,
  N9183,N9184,N9185,N9186,N9187,N9188,N9189,N9190,N9191,N9192,N9193,N9194,N9195,
  N9196,N9197,N9198,N9199,N9200,N9201,N9202,N9203,N9204,N9205,N9206,N9207,N9208,N9209,
  N9210,N9211,N9212,N9213,N9214,N9215,N9216,N9217,N9218,N9219,N9220,N9221,N9222,
  N9223,N9224,N9225,N9226,N9227,N9228,N9229,N9230,N9231,N9232,N9233,N9234,N9235,
  N9236,N9237,N9238,N9239,N9240,N9241,N9242,N9243,N9244,N9245,N9246,N9247,N9248,N9249,
  N9250,N9251,N9252,N9253,N9254,N9255,N9256,N9257,N9258,N9259,N9260,N9261,N9262,
  N9263,N9264,N9265,N9266,N9267,N9268,N9269,N9270,N9271,N9272,N9273,N9274,N9275,
  N9276,N9277,N9278,N9279,N9280,N9281,N9282,N9283,N9284,N9285,N9286,N9287,N9288,N9289,
  N9290,N9291,N9292,N9293,N9294,N9295,N9296,N9297,N9298,N9299,N9300,N9301,N9302,
  N9303,N9304,N9305,N9306,N9307,N9308,N9309,N9310,N9311,N9312,N9313,N9314,N9315,
  N9316,N9317,N9318,N9319,N9320,N9321,N9322,N9323,N9324,N9325,N9326,N9327,N9328,N9329,
  N9330,N9331,N9332,N9333,N9334,N9335,N9336,N9337,N9338,N9339,N9340,N9341,N9342,
  N9343,N9344,N9345,N9346,N9347,N9348,N9349,N9350,N9351,N9352,N9353,N9354,N9355,
  N9356,N9357,N9358,N9359,N9360,N9361,N9362,N9363,N9364,N9365,N9366,N9367,N9368,N9369,
  N9370,N9371,N9372,N9373,N9374,N9375,N9376,N9377,N9378,N9379,N9380,N9381,N9382,
  N9383,N9384,N9385,N9386,N9387,N9388,N9389,N9390,N9391,N9392,N9393,N9394,N9395,
  N9396,N9397,N9398,N9399,N9400,N9401,N9402,N9403,N9404,N9405,N9406,N9407,N9408,N9409,
  N9410,N9411,N9412,N9413,N9414,N9415,N9416,N9417,N9418,N9419,N9420,N9421,N9422,
  N9423,N9424,N9425,N9426,N9427,N9428,N9429,N9430,N9431,N9432,N9433,N9434,N9435,
  N9436,N9437,N9438,N9439,N9440,N9441,N9442,N9443,N9444,N9445,N9446,N9447,N9448,N9449,
  N9450,N9451,N9452,N9453,N9454,N9455,N9456,N9457,N9458,N9459,N9460,N9461,N9462,
  N9463,N9464,N9465,N9466,N9467,N9468,N9469,N9470,N9471,N9472,N9473,N9474,N9475,
  N9476,N9477,N9478,N9479,N9480,N9481,N9482,N9483,N9484,N9485,N9486,N9487,N9488,N9489,
  N9490,N9491,N9492,N9493,N9494,N9495,N9496,N9497,N9498,N9499,N9500,N9501,N9502,
  N9503,N9504,N9505,N9506,N9507,N9508,N9509,N9510,N9511,N9512,N9513,N9514,N9515,
  N9516,N9517,N9518,N9519,N9520,N9521,N9522,N9523,N9524,N9525,N9526,N9527,N9528,N9529,
  N9530,N9531,N9532,N9533,N9534,N9535,N9536,N9537,N9538,N9539,N9540,N9541,N9542,
  N9543,N9544,N9545,N9546,N9547,N9548,N9549,N9550,N9551,N9552,N9553,N9554,N9555,
  N9556,N9557,N9558,N9559,N9560,N9561,N9562,N9563,N9564,N9565,N9566,N9567,N9568,N9569,
  N9570,N9571,N9572,N9573,N9574,N9575,N9576,N9577,N9578,N9579,N9580,N9581,N9582,
  N9583,N9584,N9585,N9586,N9587,N9588,N9589,N9590,N9591,N9592,N9593,N9594,N9595,
  N9596,N9597,N9598,N9599,N9600,N9601,N9602,N9603,N9604,N9605,N9606,N9607,N9608,N9609,
  N9610,N9611,N9612,N9613,N9614,N9615,N9616,N9617,N9618,N9619,N9620,N9621,N9622,
  N9623,N9624,N9625,N9626,N9627,N9628,N9629,N9630,N9631,N9632,N9633,N9634,N9635,
  N9636,N9637,N9638,N9639,N9640,N9641,N9642,N9643,N9644,N9645,N9646,N9647,N9648,N9649,
  N9650,N9651,N9652,N9653,N9654,N9655,N9656,N9657,N9658,N9659,N9660,N9661,N9662,
  N9663,N9664,N9665,N9666,N9667,N9668,N9669,N9670,N9671,N9672,N9673,N9674,N9675,
  N9676,N9677,N9678,N9679,N9680,N9681,N9682,N9683,N9684,N9685,N9686,N9687,N9688,N9689,
  N9690,N9691,N9692,N9693,N9694,N9695,N9696,N9697,N9698,N9699,N9700,N9701,N9702,
  N9703,N9704,N9705,N9706,N9707,N9708,N9709,N9710,N9711,N9712,N9713,N9714,N9715,
  N9716,N9717,N9718,N9719,N9720,N9721,N9722,N9723,N9724,N9725,N9726,N9727,N9728,N9729,
  N9730,N9731,N9732,N9733,N9734,N9735,N9736,N9737,N9738,N9739,N9740,N9741,N9742,
  N9743,N9744,N9745,N9746,N9747,N9748,N9749,N9750,N9751,N9752,N9753,N9754,N9755,
  N9756,N9757,N9758,N9759,N9760,N9761,N9762,N9763,N9764,N9765,N9766,N9767,N9768,N9769,
  N9770,N9771,N9772,N9773,N9774,N9775,N9776,N9777,N9778,N9779,N9780,N9781,N9782,
  N9783,N9784,N9785,N9786,N9787,N9788,N9789,N9790,N9791,N9792,N9793,N9794,N9795,
  N9796,N9797,N9798,N9799,N9800,N9801,N9802,N9803,N9804,N9805,N9806,N9807,N9808,N9809,
  N9810,N9811,N9812,N9813,N9814,N9815,N9816,N9817,N9818,N9819,N9820,N9821,N9822,
  N9823,N9824,N9825,N9826,N9827,N9828,N9829,N9830,N9831,N9832,N9833,N9834,N9835,
  N9836,N9837,N9838,N9839,N9840,N9841,N9842,N9843,N9844,N9845,N9846,N9847,N9848,N9849,
  N9850,N9851,N9852,N9853,N9854,N9855,N9856,N9857,N9858,N9859,N9860,N9861,N9862,
  N9863,N9864,N9865,N9866,N9867,N9868,N9869,N9870,N9871,N9872,N9873,N9874,N9875,
  N9876,N9877,N9878,N9879,N9880,N9881,N9882,N9883,N9884,N9885,N9886,N9887,N9888,N9889,
  N9890,N9891,N9892,N9893,N9894,N9895,N9896,N9897,N9898,N9899,N9900,N9901,N9902,
  N9903,N9904,N9905,N9906,N9907,N9908,N9909,N9910,N9911,N9912,N9913,N9914,N9915,
  N9916,N9917,N9918,N9919,N9920,N9921,N9922,N9923,N9924,N9925,N9926,N9927,N9928,N9929,
  N9930,N9931,N9932,N9933,N9934,N9935,N9936,N9937,N9938,N9939,N9940,N9941,N9942,
  N9943,N9944,N9945,N9946,N9947,N9948,N9949,N9950,N9951,N9952,N9953,N9954,N9955,
  N9956,N9957,N9958,N9959,N9960,N9961,N9962,N9963,N9964,N9965,N9966,N9967,N9968,N9969,
  N9970,N9971,N9972,N9973,N9974,N9975,N9976,N9977,N9978,N9979,N9980,N9981,N9982,
  N9983,N9984,N9985,N9986,N9987,N9988,N9989,N9990,N9991,N9992,N9993,N9994,N9995,
  N9996,N9997,N9998,N9999,N10000,N10001,N10002,N10003,N10004,N10005,N10006,N10007,
  N10008,N10009,N10010,N10011,N10012,N10013,N10014,N10015,N10016,N10017,N10018,N10019,
  N10020,N10021,N10022,N10023,N10024,N10025,N10026,N10027,N10028,N10029,N10030,
  N10031,N10032,N10033,N10034,N10035,N10036,N10037,N10038,N10039,N10040,N10041,
  N10042,N10043,N10044,N10045,N10046,N10047,N10048,N10049,N10050,N10051,N10052,N10053,
  N10054,N10055,N10056,N10057,N10058,N10059,N10060,N10061,N10062,N10063,N10064,
  N10065,N10066,N10067,N10068,N10069,N10070,N10071,N10072,N10073,N10074,N10075,N10076,
  N10077,N10078,N10079,N10080,N10081,N10082,N10083,N10084,N10085,N10086,N10087,
  N10088,N10089,N10090,N10091,N10092,N10093,N10094,N10095,N10096,N10097,N10098,N10099,
  N10100,N10101,N10102,N10103,N10104,N10105,N10106,N10107,N10108,N10109,N10110,
  N10111,N10112,N10113,N10114,N10115,N10116,N10117,N10118,N10119,N10120,N10121,
  N10122,N10123,N10124,N10125,N10126,N10127,N10128,N10129,N10130,N10131,N10132,N10133,
  N10134,N10135,N10136,N10137,N10138,N10139,N10140,N10141,N10142,N10143,N10144,
  N10145,N10146,N10147,N10148,N10149,N10150,N10151,N10152,N10153,N10154,N10155,N10156,
  N10157,N10158,N10159,N10160,N10161,N10162,N10163,N10164,N10165,N10166,N10167,
  N10168,N10169,N10170,N10171,N10172,N10173,N10174,N10175,N10176,N10177,N10178,N10179,
  N10180,N10181,N10182,N10183,N10184,N10185,N10186,N10187,N10188,N10189,N10190,
  N10191,N10192,N10193,N10194,N10195,N10196,N10197,N10198,N10199,N10200,N10201,
  N10202,N10203,N10204,N10205,N10206,N10207,N10208,N10209,N10210,N10211,N10212,N10213,
  N10214,N10215,N10216,N10217,N10218,N10219,N10220,N10221,N10222,N10223,N10224,
  N10225,N10226,N10227,N10228,N10229,N10230,N10231,N10232,N10233,N10234,N10235,N10236,
  N10237,N10238,N10239,N10240,N10241,N10242,N10243,N10244,N10245,N10246,N10247,
  N10248,N10249,N10250,N10251,N10252,N10253,N10254,N10255,N10256,N10257,N10258,N10259,
  N10260,N10261,N10262,N10263,N10264,N10265,N10266,N10267,N10268,N10269,N10270,
  N10271,N10272,N10273,N10274,N10275,N10276,N10277,N10278,N10279,N10280,N10281,
  N10282,N10283,N10284,N10285,N10286,N10287,N10288,N10289,N10290,N10291,N10292,N10293,
  N10294,N10295,N10296,N10297,N10298,N10299,N10300,N10301,N10302,N10303,N10304,
  N10305,N10306,N10307,N10308,N10309,N10310,N10311,N10312,N10313,N10314,N10315,N10316,
  N10317,N10318,N10319,N10320,N10321,N10322,N10323,N10324,N10325,N10326,N10327,
  N10328,N10329,N10330,N10331,N10332,N10333,N10334,N10335,N10336,N10337,N10338,N10339,
  N10340,N10341,N10342,N10343,N10344,N10345,N10346,N10347,N10348,N10349,N10350,
  N10351,N10352,N10353,N10354,N10355,N10356,N10357,N10358,N10359,N10360,N10361,
  N10362,N10363,N10364,N10365,N10366,N10367,N10368,N10369,N10370,N10371,N10372,N10373,
  N10374,N10375,N10376,N10377,N10378,N10379,N10380,N10381,N10382,N10383,N10384,
  N10385,N10386,N10387,N10388,N10389,N10390,N10391,N10392,N10393,N10394,N10395,N10396,
  N10397,N10398,N10399,N10400,N10401,N10402,N10403,N10404,N10405,N10406,N10407,
  N10408,N10409,N10410,N10411,N10412,N10413,N10414,N10415,N10416,N10417,N10418,N10419,
  N10420,N10421,N10422,N10423,N10424,N10425,N10426,N10427,N10428,N10429,N10430,
  N10431,N10432,N10433,N10434,N10435,N10436,N10437,N10438,N10439,N10440,N10441,
  N10442,N10443,N10444,N10445,N10446,N10447,N10448,N10449,N10450,N10451,N10452,N10453,
  N10454,N10455,N10456,N10457,N10458,N10459,N10460,N10461,N10462,N10463,N10464,
  N10465,N10466,N10467,N10468,N10469,N10470,N10471,N10472,N10473,N10474,N10475,N10476,
  N10477,N10478,N10479,N10480,N10481,N10482,N10483,N10484,N10485,N10486,N10487,
  N10488,N10489,N10490,N10491,N10492,N10493,N10494,N10495,N10496,N10497,N10498,N10499,
  N10500,N10501,N10502,N10503,N10504,N10505,N10506,N10507,N10508,N10509,N10510,
  N10511,N10512,N10513,N10514,N10515,N10516,N10517,N10518,N10519,N10520,N10521,
  N10522,N10523,N10524,N10525,N10526,N10527,N10528,N10529,N10530,N10531,N10532,N10533,
  N10534,N10535,N10536,N10537,N10538,N10539,N10540,N10541,N10542,N10543,N10544,
  N10545,N10546,N10547,N10548,N10549,N10550,N10551,N10552,N10553,N10554,N10555,N10556,
  N10557,N10558,N10559,N10560,N10561,N10562,N10563,N10564,N10565,N10566,N10567,
  N10568,N10569,N10570,N10571,N10572,N10573,N10574,N10575,N10576,N10577,N10578,N10579,
  N10580,N10581,N10582,N10583,N10584,N10585,N10586,N10587,N10588,N10589,N10590,
  N10591,N10592,N10593,N10594,N10595,N10596,N10597,N10598,N10599,N10600,N10601,
  N10602,N10603,N10604,N10605,N10606,N10607,N10608,N10609,N10610,N10611,N10612,N10613,
  N10614,N10615,N10616,N10617,N10618,N10619,N10620,N10621,N10622,N10623,N10624,
  N10625,N10626,N10627,N10628,N10629,N10630,N10631,N10632,N10633,N10634,N10635,N10636,
  N10637,N10638,N10639,N10640,N10641,N10642,N10643,N10644,N10645,N10646,N10647,
  N10648,N10649,N10650,N10651,N10652,N10653,N10654,N10655,N10656,N10657,N10658,N10659,
  N10660,N10661,N10662,N10663,N10664,N10665,N10666,N10667,N10668,N10669,N10670,
  N10671,N10672,N10673,N10674,N10675,N10676,N10677,N10678,N10679,N10680,N10681,
  N10682,N10683,N10684,N10685,N10686,N10687,N10688,N10689,N10690,N10691,N10692,N10693,
  N10694,N10695,N10696,N10697,N10698,N10699,N10700,N10701,N10702,N10703,N10704,
  N10705,N10706,N10707,N10708,N10709,N10710,N10711,N10712,N10713,N10714,N10715,N10716,
  N10717,N10718,N10719,N10720,N10721,N10722,N10723,N10724,N10725,N10726,N10727,
  N10728,N10729,N10730,N10731,N10732,N10733,N10734,N10735,N10736,N10737,N10738,N10739,
  N10740,N10741,N10742,N10743,N10744,N10745,N10746,N10747,N10748,N10749,N10750,
  N10751,N10752,N10753,N10754,N10755,N10756,N10757,N10758,N10759,N10760,N10761,
  N10762,N10763,N10764,N10765,N10766,N10767,N10768,N10769,N10770,N10771,N10772,N10773,
  N10774,N10775,N10776,N10777,N10778,N10779,N10780,N10781,N10782,N10783,N10784,
  N10785,N10786,N10787,N10788,N10789,N10790,N10791,N10792,N10793,N10794,N10795,N10796,
  N10797,N10798,N10799,N10800,N10801,N10802,N10803,N10804,N10805,N10806,N10807,
  N10808,N10809,N10810,N10811,N10812,N10813,N10814,N10815,N10816,N10817,N10818,N10819,
  N10820,N10821,N10822,N10823,N10824,N10825,N10826,N10827,N10828,N10829,N10830,
  N10831,N10832,N10833,N10834,N10835,N10836,N10837,N10838,N10839,N10840,N10841,
  N10842,N10843,N10844,N10845,N10846,N10847,N10848,N10849,N10850,N10851,N10852,N10853,
  N10854,N10855,N10856,N10857,N10858,N10859,N10860,N10861,N10862,N10863,N10864,
  N10865,N10866,N10867,N10868,N10869,N10870,N10871,N10872,N10873,N10874,N10875,N10876,
  N10877,N10878,N10879,N10880,N10881,N10882,N10883,N10884,N10885,N10886,N10887,
  N10888,N10889,N10890,N10891,N10892,N10893,N10894,N10895,N10896,N10897,N10898,N10899,
  N10900,N10901,N10902,N10903,N10904,N10905,N10906,N10907,N10908,N10909,N10910,
  N10911,N10912,N10913,N10914,N10915,N10916,N10917,N10918,N10919,N10920,N10921,
  N10922,N10923,N10924,N10925,N10926,N10927,N10928,N10929,N10930,N10931,N10932,N10933,
  N10934,N10935,N10936,N10937,N10938,N10939,N10940,N10941,N10942,N10943,N10944,
  N10945,N10946,N10947,N10948,N10949,N10950,N10951,N10952,N10953,N10954,N10955,N10956,
  N10957,N10958,N10959,N10960,N10961,N10962,N10963,N10964,N10965,N10966,N10967,
  N10968,N10969,N10970,N10971,N10972,N10973,N10974,N10975,N10976,N10977,N10978,N10979,
  N10980,N10981,N10982,N10983,N10984,N10985,N10986,N10987,N10988,N10989,N10990,
  N10991,N10992,N10993,N10994,N10995,N10996,N10997,N10998,N10999,N11000,N11001,
  N11002,N11003,N11004,N11005,N11006,N11007,N11008,N11009,N11010,N11011,N11012,N11013,
  N11014,N11015,N11016,N11017,N11018,N11019,N11020,N11021,N11022,N11023,N11024,
  N11025,N11026,N11027,N11028,N11029,N11030,N11031,N11032,N11033,N11034,N11035,N11036,
  N11037,N11038,N11039,N11040,N11041,N11042,N11043,N11044,N11045,N11046,N11047,
  N11048,N11049,N11050,N11051,N11052,N11053,N11054,N11055,N11056,N11057,N11058,N11059,
  N11060,N11061,N11062,N11063,N11064,N11065,N11066,N11067,N11068,N11069,N11070,
  N11071,N11072,N11073,N11074,N11075,N11076,N11077,N11078,N11079,N11080,N11081,
  N11082,N11083,N11084,N11085,N11086,N11087,N11088,N11089,N11090,N11091,N11092,N11093,
  N11094,N11095,N11096,N11097,N11098,N11099,N11100,N11101,N11102,N11103,N11104,
  N11105,N11106,N11107,N11108,N11109,N11110,N11111,N11112,N11113,N11114,N11115,N11116,
  N11117,N11118,N11119,N11120,N11121,N11122,N11123,N11124,N11125,N11126,N11127,
  N11128,N11129,N11130,N11131,N11132,N11133,N11134,N11135,N11136,N11137,N11138,N11139,
  N11140,N11141,N11142,N11143,N11144,N11145,N11146,N11147,N11148,N11149,N11150,
  N11151,N11152,N11153,N11154,N11155,N11156,N11157,N11158,N11159,N11160,N11161,
  N11162,N11163,N11164,N11165,N11166,N11167,N11168,N11169,N11170,N11171,N11172,N11173,
  N11174,N11175,N11176,N11177,N11178,N11179,N11180,N11181,N11182,N11183,N11184,
  N11185,N11186,N11187,N11188,N11189,N11190,N11191,N11192,N11193,N11194,N11195,N11196,
  N11197,N11198,N11199,N11200,N11201,N11202,N11203,N11204,N11205,N11206,N11207,
  N11208,N11209,N11210,N11211,N11212,N11213,N11214,N11215,N11216,N11217,N11218,N11219,
  N11220,N11221,N11222,N11223,N11224,N11225,N11226,N11227,N11228,N11229,N11230,
  N11231,N11232,N11233,N11234,N11235,N11236,N11237,N11238,N11239,N11240,N11241,
  N11242,N11243,N11244,N11245,N11246,N11247,N11248,N11249,N11250,N11251,N11252,N11253,
  N11254,N11255,N11256,N11257,N11258,N11259,N11260,N11261,N11262,N11263,N11264,
  N11265,N11266,N11267,N11268,N11269,N11270,N11271,N11272,N11273,N11274,N11275,N11276,
  N11277,N11278,N11279,N11280,N11281,N11282,N11283,N11284,N11285,N11286,N11287,
  N11288,N11289,N11290,N11291,N11292,N11293,N11294,N11295,N11296,N11297,N11298,N11299,
  N11300,N11301,N11302,N11303,N11304,N11305,N11306,N11307,N11308,N11309,N11310,
  N11311,N11312,N11313,N11314,N11315,N11316,N11317,N11318,N11319,N11320,N11321,
  N11322,N11323,N11324,N11325,N11326,N11327,N11328,N11329,N11330,N11331,N11332,N11333,
  N11334,N11335,N11336,N11337,N11338,N11339,N11340,N11341,N11342,N11343,N11344,
  N11345,N11346,N11347,N11348,N11349,N11350,N11351,N11352,N11353,N11354,N11355,N11356,
  N11357,N11358,N11359,N11360,N11361,N11362,N11363,N11364,N11365,N11366,N11367,
  N11368,N11369,N11370,N11371,N11372,N11373,N11374,N11375,N11376,N11377,N11378,N11379,
  N11380,N11381,N11382,N11383,N11384,N11385,N11386,N11387,N11388,N11389,N11390,
  N11391,N11392,N11393,N11394,N11395,N11396,N11397,N11398,N11399,N11400,N11401,
  N11402,N11403,N11404,N11405,N11406,N11407,N11408,N11409,N11410,N11411,N11412,N11413,
  N11414,N11415,N11416,N11417,N11418,N11419,N11420,N11421,N11422,N11423,N11424,
  N11425,N11426,N11427,N11428,N11429,N11430,N11431,N11432,N11433,N11434,N11435,N11436,
  N11437,N11438,N11439,N11440,N11441,N11442,N11443,N11444,N11445,N11446,N11447,
  N11448,N11449,N11450,N11451,N11452,N11453,N11454,N11455,N11456,N11457,N11458,N11459,
  N11460,N11461,N11462,N11463,N11464,N11465,N11466,N11467,N11468,N11469,N11470,
  N11471,N11472,N11473,N11474,N11475,N11476,N11477,N11478,N11479,N11480,N11481,
  N11482,N11483,N11484,N11485,N11486,N11487,N11488,N11489,N11490,N11491,N11492,N11493,
  N11494,N11495,N11496,N11497,N11498,N11499,N11500,N11501,N11502,N11503,N11504,
  N11505,N11506,N11507,N11508,N11509,N11510,N11511,N11512,N11513,N11514,N11515,N11516,
  N11517,N11518,N11519,N11520,N11521,N11522,N11523,N11524,N11525,N11526,N11527,
  N11528,N11529,N11530,N11531,N11532,N11533,N11534,N11535,N11536,N11537,N11538,N11539,
  N11540,N11541,N11542,N11543,N11544,N11545,N11546,N11547,N11548,N11549,N11550,
  N11551,N11552,N11553,N11554,N11555,N11556,N11557,N11558,N11559,N11560,N11561,
  N11562,N11563,N11564,N11565,N11566,N11567,N11568,N11569,N11570,N11571,N11572,N11573,
  N11574,N11575,N11576,N11577,N11578,N11579,N11580,N11581,N11582,N11583,N11584,
  N11585,N11586,N11587,N11588,N11589,N11590,N11591,N11592,N11593,N11594,N11595,N11596,
  N11597,N11598,N11599,N11600,N11601,N11602,N11603,N11604,N11605,N11606,N11607,
  N11608,N11609,N11610,N11611,N11612,N11613,N11614,N11615,N11616,N11617,N11618,N11619,
  N11620,N11621,N11622,N11623,N11624,N11625,N11626,N11627,N11628,N11629,N11630,
  N11631,N11632,N11633,N11634,N11635,N11636,N11637,N11638,N11639,N11640,N11641,
  N11642,N11643,N11644,N11645,N11646,N11647,N11648,N11649,N11650,N11651,N11652,N11653,
  N11654,N11655,N11656,N11657,N11658,N11659,N11660,N11661,N11662,N11663,N11664,
  N11665,N11666,N11667,N11668,N11669,N11670,N11671,N11672,N11673,N11674,N11675,N11676,
  N11677,N11678,N11679,N11680,N11681,N11682,N11683,N11684,N11685,N11686,N11687,
  N11688,N11689,N11690,N11691,N11692,N11693,N11694,N11695,N11696,N11697,N11698,N11699,
  N11700,N11701,N11702,N11703,N11704,N11705,N11706,N11707,N11708,N11709,N11710,
  N11711,N11712,N11713,N11714,N11715,N11716,N11717,N11718,N11719,N11720,N11721,
  N11722,N11723,N11724,N11725,N11726,N11727,N11728,N11729,N11730,N11731,N11732,N11733,
  N11734,N11735,N11736,N11737,N11738,N11739,N11740,N11741,N11742,N11743,N11744,
  N11745,N11746,N11747,N11748,N11749,N11750,N11751,N11752,N11753,N11754,N11755,N11756,
  N11757,N11758,N11759,N11760,N11761,N11762,N11763,N11764,N11765,N11766,N11767,
  N11768,N11769,N11770,N11771,N11772,N11773,N11774,N11775,N11776,N11777,N11778,N11779,
  N11780,N11781,N11782,N11783,N11784,N11785,N11786,N11787,N11788,N11789,N11790,
  N11791,N11792,N11793,N11794,N11795,N11796,N11797,N11798,N11799,N11800,N11801,
  N11802,N11803,N11804,N11805,N11806,N11807,N11808,N11809,N11810,N11811,N11812,N11813,
  N11814,N11815,N11816,N11817,N11818,N11819,N11820,N11821,N11822,N11823,N11824,
  N11825,N11826,N11827,N11828,N11829,N11830,N11831,N11832,N11833,N11834,N11835,N11836,
  N11837,N11838,N11839,N11840,N11841,N11842,N11843,N11844,N11845,N11846,N11847,
  N11848,N11849,N11850,N11851,N11852,N11853,N11854,N11855,N11856,N11857,N11858,N11859,
  N11860,N11861,N11862,N11863,N11864,N11865,N11866,N11867,N11868,N11869,N11870,
  N11871,N11872,N11873,N11874,N11875,N11876,N11877,N11878,N11879,N11880,N11881,
  N11882,N11883,N11884,N11885,N11886,N11887,N11888,N11889,N11890,N11891,N11892,N11893,
  N11894,N11895,N11896,N11897,N11898,N11899,N11900,N11901,N11902,N11903,N11904,
  N11905,N11906,N11907,N11908,N11909,N11910,N11911,N11912,N11913,N11914,N11915,N11916,
  N11917,N11918,N11919,N11920,N11921,N11922,N11923,N11924,N11925,N11926,N11927,
  N11928,N11929,N11930,N11931,N11932,N11933,N11934,N11935,N11936,N11937,N11938,N11939,
  N11940,N11941,N11942,N11943,N11944,N11945,N11946,N11947,N11948,N11949,N11950,
  N11951,N11952,N11953,N11954,N11955,N11956,N11957,N11958,N11959,N11960,N11961,
  N11962,N11963,N11964,N11965,N11966,N11967,N11968,N11969,N11970,N11971,N11972,N11973,
  N11974,N11975,N11976,N11977,N11978,N11979,N11980,N11981,N11982,N11983,N11984,
  N11985,N11986,N11987,N11988,N11989,N11990,N11991,N11992,N11993,N11994,N11995,N11996,
  N11997,N11998,N11999,N12000,N12001,N12002,N12003,N12004,N12005,N12006,N12007,
  N12008,N12009,N12010,N12011,N12012,N12013,N12014,N12015,N12016,N12017,N12018,N12019,
  N12020,N12021,N12022,N12023,N12024,N12025,N12026,N12027,N12028,N12029,N12030,
  N12031,N12032,N12033,N12034,N12035,N12036,N12037,N12038,N12039,N12040,N12041,
  N12042,N12043,N12044,N12045,N12046,N12047,N12048,N12049,N12050,N12051,N12052,N12053,
  N12054,N12055,N12056,N12057,N12058,N12059,N12060,N12061,N12062,N12063,N12064,
  N12065,N12066,N12067,N12068,N12069,N12070,N12071,N12072,N12073,N12074,N12075,N12076,
  N12077,N12078,N12079,N12080,N12081,N12082,N12083,N12084,N12085,N12086,N12087,
  N12088,N12089,N12090,N12091,N12092,N12093,N12094,N12095,N12096,N12097,N12098,N12099,
  N12100,N12101,N12102,N12103,N12104,N12105,N12106,N12107,N12108,N12109,N12110,
  N12111,N12112,N12113,N12114,N12115,N12116,N12117,N12118,N12119,N12120,N12121,
  N12122,N12123,N12124,N12125,N12126,N12127,N12128,N12129,N12130,N12131,N12132,N12133,
  N12134,N12135,N12136,N12137,N12138,N12139,N12140,N12141,N12142,N12143,N12144,
  N12145,N12146,N12147,N12148,N12149,N12150,N12151,N12152,N12153,N12154,N12155,N12156,
  N12157,N12158,N12159,N12160,N12161,N12162,N12163,N12164,N12165,N12166,N12167,
  N12168,N12169,N12170,N12171,N12172,N12173,N12174,N12175,N12176,N12177,N12178,N12179,
  N12180,N12181,N12182,N12183,N12184,N12185,N12186,N12187,N12188,N12189,N12190,
  N12191,N12192,N12193,N12194,N12195,N12196,N12197,N12198,N12199,N12200,N12201,
  N12202,N12203,N12204,N12205,N12206,N12207,N12208,N12209,N12210,N12211,N12212,N12213,
  N12214,N12215,N12216,N12217,N12218,N12219,N12220,N12221,N12222,N12223,N12224,
  N12225,N12226,N12227,N12228,N12229,N12230,N12231,N12232,N12233,N12234,N12235,N12236,
  N12237,N12238,N12239,N12240,N12241,N12242,N12243,N12244,N12245,N12246,N12247,
  N12248,N12249,N12250,N12251,N12252,N12253,N12254,N12255,N12256,N12257,N12258,N12259,
  N12260,N12261,N12262,N12263,N12264,N12265,N12266,N12267,N12268,N12269,N12270,
  N12271,N12272,N12273,N12274,N12275,N12276,N12277,N12278,N12279,N12280,N12281,
  N12282,N12283,N12284,N12285,N12286,N12287,N12288,N12289,N12290,N12291,N12292,N12293,
  N12294,N12295,N12296,N12297,N12298,N12299,N12300,N12301,N12302,N12303,N12304,
  N12305,N12306,N12307,N12308,N12309,N12310,N12311,N12312,N12313,N12314,N12315,N12316,
  N12317,N12318,N12319,N12320,N12321,N12322,N12323,N12324,N12325,N12326,N12327,
  N12328,N12329,N12330,N12331,N12332,N12333,N12334,N12335,N12336,N12337,N12338,N12339,
  N12340,N12341,N12342,N12343,N12344,N12345,N12346,N12347,N12348,N12349,N12350,
  N12351,N12352,N12353,N12354,N12355,N12356,N12357,N12358,N12359,N12360,N12361,
  N12362,N12363,N12364,N12365,N12366,N12367,N12368,N12369,N12370,N12371,N12372,N12373,
  N12374,N12375,N12376,N12377,N12378,N12379,N12380,N12381,N12382,N12383,N12384,
  N12385,N12386,N12387,N12388,N12389,N12390,N12391,N12392,N12393,N12394,N12395,N12396,
  N12397,N12398,N12399,N12400,N12401,N12402,N12403,N12404,N12405,N12406,N12407,
  N12408,N12409,N12410,N12411,N12412,N12413,N12414,N12415,N12416,N12417,N12418,N12419,
  N12420,N12421,N12422,N12423,N12424,N12425,N12426,N12427,N12428,N12429,N12430,
  N12431,N12432,N12433,N12434,N12435,N12436,N12437,N12438,N12439,N12440,N12441,
  N12442,N12443,N12444,N12445,N12446,N12447,N12448,N12449,N12450,N12451,N12452,N12453,
  N12454,N12455,N12456,N12457,N12458,N12459,N12460,N12461,N12462,N12463,N12464,
  N12465,N12466,N12467,N12468,N12469,N12470,N12471,N12472,N12473,N12474,N12475,N12476,
  N12477,N12478,N12479,N12480,N12481,N12482,N12483,N12484,N12485,N12486,N12487,
  N12488,N12489,N12490,N12491,N12492,N12493,N12494,N12495,N12496,N12497,N12498,N12499,
  N12500,N12501,N12502,N12503,N12504,N12505,N12506,N12507,N12508,N12509,N12510,
  N12511,N12512,N12513,N12514,N12515,N12516,N12517,N12518,N12519,N12520,N12521,
  N12522,N12523,N12524,N12525,N12526,N12527,N12528,N12529,N12530,N12531,N12532,N12533,
  N12534,N12535,N12536,N12537,N12538,N12539,N12540,N12541,N12542,N12543,N12544,
  N12545,N12546,N12547,N12548,N12549,N12550,N12551,N12552,N12553,N12554,N12555,N12556,
  N12557,N12558,N12559,N12560,N12561,N12562,N12563,N12564,N12565,N12566,N12567,
  N12568,N12569,N12570,N12571,N12572,N12573,N12574,N12575,N12576,N12577,N12578,N12579,
  N12580,N12581,N12582,N12583,N12584,N12585,N12586,N12587,N12588,N12589,N12590,
  N12591,N12592,N12593,N12594,N12595,N12596,N12597,N12598,N12599,N12600,N12601,
  N12602,N12603,N12604,N12605,N12606,N12607,N12608,N12609,N12610,N12611,N12612,N12613,
  N12614,N12615,N12616,N12617,N12618,N12619,N12620,N12621,N12622,N12623,N12624,
  N12625,N12626,N12627,N12628,N12629,N12630,N12631,N12632,N12633,N12634,N12635,N12636,
  N12637,N12638,N12639,N12640,N12641,N12642,N12643,N12644,N12645,N12646,N12647,
  N12648,N12649,N12650,N12651,N12652,N12653,N12654,N12655,N12656,N12657,N12658,N12659,
  N12660,N12661,N12662,N12663,N12664,N12665,N12666,N12667,N12668,N12669,N12670,
  N12671,N12672,N12673,N12674,N12675,N12676,N12677,N12678,N12679,N12680,N12681,
  N12682,N12683,N12684,N12685,N12686,N12687,N12688,N12689,N12690,N12691,N12692,N12693,
  N12694,N12695,N12696,N12697,N12698,N12699,N12700,N12701,N12702,N12703,N12704,
  N12705,N12706,N12707,N12708,N12709,N12710,N12711,N12712,N12713,N12714,N12715,N12716,
  N12717,N12718,N12719,N12720,N12721,N12722,N12723,N12724,N12725,N12726,N12727,
  N12728,N12729,N12730,N12731,N12732,N12733,N12734,N12735,N12736,N12737,N12738,N12739,
  N12740,N12741,N12742,N12743,N12744,N12745,N12746,N12747,N12748,N12749,N12750,
  N12751,N12752,N12753,N12754,N12755,N12756,N12757,N12758,N12759,N12760,N12761,
  N12762,N12763,N12764,N12765,N12766,N12767,N12768,N12769,N12770,N12771,N12772,N12773,
  N12774,N12775,N12776,N12777,N12778,N12779,N12780,N12781,N12782,N12783,N12784,
  N12785,N12786,N12787,N12788,N12789,N12790,N12791,N12792,N12793,N12794,N12795,N12796,
  N12797,N12798,N12799,N12800,N12801,N12802,N12803,N12804,N12805,N12806,N12807,
  N12808,N12809,N12810,N12811,N12812,N12813,N12814,N12815,N12816,N12817,N12818,N12819,
  N12820,N12821,N12822,N12823,N12824,N12825,N12826,N12827,N12828,N12829,N12830,
  N12831,N12832,N12833,N12834,N12835,N12836,N12837,N12838,N12839,N12840,N12841,
  N12842,N12843,N12844,N12845,N12846,N12847,N12848,N12849,N12850,N12851,N12852,N12853,
  N12854,N12855,N12856,N12857,N12858,N12859,N12860,N12861,N12862,N12863,N12864,
  N12865,N12866,N12867,N12868,N12869,N12870,N12871,N12872,N12873,N12874,N12875,N12876,
  N12877,N12878,N12879,N12880,N12881,N12882,N12883,N12884,N12885,N12886,N12887,
  N12888,N12889,N12890,N12891,N12892,N12893,N12894,N12895,N12896,N12897,N12898,N12899,
  N12900,N12901,N12902,N12903,N12904,N12905,N12906,N12907,N12908,N12909,N12910,
  N12911,N12912,N12913,N12914,N12915,N12916,N12917,N12918,N12919,N12920,N12921,
  N12922,N12923,N12924,N12925,N12926,N12927,N12928,N12929,N12930,N12931,N12932,N12933,
  N12934,N12935,N12936,N12937,N12938,N12939,N12940,N12941,N12942,N12943,N12944,
  N12945,N12946,N12947,N12948,N12949,N12950,N12951,N12952,N12953,N12954,N12955,N12956,
  N12957,N12958,N12959,N12960,N12961,N12962,N12963,N12964,N12965,N12966,N12967,
  N12968,N12969,N12970,N12971,N12972,N12973,N12974,N12975,N12976,N12977,N12978,N12979,
  N12980,N12981,N12982,N12983,N12984,N12985,N12986,N12987,N12988,N12989,N12990,
  N12991,N12992,N12993,N12994,N12995,N12996,N12997,N12998,N12999,N13000,N13001,
  N13002,N13003,N13004,N13005,N13006,N13007,N13008,N13009,N13010,N13011,N13012,N13013,
  N13014,N13015,N13016,N13017,N13018,N13019,N13020,N13021,N13022,N13023,N13024,
  N13025,N13026,N13027,N13028,N13029,N13030,N13031,N13032,N13033,N13034,N13035,N13036,
  N13037,N13038,N13039,N13040,N13041,N13042,N13043,N13044,N13045,N13046,N13047,
  N13048,N13049,N13050,N13051,N13052,N13053,N13054,N13055,N13056,N13057,N13058,N13059,
  N13060,N13061,N13062,N13063,N13064,N13065,N13066,N13067,N13068,N13069,N13070,
  N13071,N13072,N13073,N13074,N13075,N13076,N13077,N13078,N13079,N13080,N13081,
  N13082,N13083,N13084,N13085,N13086,N13087,N13088,N13089,N13090,N13091,N13092,N13093,
  N13094,N13095,N13096,N13097,N13098,N13099,N13100,N13101,N13102,N13103,N13104,
  N13105,N13106,N13107,N13108,N13109,N13110,N13111,N13112,N13113,N13114,N13115,N13116,
  N13117,N13118,N13119,N13120,N13121,N13122,N13123,N13124,N13125,N13126,N13127,
  N13128,N13129,N13130,N13131,N13132,N13133,N13134,N13135,N13136,N13137,N13138,N13139,
  N13140,N13141,N13142,N13143,N13144,N13145,N13146,N13147,N13148,N13149,N13150,
  N13151,N13152,N13153,N13154,N13155,N13156,N13157,N13158,N13159,N13160,N13161,
  N13162,N13163,N13164,N13165,N13166,N13167,N13168,N13169,N13170,N13171,N13172,N13173,
  N13174,N13175,N13176,N13177,N13178,N13179,N13180,N13181,N13182,N13183,N13184,
  N13185,N13186,N13187,N13188,N13189,N13190,N13191,N13192,N13193,N13194,N13195,N13196,
  N13197,N13198,N13199,N13200,N13201,N13202,N13203,N13204,N13205,N13206,N13207,
  N13208,N13209,N13210,N13211,N13212,N13213,N13214,N13215,N13216,N13217,N13218,N13219,
  N13220,N13221,N13222,N13223,N13224,N13225,N13226,N13227,N13228,N13229,N13230,
  N13231,N13232,N13233,N13234,N13235,N13236,N13237,N13238,N13239,N13240,N13241,
  N13242,N13243,N13244,N13245,N13246,N13247,N13248,N13249,N13250,N13251,N13252,N13253,
  N13254,N13255,N13256,N13257,N13258,N13259,N13260,N13261,N13262,N13263,N13264,
  N13265,N13266,N13267,N13268,N13269,N13270,N13271,N13272,N13273,N13274,N13275,N13276,
  N13277,N13278,N13279,N13280,N13281,N13282,N13283,N13284,N13285,N13286,N13287,
  N13288,N13289,N13290,N13291,N13292,N13293,N13294,N13295,N13296,N13297,N13298,N13299,
  N13300,N13301,N13302,N13303,N13304,N13305,N13306,N13307,N13308,N13309,N13310,
  N13311,N13312,N13313,N13314,N13315,N13316,N13317,N13318,N13319,N13320,N13321,
  N13322,N13323,N13324,N13325,N13326,N13327,N13328,N13329,N13330,N13331,N13332,N13333,
  N13334,N13335,N13336,N13337,N13338,N13339,N13340,N13341,N13342,N13343,N13344,
  N13345,N13346,N13347,N13348,N13349,N13350,N13351,N13352,N13353,N13354,N13355,N13356,
  N13357,N13358,N13359,N13360,N13361,N13362,N13363,N13364,N13365,N13366,N13367,
  N13368,N13369,N13370,N13371,N13372,N13373,N13374,N13375,N13376,N13377,N13378,N13379,
  N13380,N13381,N13382,N13383,N13384,N13385,N13386,N13387,N13388,N13389,N13390,
  N13391,N13392,N13393,N13394,N13395,N13396,N13397,N13398,N13399,N13400,N13401,
  N13402,N13403,N13404,N13405,N13406,N13407,N13408,N13409,N13410,N13411,N13412,N13413,
  N13414,N13415,N13416,N13417,N13418,N13419,N13420,N13421,N13422,N13423,N13424,
  N13425,N13426,N13427,N13428,N13429,N13430,N13431,N13432,N13433,N13434,N13435,N13436,
  N13437,N13438,N13439,N13440,N13441,N13442,N13443,N13444,N13445,N13446,N13447,
  N13448,N13449,N13450,N13451,N13452,N13453,N13454,N13455,N13456,N13457,N13458,N13459,
  N13460,N13461,N13462,N13463,N13464,N13465,N13466,N13467,N13468,N13469,N13470,
  N13471,N13472,N13473,N13474,N13475,N13476,N13477,N13478,N13479,N13480,N13481,
  N13482,N13483,N13484,N13485,N13486,N13487,N13488,N13489,N13490,N13491,N13492,N13493,
  N13494,N13495,N13496,N13497,N13498,N13499,N13500,N13501,N13502,N13503,N13504,
  N13505,N13506,N13507,N13508,N13509,N13510,N13511,N13512,N13513,N13514,N13515,N13516,
  N13517,N13518,N13519,N13520,N13521,N13522,N13523,N13524,N13525,N13526,N13527,
  N13528,N13529,N13530,N13531,N13532,N13533,N13534,N13535,N13536,N13537,N13538,N13539,
  N13540,N13541,N13542,N13543,N13544,N13545,N13546,N13547,N13548,N13549,N13550,
  N13551,N13552,N13553,N13554,N13555,N13556,N13557,N13558,N13559,N13560,N13561,
  N13562,N13563,N13564,N13565,N13566,N13567,N13568,N13569,N13570,N13571,N13572,N13573,
  N13574,N13575,N13576,N13577,N13578,N13579,N13580,N13581,N13582,N13583,N13584,
  N13585,N13586,N13587,N13588,N13589,N13590,N13591,N13592,N13593,N13594,N13595,N13596,
  N13597,N13598,N13599,N13600,N13601,N13602,N13603,N13604,N13605,N13606,N13607,
  N13608,N13609,N13610,N13611,N13612,N13613,N13614,N13615,N13616,N13617,N13618,N13619,
  N13620,N13621,N13622,N13623,N13624,N13625,N13626,N13627,N13628,N13629,N13630,
  N13631,N13632,N13633,N13634,N13635,N13636,N13637,N13638,N13639,N13640,N13641,
  N13642,N13643,N13644,N13645,N13646,N13647,N13648,N13649,N13650,N13651,N13652,N13653,
  N13654,N13655,N13656,N13657,N13658,N13659,N13660,N13661,N13662,N13663,N13664,
  N13665,N13666,N13667,N13668,N13669,N13670,N13671,N13672,N13673,N13674,N13675,N13676,
  N13677,N13678,N13679,N13680,N13681,N13682,N13683,N13684,N13685,N13686,N13687,
  N13688,N13689,N13690,N13691,N13692,N13693,N13694,N13695,N13696,N13697,N13698,N13699,
  N13700,N13701,N13702,N13703,N13704,N13705,N13706,N13707,N13708,N13709,N13710,
  N13711,N13712,N13713,N13714,N13715,N13716,N13717,N13718,N13719,N13720,N13721,
  N13722,N13723,N13724,N13725,N13726,N13727,N13728,N13729,N13730,N13731,N13732,N13733,
  N13734,N13735,N13736,N13737,N13738,N13739,N13740,N13741,N13742,N13743,N13744,
  N13745,N13746,N13747,N13748,N13749,N13750,N13751,N13752,N13753,N13754,N13755,N13756,
  N13757,N13758,N13759,N13760,N13761,N13762,N13763,N13764,N13765,N13766,N13767,
  N13768,N13769,N13770,N13771,N13772,N13773,N13774,N13775,N13776,N13777,N13778,N13779,
  N13780,N13781,N13782,N13783,N13784,N13785,N13786,N13787,N13788,N13789,N13790,
  N13791,N13792,N13793,N13794,N13795,N13796,N13797,N13798,N13799,N13800,N13801,
  N13802,N13803,N13804,N13805,N13806,N13807,N13808,N13809,N13810,N13811,N13812,N13813,
  N13814,N13815,N13816,N13817,N13818,N13819,N13820,N13821,N13822,N13823,N13824,
  N13825,N13826,N13827,N13828,N13829,N13830,N13831,N13832,N13833,N13834,N13835,N13836,
  N13837,N13838,N13839,N13840,N13841,N13842,N13843,N13844,N13845,N13846,N13847,
  N13848,N13849,N13850,N13851,N13852,N13853,N13854,N13855,N13856,N13857,N13858,N13859,
  N13860,N13861,N13862,N13863,N13864,N13865,N13866,N13867,N13868,N13869,N13870,
  N13871,N13872,N13873,N13874,N13875,N13876,N13877,N13878,N13879,N13880,N13881,
  N13882,N13883,N13884,N13885,N13886,N13887,N13888,N13889,N13890,N13891,N13892,N13893,
  N13894,N13895,N13896,N13897,N13898,N13899,N13900,N13901,N13902,N13903,N13904,
  N13905,N13906,N13907,N13908,N13909,N13910,N13911,N13912,N13913,N13914,N13915,N13916,
  N13917,N13918,N13919,N13920,N13921,N13922,N13923,N13924,N13925,N13926,N13927,
  N13928,N13929,N13930,N13931,N13932,N13933,N13934,N13935,N13936,N13937,N13938,N13939,
  N13940,N13941,N13942,N13943,N13944,N13945,N13946,N13947,N13948,N13949,N13950,
  N13951,N13952,N13953,N13954,N13955,N13956,N13957,N13958,N13959,N13960,N13961,
  N13962,N13963,N13964,N13965,N13966,N13967,N13968,N13969,N13970,N13971,N13972,N13973,
  N13974,N13975,N13976,N13977,N13978,N13979,N13980,N13981,N13982,N13983,N13984,
  N13985,N13986,N13987,N13988,N13989,N13990,N13991,N13992,N13993,N13994,N13995,N13996,
  N13997,N13998,N13999,N14000,N14001,N14002,N14003,N14004,N14005,N14006,N14007,
  N14008,N14009,N14010,N14011,N14012,N14013,N14014,N14015,N14016,N14017,N14018,N14019,
  N14020,N14021,N14022,N14023,N14024,N14025,N14026,N14027,N14028,N14029,N14030,
  N14031,N14032,N14033,N14034,N14035,N14036,N14037,N14038,N14039,N14040,N14041,
  N14042,N14043,N14044,N14045,N14046,N14047,N14048,N14049,N14050,N14051,N14052,N14053,
  N14054,N14055,N14056,N14057,N14058,N14059,N14060,N14061,N14062,N14063,N14064,
  N14065,N14066,N14067,N14068,N14069,N14070,N14071,N14072,N14073,N14074,N14075,N14076,
  N14077,N14078,N14079,N14080,N14081,N14082,N14083,N14084,N14085,N14086,N14087,
  N14088,N14089,N14090,N14091,N14092,N14093,N14094,N14095,N14096,N14097,N14098,N14099,
  N14100,N14101,N14102,N14103,N14104,N14105,N14106,N14107,N14108,N14109,N14110,
  N14111,N14112,N14113,N14114,N14115,N14116,N14117,N14118,N14119,N14120,N14121,
  N14122,N14123,N14124,N14125,N14126,N14127,N14128,N14129,N14130,N14131,N14132,N14133,
  N14134,N14135,N14136,N14137,N14138,N14139,N14140,N14141,N14142,N14143,N14144,
  N14145,N14146,N14147,N14148,N14149,N14150,N14151,N14152,N14153,N14154,N14155,N14156,
  N14157,N14158,N14159,N14160,N14161,N14162,N14163,N14164,N14165,N14166,N14167,
  N14168,N14169,N14170,N14171,N14172,N14173,N14174,N14175,N14176,N14177,N14178,N14179,
  N14180,N14181,N14182,N14183,N14184,N14185,N14186,N14187,N14188,N14189,N14190,
  N14191,N14192,N14193,N14194,N14195,N14196,N14197,N14198,N14199,N14200,N14201,
  N14202,N14203,N14204,N14205,N14206,N14207,N14208,N14209,N14210,N14211,N14212,N14213,
  N14214,N14215,N14216,N14217,N14218,N14219,N14220,N14221,N14222,N14223,N14224,
  N14225,N14226,N14227,N14228,N14229,N14230,N14231,N14232,N14233,N14234,N14235,N14236,
  N14237,N14238,N14239,N14240,N14241,N14242,N14243,N14244,N14245,N14246,N14247,
  N14248,N14249,N14250,N14251,N14252,N14253,N14254,N14255,N14256,N14257,N14258,N14259,
  N14260,N14261,N14262,N14263,N14264,N14265,N14266,N14267,N14268,N14269,N14270,
  N14271,N14272,N14273,N14274,N14275,N14276,N14277,N14278,N14279,N14280,N14281,
  N14282,N14283,N14284,N14285,N14286,N14287,N14288,N14289,N14290,N14291,N14292,N14293,
  N14294,N14295,N14296,N14297,N14298,N14299,N14300,N14301,N14302,N14303,N14304,
  N14305,N14306,N14307,N14308,N14309,N14310,N14311,N14312,N14313,N14314,N14315,N14316,
  N14317,N14318,N14319,N14320,N14321,N14322,N14323,N14324,N14325,N14326,N14327,
  N14328,N14329,N14330,N14331,N14332,N14333,N14334,N14335,N14336,N14337,N14338,N14339,
  N14340,N14341,N14342,N14343,N14344,N14345,N14346,N14347,N14348,N14349,N14350,
  N14351,N14352,N14353,N14354,N14355,N14356,N14357,N14358,N14359,N14360,N14361,
  N14362,N14363,N14364,N14365,N14366,N14367,N14368,N14369,N14370,N14371,N14372,N14373,
  N14374,N14375,N14376,N14377,N14378,N14379,N14380,N14381,N14382,N14383,N14384,
  N14385,N14386,N14387,N14388,N14389,N14390,N14391,N14392,N14393,N14394,N14395,N14396,
  N14397,N14398,N14399,N14400,N14401,N14402,N14403,N14404,N14405,N14406,N14407,
  N14408,N14409,N14410,N14411,N14412,N14413,N14414,N14415,N14416,N14417,N14418,N14419,
  N14420,N14421,N14422,N14423,N14424,N14425,N14426,N14427,N14428,N14429,N14430,
  N14431,N14432,N14433,N14434,N14435,N14436,N14437,N14438,N14439,N14440,N14441,
  N14442,N14443,N14444,N14445,N14446,N14447,N14448,N14449,N14450,N14451,N14452,N14453,
  N14454,N14455,N14456,N14457,N14458,N14459,N14460,N14461,N14462,N14463,N14464,
  N14465,N14466,N14467,N14468,N14469,N14470,N14471,N14472,N14473,N14474,N14475,N14476,
  N14477,N14478,N14479,N14480,N14481,N14482,N14483,N14484,N14485,N14486,N14487,
  N14488,N14489,N14490,N14491,N14492,N14493,N14494,N14495,N14496,N14497,N14498,N14499,
  N14500,N14501,N14502,N14503,N14504,N14505,N14506,N14507,N14508,N14509,N14510,
  N14511,N14512,N14513,N14514,N14515,N14516,N14517,N14518,N14519,N14520,N14521,
  N14522,N14523,N14524,N14525,N14526,N14527,N14528,N14529,N14530,N14531,N14532,N14533,
  N14534,N14535,N14536,N14537,N14538,N14539,N14540,N14541,N14542,N14543,N14544,
  N14545,N14546,N14547,N14548,N14549,N14550,N14551,N14552,N14553,N14554,N14555,N14556,
  N14557,N14558,N14559,N14560,N14561,N14562,N14563,N14564,N14565,N14566,N14567,
  N14568,N14569,N14570,N14571,N14572,N14573,N14574,N14575,N14576,N14577,N14578,N14579,
  N14580,N14581,N14582,N14583,N14584,N14585,N14586,N14587,N14588,N14589,N14590,
  N14591,N14592,N14593,N14594,N14595,N14596,N14597,N14598,N14599,N14600,N14601,
  N14602,N14603,N14604,N14605,N14606,N14607,N14608,N14609,N14610,N14611,N14612,N14613,
  N14614,N14615,N14616,N14617,N14618,N14619,N14620,N14621,N14622,N14623,N14624,
  N14625,N14626,N14627,N14628,N14629,N14630,N14631,N14632,N14633,N14634,N14635,N14636,
  N14637,N14638,N14639,N14640,N14641,N14642,N14643,N14644,N14645,N14646,N14647,
  N14648,N14649,N14650,N14651,N14652,N14653,N14654,N14655,N14656,N14657,N14658,N14659,
  N14660,N14661,N14662,N14663,N14664,N14665,N14666,N14667,N14668,N14669,N14670,
  N14671,N14672,N14673,N14674,N14675,N14676,N14677,N14678,N14679,N14680,N14681,
  N14682,N14683,N14684,N14685,N14686,N14687,N14688,N14689,N14690,N14691,N14692,N14693,
  N14694,N14695,N14696,N14697,N14698,N14699,N14700,N14701,N14702,N14703,N14704,
  N14705,N14706,N14707,N14708,N14709,N14710,N14711,N14712,N14713,N14714,N14715,N14716,
  N14717,N14718,N14719,N14720,N14721,N14722,N14723,N14724,N14725,N14726,N14727,
  N14728,N14729,N14730,N14731,N14732,N14733,N14734,N14735,N14736,N14737,N14738,N14739,
  N14740,N14741,N14742,N14743,N14744,N14745,N14746,N14747,N14748,N14749,N14750,
  N14751,N14752,N14753,N14754,N14755,N14756,N14757,N14758,N14759,N14760,N14761,
  N14762,N14763,N14764,N14765,N14766,N14767,N14768,N14769,N14770,N14771,N14772,N14773,
  N14774,N14775,N14776,N14777,N14778,N14779,N14780,N14781,N14782,N14783,N14784,
  N14785,N14786,N14787,N14788,N14789,N14790,N14791,N14792,N14793,N14794,N14795,N14796,
  N14797,N14798,N14799,N14800,N14801,N14802,N14803,N14804,N14805,N14806,N14807,
  N14808,N14809,N14810,N14811,N14812,N14813,N14814,N14815,N14816,N14817,N14818,N14819,
  N14820,N14821,N14822,N14823,N14824,N14825,N14826,N14827,N14828,N14829,N14830,
  N14831,N14832,N14833,N14834,N14835,N14836,N14837,N14838,N14839,N14840,N14841,
  N14842,N14843,N14844,N14845,N14846,N14847,N14848,N14849,N14850,N14851,N14852,N14853,
  N14854,N14855,N14856,N14857,N14858,N14859,N14860,N14861,N14862,N14863,N14864,
  N14865,N14866,N14867,N14868,N14869,N14870,N14871,N14872,N14873,N14874,N14875,N14876,
  N14877,N14878,N14879,N14880,N14881,N14882,N14883,N14884,N14885,N14886,N14887,
  N14888,N14889,N14890,N14891,N14892,N14893,N14894,N14895,N14896,N14897,N14898,N14899,
  N14900,N14901,N14902,N14903,N14904,N14905,N14906,N14907,N14908,N14909,N14910,
  N14911,N14912,N14913,N14914,N14915,N14916,N14917,N14918,N14919,N14920,N14921,
  N14922,N14923,N14924,N14925,N14926,N14927,N14928,N14929,N14930,N14931,N14932,N14933,
  N14934,N14935,N14936,N14937,N14938,N14939,N14940,N14941,N14942,N14943,N14944,
  N14945,N14946,N14947,N14948,N14949,N14950,N14951,N14952,N14953,N14954,N14955,N14956,
  N14957,N14958,N14959,N14960,N14961,N14962,N14963,N14964,N14965,N14966,N14967,
  N14968,N14969,N14970,N14971,N14972,N14973,N14974,N14975,N14976,N14977,N14978,N14979,
  N14980,N14981,N14982,N14983,N14984,N14985,N14986,N14987,N14988,N14989,N14990,
  N14991,N14992,N14993,N14994,N14995,N14996,N14997,N14998,N14999,N15000,N15001,
  N15002,N15003,N15004,N15005,N15006,N15007,N15008,N15009,N15010,N15011,N15012,N15013,
  N15014,N15015,N15016,N15017,N15018,N15019,N15020,N15021,N15022,N15023,N15024,
  N15025,N15026,N15027,N15028,N15029,N15030,N15031,N15032,N15033,N15034,N15035,N15036,
  N15037,N15038,N15039,N15040,N15041,N15042,N15043,N15044,N15045,N15046,N15047,
  N15048,N15049,N15050,N15051,N15052,N15053,N15054,N15055,N15056,N15057,N15058,N15059,
  N15060,N15061,N15062,N15063,N15064,N15065,N15066,N15067,N15068,N15069,N15070,
  N15071,N15072,N15073,N15074,N15075,N15076,N15077,N15078,N15079,N15080,N15081,
  N15082,N15083,N15084,N15085,N15086,N15087,N15088,N15089,N15090,N15091,N15092,N15093,
  N15094,N15095,N15096,N15097,N15098,N15099,N15100,N15101,N15102,N15103,N15104,
  N15105,N15106,N15107,N15108,N15109,N15110,N15111,N15112,N15113,N15114,N15115,N15116,
  N15117,N15118,N15119,N15120,N15121,N15122,N15123,N15124,N15125,N15126,N15127,
  N15128,N15129,N15130,N15131,N15132,N15133,N15134,N15135,N15136,N15137,N15138,N15139,
  N15140,N15141,N15142,N15143,N15144,N15145,N15146,N15147,N15148,N15149,N15150,
  N15151,N15152,N15153,N15154,N15155,N15156,N15157,N15158,N15159,N15160,N15161,
  N15162,N15163,N15164,N15165,N15166,N15167,N15168,N15169,N15170,N15171,N15172,N15173,
  N15174,N15175,N15176,N15177,N15178,N15179,N15180,N15181,N15182,N15183,N15184,
  N15185,N15186,N15187,N15188,N15189,N15190,N15191,N15192,N15193,N15194,N15195,N15196,
  N15197,N15198,N15199,N15200,N15201,N15202,N15203,N15204,N15205,N15206,N15207,
  N15208,N15209,N15210,N15211,N15212,N15213,N15214,N15215,N15216,N15217,N15218,N15219,
  N15220,N15221,N15222,N15223,N15224,N15225,N15226,N15227,N15228,N15229,N15230,
  N15231,N15232,N15233,N15234,N15235,N15236,N15237,N15238,N15239,N15240,N15241,
  N15242,N15243,N15244,N15245,N15246,N15247,N15248,N15249,N15250,N15251,N15252,N15253,
  N15254,N15255,N15256,N15257,N15258,N15259,N15260,N15261,N15262,N15263,N15264,
  N15265,N15266,N15267,N15268,N15269,N15270,N15271,N15272,N15273,N15274,N15275,N15276,
  N15277,N15278,N15279,N15280,N15281,N15282,N15283,N15284,N15285,N15286,N15287,
  N15288,N15289,N15290,N15291,N15292,N15293,N15294,N15295,N15296,N15297,N15298,N15299,
  N15300,N15301,N15302,N15303,N15304,N15305,N15306,N15307,N15308,N15309,N15310,
  N15311,N15312,N15313,N15314,N15315,N15316,N15317,N15318,N15319,N15320,N15321,
  N15322,N15323,N15324,N15325,N15326,N15327,N15328,N15329,N15330,N15331,N15332,N15333,
  N15334,N15335,N15336,N15337,N15338,N15339,N15340,N15341,N15342,N15343,N15344,
  N15345,N15346,N15347,N15348,N15349,N15350,N15351,N15352,N15353,N15354,N15355,N15356,
  N15357,N15358,N15359,N15360,N15361,N15362,N15363,N15364,N15365,N15366,N15367,
  N15368,N15369,N15370,N15371,N15372,N15373,N15374,N15375,N15376,N15377,N15378,N15379,
  N15380,N15381,N15382,N15383,N15384,N15385,N15386,N15387,N15388,N15389,N15390,
  N15391,N15392,N15393,N15394,N15395,N15396,N15397,N15398,N15399,N15400,N15401,
  N15402,N15403,N15404,N15405,N15406,N15407,N15408,N15409,N15410,N15411,N15412,N15413,
  N15414,N15415,N15416,N15417,N15418,N15419,N15420,N15421,N15422,N15423,N15424,
  N15425,N15426,N15427,N15428,N15429,N15430,N15431,N15432,N15433,N15434,N15435,N15436,
  N15437,N15438,N15439,N15440,N15441,N15442,N15443,N15444,N15445,N15446,N15447,
  N15448,N15449,N15450,N15451,N15452,N15453,N15454,N15455,N15456,N15457,N15458,N15459,
  N15460,N15461,N15462,N15463,N15464,N15465,N15466,N15467,N15468,N15469,N15470,
  N15471,N15472,N15473,N15474,N15475,N15476,N15477,N15478,N15479,N15480,N15481,
  N15482,N15483,N15484,N15485,N15486,N15487,N15488,N15489,N15490,N15491,N15492,N15493,
  N15494,N15495,N15496,N15497,N15498,N15499,N15500,N15501,N15502,N15503,N15504,
  N15505,N15506,N15507,N15508,N15509,N15510,N15511,N15512,N15513,N15514,N15515,N15516,
  N15517,N15518,N15519,N15520,N15521,N15522,N15523,N15524,N15525,N15526,N15527,
  N15528,N15529,N15530,N15531,N15532,N15533,N15534,N15535,N15536,N15537,N15538,N15539,
  N15540,N15541,N15542,N15543,N15544,N15545,N15546,N15547,N15548,N15549,N15550,
  N15551,N15552,N15553,N15554,N15555,N15556,N15557,N15558,N15559,N15560,N15561,
  N15562,N15563,N15564,N15565,N15566,N15567,N15568,N15569,N15570,N15571,N15572,N15573,
  N15574,N15575,N15576,N15577,N15578,N15579,N15580,N15581,N15582,N15583,N15584,
  N15585,N15586,N15587,N15588,N15589,N15590,N15591,N15592,N15593,N15594,N15595,N15596,
  N15597,N15598,N15599,N15600,N15601,N15602,N15603,N15604,N15605,N15606,N15607,
  N15608,N15609,N15610,N15611,N15612,N15613,N15614,N15615,N15616,N15617,N15618,N15619,
  N15620,N15621,N15622,N15623,N15624,N15625,N15626,N15627,N15628,N15629,N15630,
  N15631,N15632,N15633,N15634,N15635,N15636,N15637,N15638,N15639,N15640,N15641,
  N15642,N15643,N15644,N15645,N15646,N15647,N15648,N15649,N15650,N15651,N15652,N15653,
  N15654,N15655,N15656,N15657,N15658,N15659,N15660,N15661,N15662,N15663,N15664,
  N15665,N15666,N15667,N15668,N15669,N15670,N15671,N15672,N15673,N15674,N15675,N15676,
  N15677,N15678,N15679,N15680,N15681,N15682,N15683,N15684,N15685,N15686,N15687,
  N15688,N15689,N15690,N15691,N15692,N15693,N15694,N15695,N15696,N15697,N15698,N15699,
  N15700,N15701,N15702,N15703,N15704,N15705,N15706,N15707,N15708,N15709,N15710,
  N15711,N15712,N15713,N15714,N15715,N15716,N15717,N15718,N15719,N15720,N15721,
  N15722,N15723,N15724,N15725,N15726,N15727,N15728,N15729,N15730,N15731,N15732,N15733,
  N15734,N15735,N15736,N15737,N15738,N15739,N15740,N15741,N15742,N15743,N15744,
  N15745,N15746,N15747,N15748,N15749,N15750,N15751,N15752,N15753,N15754,N15755,N15756,
  N15757,N15758,N15759,N15760,N15761,N15762,N15763,N15764,N15765,N15766,N15767,
  N15768,N15769,N15770,N15771,N15772,N15773,N15774,N15775,N15776,N15777,N15778,N15779,
  N15780,N15781,N15782,N15783,N15784,N15785,N15786,N15787,N15788,N15789,N15790,
  N15791,N15792,N15793,N15794,N15795,N15796,N15797,N15798,N15799,N15800,N15801,
  N15802,N15803,N15804,N15805,N15806,N15807,N15808,N15809,N15810,N15811,N15812,N15813,
  N15814,N15815,N15816,N15817,N15818,N15819,N15820,N15821,N15822,N15823,N15824,
  N15825,N15826,N15827,N15828,N15829,N15830,N15831,N15832,N15833,N15834,N15835,N15836,
  N15837,N15838,N15839,N15840,N15841,N15842,N15843,N15844,N15845,N15846,N15847,
  N15848,N15849,N15850,N15851,N15852,N15853,N15854,N15855,N15856,N15857,N15858,N15859,
  N15860,N15861,N15862,N15863,N15864,N15865,N15866,N15867,N15868,N15869,N15870,
  N15871,N15872,N15873,N15874,N15875,N15876,N15877,N15878,N15879,N15880,N15881,
  N15882,N15883,N15884,N15885,N15886,N15887,N15888,N15889,N15890,N15891,N15892,N15893,
  N15894,N15895,N15896,N15897,N15898,N15899,N15900,N15901,N15902,N15903,N15904,
  N15905,N15906,N15907,N15908,N15909,N15910,N15911,N15912,N15913,N15914,N15915,N15916,
  N15917,N15918,N15919,N15920,N15921,N15922,N15923,N15924,N15925,N15926,N15927,
  N15928,N15929,N15930,N15931,N15932,N15933,N15934,N15935,N15936,N15937,N15938,N15939,
  N15940,N15941,N15942,N15943,N15944,N15945,N15946,N15947,N15948,N15949,N15950,
  N15951,N15952,N15953,N15954,N15955,N15956,N15957,N15958,N15959,N15960,N15961,
  N15962,N15963,N15964,N15965,N15966,N15967,N15968,N15969,N15970,N15971,N15972,N15973,
  N15974,N15975,N15976,N15977,N15978,N15979,N15980,N15981,N15982,N15983,N15984,
  N15985,N15986,N15987,N15988,N15989,N15990,N15991,N15992,N15993,N15994,N15995,N15996,
  N15997,N15998,N15999,N16000,N16001,N16002,N16003,N16004,N16005,N16006,N16007,
  N16008,N16009,N16010,N16011,N16012,N16013,N16014,N16015,N16016,N16017,N16018,N16019,
  N16020,N16021,N16022,N16023,N16024,N16025,N16026,N16027,N16028,N16029,N16030,
  N16031,N16032,N16033,N16034,N16035,N16036,N16037,N16038,N16039,N16040,N16041,
  N16042,N16043,N16044,N16045,N16046,N16047,N16048,N16049,N16050,N16051,N16052,N16053,
  N16054,N16055,N16056,N16057,N16058,N16059,N16060,N16061,N16062,N16063,N16064,
  N16065,N16066,N16067,N16068,N16069,N16070,N16071,N16072,N16073,N16074,N16075,N16076,
  N16077,N16078,N16079,N16080,N16081,N16082,N16083,N16084,N16085,N16086,N16087,
  N16088,N16089,N16090,N16091,N16092,N16093,N16094,N16095,N16096,N16097,N16098,N16099,
  N16100,N16101,N16102,N16103,N16104,N16105,N16106,N16107,N16108,N16109,N16110,
  N16111,N16112,N16113,N16114,N16115,N16116,N16117,N16118,N16119,N16120,N16121,
  N16122,N16123,N16124,N16125,N16126,N16127,N16128,N16129,N16130,N16131,N16132,N16133,
  N16134,N16135,N16136,N16137,N16138,N16139,N16140,N16141,N16142,N16143,N16144,
  N16145,N16146,N16147,N16148,N16149,N16150,N16151,N16152,N16153,N16154,N16155,N16156,
  N16157,N16158,N16159,N16160,N16161,N16162,N16163,N16164,N16165,N16166,N16167,
  N16168,N16169,N16170,N16171,N16172,N16173,N16174,N16175,N16176,N16177,N16178,N16179,
  N16180,N16181,N16182,N16183,N16184,N16185,N16186,N16187,N16188,N16189,N16190,
  N16191,N16192,N16193,N16194,N16195,N16196,N16197,N16198,N16199,N16200,N16201,
  N16202,N16203,N16204,N16205,N16206,N16207,N16208,N16209,N16210,N16211,N16212,N16213,
  N16214,N16215,N16216,N16217,N16218,N16219,N16220,N16221,N16222,N16223,N16224,
  N16225,N16226,N16227,N16228,N16229,N16230,N16231,N16232,N16233,N16234,N16235,N16236,
  N16237,N16238,N16239,N16240,N16241,N16242,N16243,N16244,N16245,N16246,N16247,
  N16248,N16249,N16250,N16251,N16252,N16253,N16254,N16255,N16256,N16257,N16258,N16259,
  N16260,N16261,N16262,N16263,N16264,N16265,N16266,N16267,N16268,N16269,N16270,
  N16271,N16272,N16273,N16274,N16275,N16276,N16277,N16278,N16279,N16280,N16281,
  N16282,N16283,N16284,N16285,N16286,N16287,N16288,N16289,N16290,N16291,N16292,N16293,
  N16294,N16295,N16296,N16297,N16298,N16299,N16300,N16301,N16302,N16303,N16304,
  N16305,N16306,N16307,N16308,N16309,N16310,N16311,N16312,N16313,N16314,N16315,N16316,
  N16317,N16318,N16319,N16320,N16321,N16322,N16323,N16324,N16325,N16326,N16327,
  N16328,N16329,N16330,N16331,N16332,N16333,N16334,N16335,N16336,N16337,N16338,N16339,
  N16340,N16341,N16342,N16343,N16344,N16345,N16346,N16347,N16348,N16349,N16350,
  N16351,N16352,N16353,N16354,N16355,N16356,N16357,N16358,N16359,N16360,N16361,
  N16362,N16363,N16364,N16365,N16366,N16367,N16368,N16369,N16370,N16371,N16372,N16373,
  N16374,N16375,N16376,N16377,N16378,N16379,N16380,N16381,N16382,N16383,N16384,
  N16385,N16386,N16387,N16388,N16389,N16390,N16391,N16392,N16393,N16394,N16395,N16396,
  N16397,N16398,N16399,N16400,N16401,N16402,N16403,N16404,N16405,N16406,N16407,
  N16408,N16409,N16410,N16411,N16412,N16413,N16414,N16415,N16416,N16417,N16418,N16419,
  N16420,N16421,N16422,N16423,N16424,N16425,N16426,N16427,N16428,N16429,N16430,
  N16431,N16432,N16433,N16434,N16435,N16436,N16437,N16438,N16439,N16440,N16441,
  N16442,N16443,N16444,N16445,N16446,N16447,N16448,N16449,N16450,N16451,N16452,N16453,
  N16454,N16455,N16456,N16457,N16458,N16459,N16460,N16461,N16462,N16463,N16464,
  N16465,N16466,N16467,N16468,N16469,N16470,N16471,N16472,N16473,N16474,N16475,N16476,
  N16477,N16478,N16479,N16480,N16481,N16482,N16483,N16484,N16485,N16486,N16487,
  N16488,N16489,N16490,N16491,N16492,N16493,N16494,N16495,N16496,N16497,N16498,N16499,
  N16500,N16501,N16502,N16503,N16504,N16505,N16506,N16507,N16508,N16509,N16510,
  N16511,N16512,N16513,N16514,N16515,N16516,N16517,N16518,N16519,N16520,N16521,
  N16522,N16523,N16524,N16525,N16526,N16527,N16528,N16529,N16530,N16531,N16532,N16533,
  N16534,N16535,N16536,N16537,N16538,N16539,N16540,N16541,N16542,N16543,N16544,
  N16545,N16546,N16547,N16548,N16549,N16550,N16551,N16552,N16553,N16554,N16555,N16556,
  N16557,N16558,N16559,N16560,N16561,N16562,N16563,N16564,N16565,N16566,N16567,
  N16568,N16569,N16570,N16571,N16572,N16573,N16574,N16575,N16576,N16577,N16578,N16579,
  N16580,N16581,N16582,N16583,N16584,N16585,N16586,N16587,N16588,N16589,N16590,
  N16591,N16592,N16593,N16594,N16595,N16596,N16597,N16598,N16599,N16600,N16601,
  N16602,N16603,N16604,N16605,N16606,N16607,N16608,N16609,N16610,N16611,N16612,N16613,
  N16614,N16615,N16616,N16617,N16618,N16619,N16620,N16621,N16622,N16623,N16624,
  N16625,N16626,N16627,N16628,N16629,N16630,N16631,N16632,N16633,N16634;
  wire [1023:0] mem;
  reg mem_1023_sv2v_reg,mem_1022_sv2v_reg,mem_1021_sv2v_reg,mem_1020_sv2v_reg,
  mem_1019_sv2v_reg,mem_1018_sv2v_reg,mem_1017_sv2v_reg,mem_1016_sv2v_reg,
  mem_1015_sv2v_reg,mem_1014_sv2v_reg,mem_1013_sv2v_reg,mem_1012_sv2v_reg,mem_1011_sv2v_reg,
  mem_1010_sv2v_reg,mem_1009_sv2v_reg,mem_1008_sv2v_reg,mem_1007_sv2v_reg,
  mem_1006_sv2v_reg,mem_1005_sv2v_reg,mem_1004_sv2v_reg,mem_1003_sv2v_reg,mem_1002_sv2v_reg,
  mem_1001_sv2v_reg,mem_1000_sv2v_reg,mem_999_sv2v_reg,mem_998_sv2v_reg,
  mem_997_sv2v_reg,mem_996_sv2v_reg,mem_995_sv2v_reg,mem_994_sv2v_reg,mem_993_sv2v_reg,
  mem_992_sv2v_reg,mem_991_sv2v_reg,mem_990_sv2v_reg,mem_989_sv2v_reg,mem_988_sv2v_reg,
  mem_987_sv2v_reg,mem_986_sv2v_reg,mem_985_sv2v_reg,mem_984_sv2v_reg,
  mem_983_sv2v_reg,mem_982_sv2v_reg,mem_981_sv2v_reg,mem_980_sv2v_reg,mem_979_sv2v_reg,
  mem_978_sv2v_reg,mem_977_sv2v_reg,mem_976_sv2v_reg,mem_975_sv2v_reg,mem_974_sv2v_reg,
  mem_973_sv2v_reg,mem_972_sv2v_reg,mem_971_sv2v_reg,mem_970_sv2v_reg,mem_969_sv2v_reg,
  mem_968_sv2v_reg,mem_967_sv2v_reg,mem_966_sv2v_reg,mem_965_sv2v_reg,
  mem_964_sv2v_reg,mem_963_sv2v_reg,mem_962_sv2v_reg,mem_961_sv2v_reg,mem_960_sv2v_reg,
  mem_959_sv2v_reg,mem_958_sv2v_reg,mem_957_sv2v_reg,mem_956_sv2v_reg,mem_955_sv2v_reg,
  mem_954_sv2v_reg,mem_953_sv2v_reg,mem_952_sv2v_reg,mem_951_sv2v_reg,
  mem_950_sv2v_reg,mem_949_sv2v_reg,mem_948_sv2v_reg,mem_947_sv2v_reg,mem_946_sv2v_reg,
  mem_945_sv2v_reg,mem_944_sv2v_reg,mem_943_sv2v_reg,mem_942_sv2v_reg,mem_941_sv2v_reg,
  mem_940_sv2v_reg,mem_939_sv2v_reg,mem_938_sv2v_reg,mem_937_sv2v_reg,mem_936_sv2v_reg,
  mem_935_sv2v_reg,mem_934_sv2v_reg,mem_933_sv2v_reg,mem_932_sv2v_reg,
  mem_931_sv2v_reg,mem_930_sv2v_reg,mem_929_sv2v_reg,mem_928_sv2v_reg,mem_927_sv2v_reg,
  mem_926_sv2v_reg,mem_925_sv2v_reg,mem_924_sv2v_reg,mem_923_sv2v_reg,mem_922_sv2v_reg,
  mem_921_sv2v_reg,mem_920_sv2v_reg,mem_919_sv2v_reg,mem_918_sv2v_reg,
  mem_917_sv2v_reg,mem_916_sv2v_reg,mem_915_sv2v_reg,mem_914_sv2v_reg,mem_913_sv2v_reg,
  mem_912_sv2v_reg,mem_911_sv2v_reg,mem_910_sv2v_reg,mem_909_sv2v_reg,mem_908_sv2v_reg,
  mem_907_sv2v_reg,mem_906_sv2v_reg,mem_905_sv2v_reg,mem_904_sv2v_reg,
  mem_903_sv2v_reg,mem_902_sv2v_reg,mem_901_sv2v_reg,mem_900_sv2v_reg,mem_899_sv2v_reg,
  mem_898_sv2v_reg,mem_897_sv2v_reg,mem_896_sv2v_reg,mem_895_sv2v_reg,mem_894_sv2v_reg,
  mem_893_sv2v_reg,mem_892_sv2v_reg,mem_891_sv2v_reg,mem_890_sv2v_reg,mem_889_sv2v_reg,
  mem_888_sv2v_reg,mem_887_sv2v_reg,mem_886_sv2v_reg,mem_885_sv2v_reg,
  mem_884_sv2v_reg,mem_883_sv2v_reg,mem_882_sv2v_reg,mem_881_sv2v_reg,mem_880_sv2v_reg,
  mem_879_sv2v_reg,mem_878_sv2v_reg,mem_877_sv2v_reg,mem_876_sv2v_reg,mem_875_sv2v_reg,
  mem_874_sv2v_reg,mem_873_sv2v_reg,mem_872_sv2v_reg,mem_871_sv2v_reg,
  mem_870_sv2v_reg,mem_869_sv2v_reg,mem_868_sv2v_reg,mem_867_sv2v_reg,mem_866_sv2v_reg,
  mem_865_sv2v_reg,mem_864_sv2v_reg,mem_863_sv2v_reg,mem_862_sv2v_reg,mem_861_sv2v_reg,
  mem_860_sv2v_reg,mem_859_sv2v_reg,mem_858_sv2v_reg,mem_857_sv2v_reg,mem_856_sv2v_reg,
  mem_855_sv2v_reg,mem_854_sv2v_reg,mem_853_sv2v_reg,mem_852_sv2v_reg,
  mem_851_sv2v_reg,mem_850_sv2v_reg,mem_849_sv2v_reg,mem_848_sv2v_reg,mem_847_sv2v_reg,
  mem_846_sv2v_reg,mem_845_sv2v_reg,mem_844_sv2v_reg,mem_843_sv2v_reg,mem_842_sv2v_reg,
  mem_841_sv2v_reg,mem_840_sv2v_reg,mem_839_sv2v_reg,mem_838_sv2v_reg,
  mem_837_sv2v_reg,mem_836_sv2v_reg,mem_835_sv2v_reg,mem_834_sv2v_reg,mem_833_sv2v_reg,
  mem_832_sv2v_reg,mem_831_sv2v_reg,mem_830_sv2v_reg,mem_829_sv2v_reg,mem_828_sv2v_reg,
  mem_827_sv2v_reg,mem_826_sv2v_reg,mem_825_sv2v_reg,mem_824_sv2v_reg,
  mem_823_sv2v_reg,mem_822_sv2v_reg,mem_821_sv2v_reg,mem_820_sv2v_reg,mem_819_sv2v_reg,
  mem_818_sv2v_reg,mem_817_sv2v_reg,mem_816_sv2v_reg,mem_815_sv2v_reg,mem_814_sv2v_reg,
  mem_813_sv2v_reg,mem_812_sv2v_reg,mem_811_sv2v_reg,mem_810_sv2v_reg,mem_809_sv2v_reg,
  mem_808_sv2v_reg,mem_807_sv2v_reg,mem_806_sv2v_reg,mem_805_sv2v_reg,
  mem_804_sv2v_reg,mem_803_sv2v_reg,mem_802_sv2v_reg,mem_801_sv2v_reg,mem_800_sv2v_reg,
  mem_799_sv2v_reg,mem_798_sv2v_reg,mem_797_sv2v_reg,mem_796_sv2v_reg,mem_795_sv2v_reg,
  mem_794_sv2v_reg,mem_793_sv2v_reg,mem_792_sv2v_reg,mem_791_sv2v_reg,
  mem_790_sv2v_reg,mem_789_sv2v_reg,mem_788_sv2v_reg,mem_787_sv2v_reg,mem_786_sv2v_reg,
  mem_785_sv2v_reg,mem_784_sv2v_reg,mem_783_sv2v_reg,mem_782_sv2v_reg,mem_781_sv2v_reg,
  mem_780_sv2v_reg,mem_779_sv2v_reg,mem_778_sv2v_reg,mem_777_sv2v_reg,mem_776_sv2v_reg,
  mem_775_sv2v_reg,mem_774_sv2v_reg,mem_773_sv2v_reg,mem_772_sv2v_reg,
  mem_771_sv2v_reg,mem_770_sv2v_reg,mem_769_sv2v_reg,mem_768_sv2v_reg,mem_767_sv2v_reg,
  mem_766_sv2v_reg,mem_765_sv2v_reg,mem_764_sv2v_reg,mem_763_sv2v_reg,mem_762_sv2v_reg,
  mem_761_sv2v_reg,mem_760_sv2v_reg,mem_759_sv2v_reg,mem_758_sv2v_reg,
  mem_757_sv2v_reg,mem_756_sv2v_reg,mem_755_sv2v_reg,mem_754_sv2v_reg,mem_753_sv2v_reg,
  mem_752_sv2v_reg,mem_751_sv2v_reg,mem_750_sv2v_reg,mem_749_sv2v_reg,mem_748_sv2v_reg,
  mem_747_sv2v_reg,mem_746_sv2v_reg,mem_745_sv2v_reg,mem_744_sv2v_reg,
  mem_743_sv2v_reg,mem_742_sv2v_reg,mem_741_sv2v_reg,mem_740_sv2v_reg,mem_739_sv2v_reg,
  mem_738_sv2v_reg,mem_737_sv2v_reg,mem_736_sv2v_reg,mem_735_sv2v_reg,mem_734_sv2v_reg,
  mem_733_sv2v_reg,mem_732_sv2v_reg,mem_731_sv2v_reg,mem_730_sv2v_reg,mem_729_sv2v_reg,
  mem_728_sv2v_reg,mem_727_sv2v_reg,mem_726_sv2v_reg,mem_725_sv2v_reg,
  mem_724_sv2v_reg,mem_723_sv2v_reg,mem_722_sv2v_reg,mem_721_sv2v_reg,mem_720_sv2v_reg,
  mem_719_sv2v_reg,mem_718_sv2v_reg,mem_717_sv2v_reg,mem_716_sv2v_reg,mem_715_sv2v_reg,
  mem_714_sv2v_reg,mem_713_sv2v_reg,mem_712_sv2v_reg,mem_711_sv2v_reg,
  mem_710_sv2v_reg,mem_709_sv2v_reg,mem_708_sv2v_reg,mem_707_sv2v_reg,mem_706_sv2v_reg,
  mem_705_sv2v_reg,mem_704_sv2v_reg,mem_703_sv2v_reg,mem_702_sv2v_reg,mem_701_sv2v_reg,
  mem_700_sv2v_reg,mem_699_sv2v_reg,mem_698_sv2v_reg,mem_697_sv2v_reg,mem_696_sv2v_reg,
  mem_695_sv2v_reg,mem_694_sv2v_reg,mem_693_sv2v_reg,mem_692_sv2v_reg,
  mem_691_sv2v_reg,mem_690_sv2v_reg,mem_689_sv2v_reg,mem_688_sv2v_reg,mem_687_sv2v_reg,
  mem_686_sv2v_reg,mem_685_sv2v_reg,mem_684_sv2v_reg,mem_683_sv2v_reg,mem_682_sv2v_reg,
  mem_681_sv2v_reg,mem_680_sv2v_reg,mem_679_sv2v_reg,mem_678_sv2v_reg,
  mem_677_sv2v_reg,mem_676_sv2v_reg,mem_675_sv2v_reg,mem_674_sv2v_reg,mem_673_sv2v_reg,
  mem_672_sv2v_reg,mem_671_sv2v_reg,mem_670_sv2v_reg,mem_669_sv2v_reg,mem_668_sv2v_reg,
  mem_667_sv2v_reg,mem_666_sv2v_reg,mem_665_sv2v_reg,mem_664_sv2v_reg,
  mem_663_sv2v_reg,mem_662_sv2v_reg,mem_661_sv2v_reg,mem_660_sv2v_reg,mem_659_sv2v_reg,
  mem_658_sv2v_reg,mem_657_sv2v_reg,mem_656_sv2v_reg,mem_655_sv2v_reg,mem_654_sv2v_reg,
  mem_653_sv2v_reg,mem_652_sv2v_reg,mem_651_sv2v_reg,mem_650_sv2v_reg,mem_649_sv2v_reg,
  mem_648_sv2v_reg,mem_647_sv2v_reg,mem_646_sv2v_reg,mem_645_sv2v_reg,
  mem_644_sv2v_reg,mem_643_sv2v_reg,mem_642_sv2v_reg,mem_641_sv2v_reg,mem_640_sv2v_reg,
  mem_639_sv2v_reg,mem_638_sv2v_reg,mem_637_sv2v_reg,mem_636_sv2v_reg,mem_635_sv2v_reg,
  mem_634_sv2v_reg,mem_633_sv2v_reg,mem_632_sv2v_reg,mem_631_sv2v_reg,
  mem_630_sv2v_reg,mem_629_sv2v_reg,mem_628_sv2v_reg,mem_627_sv2v_reg,mem_626_sv2v_reg,
  mem_625_sv2v_reg,mem_624_sv2v_reg,mem_623_sv2v_reg,mem_622_sv2v_reg,mem_621_sv2v_reg,
  mem_620_sv2v_reg,mem_619_sv2v_reg,mem_618_sv2v_reg,mem_617_sv2v_reg,mem_616_sv2v_reg,
  mem_615_sv2v_reg,mem_614_sv2v_reg,mem_613_sv2v_reg,mem_612_sv2v_reg,
  mem_611_sv2v_reg,mem_610_sv2v_reg,mem_609_sv2v_reg,mem_608_sv2v_reg,mem_607_sv2v_reg,
  mem_606_sv2v_reg,mem_605_sv2v_reg,mem_604_sv2v_reg,mem_603_sv2v_reg,mem_602_sv2v_reg,
  mem_601_sv2v_reg,mem_600_sv2v_reg,mem_599_sv2v_reg,mem_598_sv2v_reg,
  mem_597_sv2v_reg,mem_596_sv2v_reg,mem_595_sv2v_reg,mem_594_sv2v_reg,mem_593_sv2v_reg,
  mem_592_sv2v_reg,mem_591_sv2v_reg,mem_590_sv2v_reg,mem_589_sv2v_reg,mem_588_sv2v_reg,
  mem_587_sv2v_reg,mem_586_sv2v_reg,mem_585_sv2v_reg,mem_584_sv2v_reg,
  mem_583_sv2v_reg,mem_582_sv2v_reg,mem_581_sv2v_reg,mem_580_sv2v_reg,mem_579_sv2v_reg,
  mem_578_sv2v_reg,mem_577_sv2v_reg,mem_576_sv2v_reg,mem_575_sv2v_reg,mem_574_sv2v_reg,
  mem_573_sv2v_reg,mem_572_sv2v_reg,mem_571_sv2v_reg,mem_570_sv2v_reg,mem_569_sv2v_reg,
  mem_568_sv2v_reg,mem_567_sv2v_reg,mem_566_sv2v_reg,mem_565_sv2v_reg,
  mem_564_sv2v_reg,mem_563_sv2v_reg,mem_562_sv2v_reg,mem_561_sv2v_reg,mem_560_sv2v_reg,
  mem_559_sv2v_reg,mem_558_sv2v_reg,mem_557_sv2v_reg,mem_556_sv2v_reg,mem_555_sv2v_reg,
  mem_554_sv2v_reg,mem_553_sv2v_reg,mem_552_sv2v_reg,mem_551_sv2v_reg,
  mem_550_sv2v_reg,mem_549_sv2v_reg,mem_548_sv2v_reg,mem_547_sv2v_reg,mem_546_sv2v_reg,
  mem_545_sv2v_reg,mem_544_sv2v_reg,mem_543_sv2v_reg,mem_542_sv2v_reg,mem_541_sv2v_reg,
  mem_540_sv2v_reg,mem_539_sv2v_reg,mem_538_sv2v_reg,mem_537_sv2v_reg,mem_536_sv2v_reg,
  mem_535_sv2v_reg,mem_534_sv2v_reg,mem_533_sv2v_reg,mem_532_sv2v_reg,
  mem_531_sv2v_reg,mem_530_sv2v_reg,mem_529_sv2v_reg,mem_528_sv2v_reg,mem_527_sv2v_reg,
  mem_526_sv2v_reg,mem_525_sv2v_reg,mem_524_sv2v_reg,mem_523_sv2v_reg,mem_522_sv2v_reg,
  mem_521_sv2v_reg,mem_520_sv2v_reg,mem_519_sv2v_reg,mem_518_sv2v_reg,
  mem_517_sv2v_reg,mem_516_sv2v_reg,mem_515_sv2v_reg,mem_514_sv2v_reg,mem_513_sv2v_reg,
  mem_512_sv2v_reg,mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,
  mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,
  mem_503_sv2v_reg,mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,
  mem_498_sv2v_reg,mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,
  mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,
  mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,
  mem_484_sv2v_reg,mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,
  mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,
  mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,
  mem_470_sv2v_reg,mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,
  mem_465_sv2v_reg,mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,
  mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,
  mem_451_sv2v_reg,mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,
  mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,
  mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,
  mem_437_sv2v_reg,mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,
  mem_432_sv2v_reg,mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,
  mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,
  mem_423_sv2v_reg,mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,
  mem_418_sv2v_reg,mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,
  mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,
  mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,
  mem_404_sv2v_reg,mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,
  mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,
  mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,
  mem_390_sv2v_reg,mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,
  mem_385_sv2v_reg,mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,
  mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,
  mem_371_sv2v_reg,mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,
  mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,
  mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,
  mem_357_sv2v_reg,mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,
  mem_352_sv2v_reg,mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,
  mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,
  mem_343_sv2v_reg,mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,
  mem_338_sv2v_reg,mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,
  mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,
  mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,
  mem_324_sv2v_reg,mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,
  mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,
  mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,
  mem_310_sv2v_reg,mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,
  mem_305_sv2v_reg,mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,
  mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,
  mem_291_sv2v_reg,mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,
  mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,
  mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,
  mem_277_sv2v_reg,mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,
  mem_272_sv2v_reg,mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,
  mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,
  mem_263_sv2v_reg,mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,
  mem_258_sv2v_reg,mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,
  mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,
  mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,
  mem_244_sv2v_reg,mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,
  mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,
  mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,
  mem_230_sv2v_reg,mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,
  mem_225_sv2v_reg,mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,
  mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,
  mem_211_sv2v_reg,mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,
  mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,
  mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,
  mem_197_sv2v_reg,mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,
  mem_192_sv2v_reg,mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,
  mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,
  mem_183_sv2v_reg,mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,
  mem_178_sv2v_reg,mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,
  mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,
  mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,
  mem_164_sv2v_reg,mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,
  mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,
  mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,
  mem_150_sv2v_reg,mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,
  mem_145_sv2v_reg,mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,
  mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,
  mem_131_sv2v_reg,mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,
  mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,
  mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,
  mem_117_sv2v_reg,mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,
  mem_112_sv2v_reg,mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,
  mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,
  mem_103_sv2v_reg,mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,
  mem_98_sv2v_reg,mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,
  mem_93_sv2v_reg,mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,
  mem_88_sv2v_reg,mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,
  mem_83_sv2v_reg,mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,
  mem_78_sv2v_reg,mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,
  mem_73_sv2v_reg,mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,
  mem_68_sv2v_reg,mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,
  mem_63_sv2v_reg,mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,
  mem_58_sv2v_reg,mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,
  mem_53_sv2v_reg,mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,
  mem_48_sv2v_reg,mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,
  mem_43_sv2v_reg,mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,
  mem_38_sv2v_reg,mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,
  mem_33_sv2v_reg,mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,
  mem_28_sv2v_reg,mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,
  mem_23_sv2v_reg,mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,
  mem_18_sv2v_reg,mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,
  mem_13_sv2v_reg,mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,
  mem_8_sv2v_reg,mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,
  mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[1023] = mem_1023_sv2v_reg;
  assign mem[1022] = mem_1022_sv2v_reg;
  assign mem[1021] = mem_1021_sv2v_reg;
  assign mem[1020] = mem_1020_sv2v_reg;
  assign mem[1019] = mem_1019_sv2v_reg;
  assign mem[1018] = mem_1018_sv2v_reg;
  assign mem[1017] = mem_1017_sv2v_reg;
  assign mem[1016] = mem_1016_sv2v_reg;
  assign mem[1015] = mem_1015_sv2v_reg;
  assign mem[1014] = mem_1014_sv2v_reg;
  assign mem[1013] = mem_1013_sv2v_reg;
  assign mem[1012] = mem_1012_sv2v_reg;
  assign mem[1011] = mem_1011_sv2v_reg;
  assign mem[1010] = mem_1010_sv2v_reg;
  assign mem[1009] = mem_1009_sv2v_reg;
  assign mem[1008] = mem_1008_sv2v_reg;
  assign mem[1007] = mem_1007_sv2v_reg;
  assign mem[1006] = mem_1006_sv2v_reg;
  assign mem[1005] = mem_1005_sv2v_reg;
  assign mem[1004] = mem_1004_sv2v_reg;
  assign mem[1003] = mem_1003_sv2v_reg;
  assign mem[1002] = mem_1002_sv2v_reg;
  assign mem[1001] = mem_1001_sv2v_reg;
  assign mem[1000] = mem_1000_sv2v_reg;
  assign mem[999] = mem_999_sv2v_reg;
  assign mem[998] = mem_998_sv2v_reg;
  assign mem[997] = mem_997_sv2v_reg;
  assign mem[996] = mem_996_sv2v_reg;
  assign mem[995] = mem_995_sv2v_reg;
  assign mem[994] = mem_994_sv2v_reg;
  assign mem[993] = mem_993_sv2v_reg;
  assign mem[992] = mem_992_sv2v_reg;
  assign mem[991] = mem_991_sv2v_reg;
  assign mem[990] = mem_990_sv2v_reg;
  assign mem[989] = mem_989_sv2v_reg;
  assign mem[988] = mem_988_sv2v_reg;
  assign mem[987] = mem_987_sv2v_reg;
  assign mem[986] = mem_986_sv2v_reg;
  assign mem[985] = mem_985_sv2v_reg;
  assign mem[984] = mem_984_sv2v_reg;
  assign mem[983] = mem_983_sv2v_reg;
  assign mem[982] = mem_982_sv2v_reg;
  assign mem[981] = mem_981_sv2v_reg;
  assign mem[980] = mem_980_sv2v_reg;
  assign mem[979] = mem_979_sv2v_reg;
  assign mem[978] = mem_978_sv2v_reg;
  assign mem[977] = mem_977_sv2v_reg;
  assign mem[976] = mem_976_sv2v_reg;
  assign mem[975] = mem_975_sv2v_reg;
  assign mem[974] = mem_974_sv2v_reg;
  assign mem[973] = mem_973_sv2v_reg;
  assign mem[972] = mem_972_sv2v_reg;
  assign mem[971] = mem_971_sv2v_reg;
  assign mem[970] = mem_970_sv2v_reg;
  assign mem[969] = mem_969_sv2v_reg;
  assign mem[968] = mem_968_sv2v_reg;
  assign mem[967] = mem_967_sv2v_reg;
  assign mem[966] = mem_966_sv2v_reg;
  assign mem[965] = mem_965_sv2v_reg;
  assign mem[964] = mem_964_sv2v_reg;
  assign mem[963] = mem_963_sv2v_reg;
  assign mem[962] = mem_962_sv2v_reg;
  assign mem[961] = mem_961_sv2v_reg;
  assign mem[960] = mem_960_sv2v_reg;
  assign mem[959] = mem_959_sv2v_reg;
  assign mem[958] = mem_958_sv2v_reg;
  assign mem[957] = mem_957_sv2v_reg;
  assign mem[956] = mem_956_sv2v_reg;
  assign mem[955] = mem_955_sv2v_reg;
  assign mem[954] = mem_954_sv2v_reg;
  assign mem[953] = mem_953_sv2v_reg;
  assign mem[952] = mem_952_sv2v_reg;
  assign mem[951] = mem_951_sv2v_reg;
  assign mem[950] = mem_950_sv2v_reg;
  assign mem[949] = mem_949_sv2v_reg;
  assign mem[948] = mem_948_sv2v_reg;
  assign mem[947] = mem_947_sv2v_reg;
  assign mem[946] = mem_946_sv2v_reg;
  assign mem[945] = mem_945_sv2v_reg;
  assign mem[944] = mem_944_sv2v_reg;
  assign mem[943] = mem_943_sv2v_reg;
  assign mem[942] = mem_942_sv2v_reg;
  assign mem[941] = mem_941_sv2v_reg;
  assign mem[940] = mem_940_sv2v_reg;
  assign mem[939] = mem_939_sv2v_reg;
  assign mem[938] = mem_938_sv2v_reg;
  assign mem[937] = mem_937_sv2v_reg;
  assign mem[936] = mem_936_sv2v_reg;
  assign mem[935] = mem_935_sv2v_reg;
  assign mem[934] = mem_934_sv2v_reg;
  assign mem[933] = mem_933_sv2v_reg;
  assign mem[932] = mem_932_sv2v_reg;
  assign mem[931] = mem_931_sv2v_reg;
  assign mem[930] = mem_930_sv2v_reg;
  assign mem[929] = mem_929_sv2v_reg;
  assign mem[928] = mem_928_sv2v_reg;
  assign mem[927] = mem_927_sv2v_reg;
  assign mem[926] = mem_926_sv2v_reg;
  assign mem[925] = mem_925_sv2v_reg;
  assign mem[924] = mem_924_sv2v_reg;
  assign mem[923] = mem_923_sv2v_reg;
  assign mem[922] = mem_922_sv2v_reg;
  assign mem[921] = mem_921_sv2v_reg;
  assign mem[920] = mem_920_sv2v_reg;
  assign mem[919] = mem_919_sv2v_reg;
  assign mem[918] = mem_918_sv2v_reg;
  assign mem[917] = mem_917_sv2v_reg;
  assign mem[916] = mem_916_sv2v_reg;
  assign mem[915] = mem_915_sv2v_reg;
  assign mem[914] = mem_914_sv2v_reg;
  assign mem[913] = mem_913_sv2v_reg;
  assign mem[912] = mem_912_sv2v_reg;
  assign mem[911] = mem_911_sv2v_reg;
  assign mem[910] = mem_910_sv2v_reg;
  assign mem[909] = mem_909_sv2v_reg;
  assign mem[908] = mem_908_sv2v_reg;
  assign mem[907] = mem_907_sv2v_reg;
  assign mem[906] = mem_906_sv2v_reg;
  assign mem[905] = mem_905_sv2v_reg;
  assign mem[904] = mem_904_sv2v_reg;
  assign mem[903] = mem_903_sv2v_reg;
  assign mem[902] = mem_902_sv2v_reg;
  assign mem[901] = mem_901_sv2v_reg;
  assign mem[900] = mem_900_sv2v_reg;
  assign mem[899] = mem_899_sv2v_reg;
  assign mem[898] = mem_898_sv2v_reg;
  assign mem[897] = mem_897_sv2v_reg;
  assign mem[896] = mem_896_sv2v_reg;
  assign mem[895] = mem_895_sv2v_reg;
  assign mem[894] = mem_894_sv2v_reg;
  assign mem[893] = mem_893_sv2v_reg;
  assign mem[892] = mem_892_sv2v_reg;
  assign mem[891] = mem_891_sv2v_reg;
  assign mem[890] = mem_890_sv2v_reg;
  assign mem[889] = mem_889_sv2v_reg;
  assign mem[888] = mem_888_sv2v_reg;
  assign mem[887] = mem_887_sv2v_reg;
  assign mem[886] = mem_886_sv2v_reg;
  assign mem[885] = mem_885_sv2v_reg;
  assign mem[884] = mem_884_sv2v_reg;
  assign mem[883] = mem_883_sv2v_reg;
  assign mem[882] = mem_882_sv2v_reg;
  assign mem[881] = mem_881_sv2v_reg;
  assign mem[880] = mem_880_sv2v_reg;
  assign mem[879] = mem_879_sv2v_reg;
  assign mem[878] = mem_878_sv2v_reg;
  assign mem[877] = mem_877_sv2v_reg;
  assign mem[876] = mem_876_sv2v_reg;
  assign mem[875] = mem_875_sv2v_reg;
  assign mem[874] = mem_874_sv2v_reg;
  assign mem[873] = mem_873_sv2v_reg;
  assign mem[872] = mem_872_sv2v_reg;
  assign mem[871] = mem_871_sv2v_reg;
  assign mem[870] = mem_870_sv2v_reg;
  assign mem[869] = mem_869_sv2v_reg;
  assign mem[868] = mem_868_sv2v_reg;
  assign mem[867] = mem_867_sv2v_reg;
  assign mem[866] = mem_866_sv2v_reg;
  assign mem[865] = mem_865_sv2v_reg;
  assign mem[864] = mem_864_sv2v_reg;
  assign mem[863] = mem_863_sv2v_reg;
  assign mem[862] = mem_862_sv2v_reg;
  assign mem[861] = mem_861_sv2v_reg;
  assign mem[860] = mem_860_sv2v_reg;
  assign mem[859] = mem_859_sv2v_reg;
  assign mem[858] = mem_858_sv2v_reg;
  assign mem[857] = mem_857_sv2v_reg;
  assign mem[856] = mem_856_sv2v_reg;
  assign mem[855] = mem_855_sv2v_reg;
  assign mem[854] = mem_854_sv2v_reg;
  assign mem[853] = mem_853_sv2v_reg;
  assign mem[852] = mem_852_sv2v_reg;
  assign mem[851] = mem_851_sv2v_reg;
  assign mem[850] = mem_850_sv2v_reg;
  assign mem[849] = mem_849_sv2v_reg;
  assign mem[848] = mem_848_sv2v_reg;
  assign mem[847] = mem_847_sv2v_reg;
  assign mem[846] = mem_846_sv2v_reg;
  assign mem[845] = mem_845_sv2v_reg;
  assign mem[844] = mem_844_sv2v_reg;
  assign mem[843] = mem_843_sv2v_reg;
  assign mem[842] = mem_842_sv2v_reg;
  assign mem[841] = mem_841_sv2v_reg;
  assign mem[840] = mem_840_sv2v_reg;
  assign mem[839] = mem_839_sv2v_reg;
  assign mem[838] = mem_838_sv2v_reg;
  assign mem[837] = mem_837_sv2v_reg;
  assign mem[836] = mem_836_sv2v_reg;
  assign mem[835] = mem_835_sv2v_reg;
  assign mem[834] = mem_834_sv2v_reg;
  assign mem[833] = mem_833_sv2v_reg;
  assign mem[832] = mem_832_sv2v_reg;
  assign mem[831] = mem_831_sv2v_reg;
  assign mem[830] = mem_830_sv2v_reg;
  assign mem[829] = mem_829_sv2v_reg;
  assign mem[828] = mem_828_sv2v_reg;
  assign mem[827] = mem_827_sv2v_reg;
  assign mem[826] = mem_826_sv2v_reg;
  assign mem[825] = mem_825_sv2v_reg;
  assign mem[824] = mem_824_sv2v_reg;
  assign mem[823] = mem_823_sv2v_reg;
  assign mem[822] = mem_822_sv2v_reg;
  assign mem[821] = mem_821_sv2v_reg;
  assign mem[820] = mem_820_sv2v_reg;
  assign mem[819] = mem_819_sv2v_reg;
  assign mem[818] = mem_818_sv2v_reg;
  assign mem[817] = mem_817_sv2v_reg;
  assign mem[816] = mem_816_sv2v_reg;
  assign mem[815] = mem_815_sv2v_reg;
  assign mem[814] = mem_814_sv2v_reg;
  assign mem[813] = mem_813_sv2v_reg;
  assign mem[812] = mem_812_sv2v_reg;
  assign mem[811] = mem_811_sv2v_reg;
  assign mem[810] = mem_810_sv2v_reg;
  assign mem[809] = mem_809_sv2v_reg;
  assign mem[808] = mem_808_sv2v_reg;
  assign mem[807] = mem_807_sv2v_reg;
  assign mem[806] = mem_806_sv2v_reg;
  assign mem[805] = mem_805_sv2v_reg;
  assign mem[804] = mem_804_sv2v_reg;
  assign mem[803] = mem_803_sv2v_reg;
  assign mem[802] = mem_802_sv2v_reg;
  assign mem[801] = mem_801_sv2v_reg;
  assign mem[800] = mem_800_sv2v_reg;
  assign mem[799] = mem_799_sv2v_reg;
  assign mem[798] = mem_798_sv2v_reg;
  assign mem[797] = mem_797_sv2v_reg;
  assign mem[796] = mem_796_sv2v_reg;
  assign mem[795] = mem_795_sv2v_reg;
  assign mem[794] = mem_794_sv2v_reg;
  assign mem[793] = mem_793_sv2v_reg;
  assign mem[792] = mem_792_sv2v_reg;
  assign mem[791] = mem_791_sv2v_reg;
  assign mem[790] = mem_790_sv2v_reg;
  assign mem[789] = mem_789_sv2v_reg;
  assign mem[788] = mem_788_sv2v_reg;
  assign mem[787] = mem_787_sv2v_reg;
  assign mem[786] = mem_786_sv2v_reg;
  assign mem[785] = mem_785_sv2v_reg;
  assign mem[784] = mem_784_sv2v_reg;
  assign mem[783] = mem_783_sv2v_reg;
  assign mem[782] = mem_782_sv2v_reg;
  assign mem[781] = mem_781_sv2v_reg;
  assign mem[780] = mem_780_sv2v_reg;
  assign mem[779] = mem_779_sv2v_reg;
  assign mem[778] = mem_778_sv2v_reg;
  assign mem[777] = mem_777_sv2v_reg;
  assign mem[776] = mem_776_sv2v_reg;
  assign mem[775] = mem_775_sv2v_reg;
  assign mem[774] = mem_774_sv2v_reg;
  assign mem[773] = mem_773_sv2v_reg;
  assign mem[772] = mem_772_sv2v_reg;
  assign mem[771] = mem_771_sv2v_reg;
  assign mem[770] = mem_770_sv2v_reg;
  assign mem[769] = mem_769_sv2v_reg;
  assign mem[768] = mem_768_sv2v_reg;
  assign mem[767] = mem_767_sv2v_reg;
  assign mem[766] = mem_766_sv2v_reg;
  assign mem[765] = mem_765_sv2v_reg;
  assign mem[764] = mem_764_sv2v_reg;
  assign mem[763] = mem_763_sv2v_reg;
  assign mem[762] = mem_762_sv2v_reg;
  assign mem[761] = mem_761_sv2v_reg;
  assign mem[760] = mem_760_sv2v_reg;
  assign mem[759] = mem_759_sv2v_reg;
  assign mem[758] = mem_758_sv2v_reg;
  assign mem[757] = mem_757_sv2v_reg;
  assign mem[756] = mem_756_sv2v_reg;
  assign mem[755] = mem_755_sv2v_reg;
  assign mem[754] = mem_754_sv2v_reg;
  assign mem[753] = mem_753_sv2v_reg;
  assign mem[752] = mem_752_sv2v_reg;
  assign mem[751] = mem_751_sv2v_reg;
  assign mem[750] = mem_750_sv2v_reg;
  assign mem[749] = mem_749_sv2v_reg;
  assign mem[748] = mem_748_sv2v_reg;
  assign mem[747] = mem_747_sv2v_reg;
  assign mem[746] = mem_746_sv2v_reg;
  assign mem[745] = mem_745_sv2v_reg;
  assign mem[744] = mem_744_sv2v_reg;
  assign mem[743] = mem_743_sv2v_reg;
  assign mem[742] = mem_742_sv2v_reg;
  assign mem[741] = mem_741_sv2v_reg;
  assign mem[740] = mem_740_sv2v_reg;
  assign mem[739] = mem_739_sv2v_reg;
  assign mem[738] = mem_738_sv2v_reg;
  assign mem[737] = mem_737_sv2v_reg;
  assign mem[736] = mem_736_sv2v_reg;
  assign mem[735] = mem_735_sv2v_reg;
  assign mem[734] = mem_734_sv2v_reg;
  assign mem[733] = mem_733_sv2v_reg;
  assign mem[732] = mem_732_sv2v_reg;
  assign mem[731] = mem_731_sv2v_reg;
  assign mem[730] = mem_730_sv2v_reg;
  assign mem[729] = mem_729_sv2v_reg;
  assign mem[728] = mem_728_sv2v_reg;
  assign mem[727] = mem_727_sv2v_reg;
  assign mem[726] = mem_726_sv2v_reg;
  assign mem[725] = mem_725_sv2v_reg;
  assign mem[724] = mem_724_sv2v_reg;
  assign mem[723] = mem_723_sv2v_reg;
  assign mem[722] = mem_722_sv2v_reg;
  assign mem[721] = mem_721_sv2v_reg;
  assign mem[720] = mem_720_sv2v_reg;
  assign mem[719] = mem_719_sv2v_reg;
  assign mem[718] = mem_718_sv2v_reg;
  assign mem[717] = mem_717_sv2v_reg;
  assign mem[716] = mem_716_sv2v_reg;
  assign mem[715] = mem_715_sv2v_reg;
  assign mem[714] = mem_714_sv2v_reg;
  assign mem[713] = mem_713_sv2v_reg;
  assign mem[712] = mem_712_sv2v_reg;
  assign mem[711] = mem_711_sv2v_reg;
  assign mem[710] = mem_710_sv2v_reg;
  assign mem[709] = mem_709_sv2v_reg;
  assign mem[708] = mem_708_sv2v_reg;
  assign mem[707] = mem_707_sv2v_reg;
  assign mem[706] = mem_706_sv2v_reg;
  assign mem[705] = mem_705_sv2v_reg;
  assign mem[704] = mem_704_sv2v_reg;
  assign mem[703] = mem_703_sv2v_reg;
  assign mem[702] = mem_702_sv2v_reg;
  assign mem[701] = mem_701_sv2v_reg;
  assign mem[700] = mem_700_sv2v_reg;
  assign mem[699] = mem_699_sv2v_reg;
  assign mem[698] = mem_698_sv2v_reg;
  assign mem[697] = mem_697_sv2v_reg;
  assign mem[696] = mem_696_sv2v_reg;
  assign mem[695] = mem_695_sv2v_reg;
  assign mem[694] = mem_694_sv2v_reg;
  assign mem[693] = mem_693_sv2v_reg;
  assign mem[692] = mem_692_sv2v_reg;
  assign mem[691] = mem_691_sv2v_reg;
  assign mem[690] = mem_690_sv2v_reg;
  assign mem[689] = mem_689_sv2v_reg;
  assign mem[688] = mem_688_sv2v_reg;
  assign mem[687] = mem_687_sv2v_reg;
  assign mem[686] = mem_686_sv2v_reg;
  assign mem[685] = mem_685_sv2v_reg;
  assign mem[684] = mem_684_sv2v_reg;
  assign mem[683] = mem_683_sv2v_reg;
  assign mem[682] = mem_682_sv2v_reg;
  assign mem[681] = mem_681_sv2v_reg;
  assign mem[680] = mem_680_sv2v_reg;
  assign mem[679] = mem_679_sv2v_reg;
  assign mem[678] = mem_678_sv2v_reg;
  assign mem[677] = mem_677_sv2v_reg;
  assign mem[676] = mem_676_sv2v_reg;
  assign mem[675] = mem_675_sv2v_reg;
  assign mem[674] = mem_674_sv2v_reg;
  assign mem[673] = mem_673_sv2v_reg;
  assign mem[672] = mem_672_sv2v_reg;
  assign mem[671] = mem_671_sv2v_reg;
  assign mem[670] = mem_670_sv2v_reg;
  assign mem[669] = mem_669_sv2v_reg;
  assign mem[668] = mem_668_sv2v_reg;
  assign mem[667] = mem_667_sv2v_reg;
  assign mem[666] = mem_666_sv2v_reg;
  assign mem[665] = mem_665_sv2v_reg;
  assign mem[664] = mem_664_sv2v_reg;
  assign mem[663] = mem_663_sv2v_reg;
  assign mem[662] = mem_662_sv2v_reg;
  assign mem[661] = mem_661_sv2v_reg;
  assign mem[660] = mem_660_sv2v_reg;
  assign mem[659] = mem_659_sv2v_reg;
  assign mem[658] = mem_658_sv2v_reg;
  assign mem[657] = mem_657_sv2v_reg;
  assign mem[656] = mem_656_sv2v_reg;
  assign mem[655] = mem_655_sv2v_reg;
  assign mem[654] = mem_654_sv2v_reg;
  assign mem[653] = mem_653_sv2v_reg;
  assign mem[652] = mem_652_sv2v_reg;
  assign mem[651] = mem_651_sv2v_reg;
  assign mem[650] = mem_650_sv2v_reg;
  assign mem[649] = mem_649_sv2v_reg;
  assign mem[648] = mem_648_sv2v_reg;
  assign mem[647] = mem_647_sv2v_reg;
  assign mem[646] = mem_646_sv2v_reg;
  assign mem[645] = mem_645_sv2v_reg;
  assign mem[644] = mem_644_sv2v_reg;
  assign mem[643] = mem_643_sv2v_reg;
  assign mem[642] = mem_642_sv2v_reg;
  assign mem[641] = mem_641_sv2v_reg;
  assign mem[640] = mem_640_sv2v_reg;
  assign mem[639] = mem_639_sv2v_reg;
  assign mem[638] = mem_638_sv2v_reg;
  assign mem[637] = mem_637_sv2v_reg;
  assign mem[636] = mem_636_sv2v_reg;
  assign mem[635] = mem_635_sv2v_reg;
  assign mem[634] = mem_634_sv2v_reg;
  assign mem[633] = mem_633_sv2v_reg;
  assign mem[632] = mem_632_sv2v_reg;
  assign mem[631] = mem_631_sv2v_reg;
  assign mem[630] = mem_630_sv2v_reg;
  assign mem[629] = mem_629_sv2v_reg;
  assign mem[628] = mem_628_sv2v_reg;
  assign mem[627] = mem_627_sv2v_reg;
  assign mem[626] = mem_626_sv2v_reg;
  assign mem[625] = mem_625_sv2v_reg;
  assign mem[624] = mem_624_sv2v_reg;
  assign mem[623] = mem_623_sv2v_reg;
  assign mem[622] = mem_622_sv2v_reg;
  assign mem[621] = mem_621_sv2v_reg;
  assign mem[620] = mem_620_sv2v_reg;
  assign mem[619] = mem_619_sv2v_reg;
  assign mem[618] = mem_618_sv2v_reg;
  assign mem[617] = mem_617_sv2v_reg;
  assign mem[616] = mem_616_sv2v_reg;
  assign mem[615] = mem_615_sv2v_reg;
  assign mem[614] = mem_614_sv2v_reg;
  assign mem[613] = mem_613_sv2v_reg;
  assign mem[612] = mem_612_sv2v_reg;
  assign mem[611] = mem_611_sv2v_reg;
  assign mem[610] = mem_610_sv2v_reg;
  assign mem[609] = mem_609_sv2v_reg;
  assign mem[608] = mem_608_sv2v_reg;
  assign mem[607] = mem_607_sv2v_reg;
  assign mem[606] = mem_606_sv2v_reg;
  assign mem[605] = mem_605_sv2v_reg;
  assign mem[604] = mem_604_sv2v_reg;
  assign mem[603] = mem_603_sv2v_reg;
  assign mem[602] = mem_602_sv2v_reg;
  assign mem[601] = mem_601_sv2v_reg;
  assign mem[600] = mem_600_sv2v_reg;
  assign mem[599] = mem_599_sv2v_reg;
  assign mem[598] = mem_598_sv2v_reg;
  assign mem[597] = mem_597_sv2v_reg;
  assign mem[596] = mem_596_sv2v_reg;
  assign mem[595] = mem_595_sv2v_reg;
  assign mem[594] = mem_594_sv2v_reg;
  assign mem[593] = mem_593_sv2v_reg;
  assign mem[592] = mem_592_sv2v_reg;
  assign mem[591] = mem_591_sv2v_reg;
  assign mem[590] = mem_590_sv2v_reg;
  assign mem[589] = mem_589_sv2v_reg;
  assign mem[588] = mem_588_sv2v_reg;
  assign mem[587] = mem_587_sv2v_reg;
  assign mem[586] = mem_586_sv2v_reg;
  assign mem[585] = mem_585_sv2v_reg;
  assign mem[584] = mem_584_sv2v_reg;
  assign mem[583] = mem_583_sv2v_reg;
  assign mem[582] = mem_582_sv2v_reg;
  assign mem[581] = mem_581_sv2v_reg;
  assign mem[580] = mem_580_sv2v_reg;
  assign mem[579] = mem_579_sv2v_reg;
  assign mem[578] = mem_578_sv2v_reg;
  assign mem[577] = mem_577_sv2v_reg;
  assign mem[576] = mem_576_sv2v_reg;
  assign mem[575] = mem_575_sv2v_reg;
  assign mem[574] = mem_574_sv2v_reg;
  assign mem[573] = mem_573_sv2v_reg;
  assign mem[572] = mem_572_sv2v_reg;
  assign mem[571] = mem_571_sv2v_reg;
  assign mem[570] = mem_570_sv2v_reg;
  assign mem[569] = mem_569_sv2v_reg;
  assign mem[568] = mem_568_sv2v_reg;
  assign mem[567] = mem_567_sv2v_reg;
  assign mem[566] = mem_566_sv2v_reg;
  assign mem[565] = mem_565_sv2v_reg;
  assign mem[564] = mem_564_sv2v_reg;
  assign mem[563] = mem_563_sv2v_reg;
  assign mem[562] = mem_562_sv2v_reg;
  assign mem[561] = mem_561_sv2v_reg;
  assign mem[560] = mem_560_sv2v_reg;
  assign mem[559] = mem_559_sv2v_reg;
  assign mem[558] = mem_558_sv2v_reg;
  assign mem[557] = mem_557_sv2v_reg;
  assign mem[556] = mem_556_sv2v_reg;
  assign mem[555] = mem_555_sv2v_reg;
  assign mem[554] = mem_554_sv2v_reg;
  assign mem[553] = mem_553_sv2v_reg;
  assign mem[552] = mem_552_sv2v_reg;
  assign mem[551] = mem_551_sv2v_reg;
  assign mem[550] = mem_550_sv2v_reg;
  assign mem[549] = mem_549_sv2v_reg;
  assign mem[548] = mem_548_sv2v_reg;
  assign mem[547] = mem_547_sv2v_reg;
  assign mem[546] = mem_546_sv2v_reg;
  assign mem[545] = mem_545_sv2v_reg;
  assign mem[544] = mem_544_sv2v_reg;
  assign mem[543] = mem_543_sv2v_reg;
  assign mem[542] = mem_542_sv2v_reg;
  assign mem[541] = mem_541_sv2v_reg;
  assign mem[540] = mem_540_sv2v_reg;
  assign mem[539] = mem_539_sv2v_reg;
  assign mem[538] = mem_538_sv2v_reg;
  assign mem[537] = mem_537_sv2v_reg;
  assign mem[536] = mem_536_sv2v_reg;
  assign mem[535] = mem_535_sv2v_reg;
  assign mem[534] = mem_534_sv2v_reg;
  assign mem[533] = mem_533_sv2v_reg;
  assign mem[532] = mem_532_sv2v_reg;
  assign mem[531] = mem_531_sv2v_reg;
  assign mem[530] = mem_530_sv2v_reg;
  assign mem[529] = mem_529_sv2v_reg;
  assign mem[528] = mem_528_sv2v_reg;
  assign mem[527] = mem_527_sv2v_reg;
  assign mem[526] = mem_526_sv2v_reg;
  assign mem[525] = mem_525_sv2v_reg;
  assign mem[524] = mem_524_sv2v_reg;
  assign mem[523] = mem_523_sv2v_reg;
  assign mem[522] = mem_522_sv2v_reg;
  assign mem[521] = mem_521_sv2v_reg;
  assign mem[520] = mem_520_sv2v_reg;
  assign mem[519] = mem_519_sv2v_reg;
  assign mem[518] = mem_518_sv2v_reg;
  assign mem[517] = mem_517_sv2v_reg;
  assign mem[516] = mem_516_sv2v_reg;
  assign mem[515] = mem_515_sv2v_reg;
  assign mem[514] = mem_514_sv2v_reg;
  assign mem[513] = mem_513_sv2v_reg;
  assign mem[512] = mem_512_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign N1057 = (N545)? mem[1] : 
                 (N547)? mem[3] : 
                 (N549)? mem[5] : 
                 (N551)? mem[7] : 
                 (N553)? mem[9] : 
                 (N555)? mem[11] : 
                 (N557)? mem[13] : 
                 (N559)? mem[15] : 
                 (N561)? mem[17] : 
                 (N563)? mem[19] : 
                 (N565)? mem[21] : 
                 (N567)? mem[23] : 
                 (N569)? mem[25] : 
                 (N571)? mem[27] : 
                 (N573)? mem[29] : 
                 (N575)? mem[31] : 
                 (N577)? mem[33] : 
                 (N579)? mem[35] : 
                 (N581)? mem[37] : 
                 (N583)? mem[39] : 
                 (N585)? mem[41] : 
                 (N587)? mem[43] : 
                 (N589)? mem[45] : 
                 (N591)? mem[47] : 
                 (N593)? mem[49] : 
                 (N595)? mem[51] : 
                 (N597)? mem[53] : 
                 (N599)? mem[55] : 
                 (N601)? mem[57] : 
                 (N603)? mem[59] : 
                 (N605)? mem[61] : 
                 (N607)? mem[63] : 
                 (N609)? mem[65] : 
                 (N611)? mem[67] : 
                 (N613)? mem[69] : 
                 (N615)? mem[71] : 
                 (N617)? mem[73] : 
                 (N619)? mem[75] : 
                 (N621)? mem[77] : 
                 (N623)? mem[79] : 
                 (N625)? mem[81] : 
                 (N627)? mem[83] : 
                 (N629)? mem[85] : 
                 (N631)? mem[87] : 
                 (N633)? mem[89] : 
                 (N635)? mem[91] : 
                 (N637)? mem[93] : 
                 (N639)? mem[95] : 
                 (N641)? mem[97] : 
                 (N643)? mem[99] : 
                 (N645)? mem[101] : 
                 (N647)? mem[103] : 
                 (N649)? mem[105] : 
                 (N651)? mem[107] : 
                 (N653)? mem[109] : 
                 (N655)? mem[111] : 
                 (N657)? mem[113] : 
                 (N659)? mem[115] : 
                 (N661)? mem[117] : 
                 (N663)? mem[119] : 
                 (N665)? mem[121] : 
                 (N667)? mem[123] : 
                 (N669)? mem[125] : 
                 (N671)? mem[127] : 
                 (N673)? mem[129] : 
                 (N675)? mem[131] : 
                 (N677)? mem[133] : 
                 (N679)? mem[135] : 
                 (N681)? mem[137] : 
                 (N683)? mem[139] : 
                 (N685)? mem[141] : 
                 (N687)? mem[143] : 
                 (N689)? mem[145] : 
                 (N691)? mem[147] : 
                 (N693)? mem[149] : 
                 (N695)? mem[151] : 
                 (N697)? mem[153] : 
                 (N699)? mem[155] : 
                 (N701)? mem[157] : 
                 (N703)? mem[159] : 
                 (N705)? mem[161] : 
                 (N707)? mem[163] : 
                 (N709)? mem[165] : 
                 (N711)? mem[167] : 
                 (N713)? mem[169] : 
                 (N715)? mem[171] : 
                 (N717)? mem[173] : 
                 (N719)? mem[175] : 
                 (N721)? mem[177] : 
                 (N723)? mem[179] : 
                 (N725)? mem[181] : 
                 (N727)? mem[183] : 
                 (N729)? mem[185] : 
                 (N731)? mem[187] : 
                 (N733)? mem[189] : 
                 (N735)? mem[191] : 
                 (N737)? mem[193] : 
                 (N739)? mem[195] : 
                 (N741)? mem[197] : 
                 (N743)? mem[199] : 
                 (N745)? mem[201] : 
                 (N747)? mem[203] : 
                 (N749)? mem[205] : 
                 (N751)? mem[207] : 
                 (N753)? mem[209] : 
                 (N755)? mem[211] : 
                 (N757)? mem[213] : 
                 (N759)? mem[215] : 
                 (N761)? mem[217] : 
                 (N763)? mem[219] : 
                 (N765)? mem[221] : 
                 (N767)? mem[223] : 
                 (N769)? mem[225] : 
                 (N771)? mem[227] : 
                 (N773)? mem[229] : 
                 (N775)? mem[231] : 
                 (N777)? mem[233] : 
                 (N779)? mem[235] : 
                 (N781)? mem[237] : 
                 (N783)? mem[239] : 
                 (N785)? mem[241] : 
                 (N787)? mem[243] : 
                 (N789)? mem[245] : 
                 (N791)? mem[247] : 
                 (N793)? mem[249] : 
                 (N795)? mem[251] : 
                 (N797)? mem[253] : 
                 (N799)? mem[255] : 
                 (N801)? mem[257] : 
                 (N803)? mem[259] : 
                 (N805)? mem[261] : 
                 (N807)? mem[263] : 
                 (N809)? mem[265] : 
                 (N811)? mem[267] : 
                 (N813)? mem[269] : 
                 (N815)? mem[271] : 
                 (N817)? mem[273] : 
                 (N819)? mem[275] : 
                 (N821)? mem[277] : 
                 (N823)? mem[279] : 
                 (N825)? mem[281] : 
                 (N827)? mem[283] : 
                 (N829)? mem[285] : 
                 (N831)? mem[287] : 
                 (N833)? mem[289] : 
                 (N835)? mem[291] : 
                 (N837)? mem[293] : 
                 (N839)? mem[295] : 
                 (N841)? mem[297] : 
                 (N843)? mem[299] : 
                 (N845)? mem[301] : 
                 (N847)? mem[303] : 
                 (N849)? mem[305] : 
                 (N851)? mem[307] : 
                 (N853)? mem[309] : 
                 (N855)? mem[311] : 
                 (N857)? mem[313] : 
                 (N859)? mem[315] : 
                 (N861)? mem[317] : 
                 (N863)? mem[319] : 
                 (N865)? mem[321] : 
                 (N867)? mem[323] : 
                 (N869)? mem[325] : 
                 (N871)? mem[327] : 
                 (N873)? mem[329] : 
                 (N875)? mem[331] : 
                 (N877)? mem[333] : 
                 (N879)? mem[335] : 
                 (N881)? mem[337] : 
                 (N883)? mem[339] : 
                 (N885)? mem[341] : 
                 (N887)? mem[343] : 
                 (N889)? mem[345] : 
                 (N891)? mem[347] : 
                 (N893)? mem[349] : 
                 (N895)? mem[351] : 
                 (N897)? mem[353] : 
                 (N899)? mem[355] : 
                 (N901)? mem[357] : 
                 (N903)? mem[359] : 
                 (N905)? mem[361] : 
                 (N907)? mem[363] : 
                 (N909)? mem[365] : 
                 (N911)? mem[367] : 
                 (N913)? mem[369] : 
                 (N915)? mem[371] : 
                 (N917)? mem[373] : 
                 (N919)? mem[375] : 
                 (N921)? mem[377] : 
                 (N923)? mem[379] : 
                 (N925)? mem[381] : 
                 (N927)? mem[383] : 
                 (N929)? mem[385] : 
                 (N931)? mem[387] : 
                 (N933)? mem[389] : 
                 (N935)? mem[391] : 
                 (N937)? mem[393] : 
                 (N939)? mem[395] : 
                 (N941)? mem[397] : 
                 (N943)? mem[399] : 
                 (N945)? mem[401] : 
                 (N947)? mem[403] : 
                 (N949)? mem[405] : 
                 (N951)? mem[407] : 
                 (N953)? mem[409] : 
                 (N955)? mem[411] : 
                 (N957)? mem[413] : 
                 (N959)? mem[415] : 
                 (N961)? mem[417] : 
                 (N963)? mem[419] : 
                 (N965)? mem[421] : 
                 (N967)? mem[423] : 
                 (N969)? mem[425] : 
                 (N971)? mem[427] : 
                 (N973)? mem[429] : 
                 (N975)? mem[431] : 
                 (N977)? mem[433] : 
                 (N979)? mem[435] : 
                 (N981)? mem[437] : 
                 (N983)? mem[439] : 
                 (N985)? mem[441] : 
                 (N987)? mem[443] : 
                 (N989)? mem[445] : 
                 (N991)? mem[447] : 
                 (N993)? mem[449] : 
                 (N995)? mem[451] : 
                 (N997)? mem[453] : 
                 (N999)? mem[455] : 
                 (N1001)? mem[457] : 
                 (N1003)? mem[459] : 
                 (N1005)? mem[461] : 
                 (N1007)? mem[463] : 
                 (N1009)? mem[465] : 
                 (N1011)? mem[467] : 
                 (N1013)? mem[469] : 
                 (N1015)? mem[471] : 
                 (N1017)? mem[473] : 
                 (N1019)? mem[475] : 
                 (N1021)? mem[477] : 
                 (N1023)? mem[479] : 
                 (N1025)? mem[481] : 
                 (N1027)? mem[483] : 
                 (N1029)? mem[485] : 
                 (N1031)? mem[487] : 
                 (N1033)? mem[489] : 
                 (N1035)? mem[491] : 
                 (N1037)? mem[493] : 
                 (N1039)? mem[495] : 
                 (N1041)? mem[497] : 
                 (N1043)? mem[499] : 
                 (N1045)? mem[501] : 
                 (N1047)? mem[503] : 
                 (N1049)? mem[505] : 
                 (N1051)? mem[507] : 
                 (N1053)? mem[509] : 
                 (N1055)? mem[511] : 
                 (N546)? mem[513] : 
                 (N548)? mem[515] : 
                 (N550)? mem[517] : 
                 (N552)? mem[519] : 
                 (N554)? mem[521] : 
                 (N556)? mem[523] : 
                 (N558)? mem[525] : 
                 (N560)? mem[527] : 
                 (N562)? mem[529] : 
                 (N564)? mem[531] : 
                 (N566)? mem[533] : 
                 (N568)? mem[535] : 
                 (N570)? mem[537] : 
                 (N572)? mem[539] : 
                 (N574)? mem[541] : 
                 (N576)? mem[543] : 
                 (N578)? mem[545] : 
                 (N580)? mem[547] : 
                 (N582)? mem[549] : 
                 (N584)? mem[551] : 
                 (N586)? mem[553] : 
                 (N588)? mem[555] : 
                 (N590)? mem[557] : 
                 (N592)? mem[559] : 
                 (N594)? mem[561] : 
                 (N596)? mem[563] : 
                 (N598)? mem[565] : 
                 (N600)? mem[567] : 
                 (N602)? mem[569] : 
                 (N604)? mem[571] : 
                 (N606)? mem[573] : 
                 (N608)? mem[575] : 
                 (N610)? mem[577] : 
                 (N612)? mem[579] : 
                 (N614)? mem[581] : 
                 (N616)? mem[583] : 
                 (N618)? mem[585] : 
                 (N620)? mem[587] : 
                 (N622)? mem[589] : 
                 (N624)? mem[591] : 
                 (N626)? mem[593] : 
                 (N628)? mem[595] : 
                 (N630)? mem[597] : 
                 (N632)? mem[599] : 
                 (N634)? mem[601] : 
                 (N636)? mem[603] : 
                 (N638)? mem[605] : 
                 (N640)? mem[607] : 
                 (N642)? mem[609] : 
                 (N644)? mem[611] : 
                 (N646)? mem[613] : 
                 (N648)? mem[615] : 
                 (N650)? mem[617] : 
                 (N652)? mem[619] : 
                 (N654)? mem[621] : 
                 (N656)? mem[623] : 
                 (N658)? mem[625] : 
                 (N660)? mem[627] : 
                 (N662)? mem[629] : 
                 (N664)? mem[631] : 
                 (N666)? mem[633] : 
                 (N668)? mem[635] : 
                 (N670)? mem[637] : 
                 (N672)? mem[639] : 
                 (N674)? mem[641] : 
                 (N676)? mem[643] : 
                 (N678)? mem[645] : 
                 (N680)? mem[647] : 
                 (N682)? mem[649] : 
                 (N684)? mem[651] : 
                 (N686)? mem[653] : 
                 (N688)? mem[655] : 
                 (N690)? mem[657] : 
                 (N692)? mem[659] : 
                 (N694)? mem[661] : 
                 (N696)? mem[663] : 
                 (N698)? mem[665] : 
                 (N700)? mem[667] : 
                 (N702)? mem[669] : 
                 (N704)? mem[671] : 
                 (N706)? mem[673] : 
                 (N708)? mem[675] : 
                 (N710)? mem[677] : 
                 (N712)? mem[679] : 
                 (N714)? mem[681] : 
                 (N716)? mem[683] : 
                 (N718)? mem[685] : 
                 (N720)? mem[687] : 
                 (N722)? mem[689] : 
                 (N724)? mem[691] : 
                 (N726)? mem[693] : 
                 (N728)? mem[695] : 
                 (N730)? mem[697] : 
                 (N732)? mem[699] : 
                 (N734)? mem[701] : 
                 (N736)? mem[703] : 
                 (N738)? mem[705] : 
                 (N740)? mem[707] : 
                 (N742)? mem[709] : 
                 (N744)? mem[711] : 
                 (N746)? mem[713] : 
                 (N748)? mem[715] : 
                 (N750)? mem[717] : 
                 (N752)? mem[719] : 
                 (N754)? mem[721] : 
                 (N756)? mem[723] : 
                 (N758)? mem[725] : 
                 (N760)? mem[727] : 
                 (N762)? mem[729] : 
                 (N764)? mem[731] : 
                 (N766)? mem[733] : 
                 (N768)? mem[735] : 
                 (N770)? mem[737] : 
                 (N772)? mem[739] : 
                 (N774)? mem[741] : 
                 (N776)? mem[743] : 
                 (N778)? mem[745] : 
                 (N780)? mem[747] : 
                 (N782)? mem[749] : 
                 (N784)? mem[751] : 
                 (N786)? mem[753] : 
                 (N788)? mem[755] : 
                 (N790)? mem[757] : 
                 (N792)? mem[759] : 
                 (N794)? mem[761] : 
                 (N796)? mem[763] : 
                 (N798)? mem[765] : 
                 (N800)? mem[767] : 
                 (N802)? mem[769] : 
                 (N804)? mem[771] : 
                 (N806)? mem[773] : 
                 (N808)? mem[775] : 
                 (N810)? mem[777] : 
                 (N812)? mem[779] : 
                 (N814)? mem[781] : 
                 (N816)? mem[783] : 
                 (N818)? mem[785] : 
                 (N820)? mem[787] : 
                 (N822)? mem[789] : 
                 (N824)? mem[791] : 
                 (N826)? mem[793] : 
                 (N828)? mem[795] : 
                 (N830)? mem[797] : 
                 (N832)? mem[799] : 
                 (N834)? mem[801] : 
                 (N836)? mem[803] : 
                 (N838)? mem[805] : 
                 (N840)? mem[807] : 
                 (N842)? mem[809] : 
                 (N844)? mem[811] : 
                 (N846)? mem[813] : 
                 (N848)? mem[815] : 
                 (N850)? mem[817] : 
                 (N852)? mem[819] : 
                 (N854)? mem[821] : 
                 (N856)? mem[823] : 
                 (N858)? mem[825] : 
                 (N860)? mem[827] : 
                 (N862)? mem[829] : 
                 (N864)? mem[831] : 
                 (N866)? mem[833] : 
                 (N868)? mem[835] : 
                 (N870)? mem[837] : 
                 (N872)? mem[839] : 
                 (N874)? mem[841] : 
                 (N876)? mem[843] : 
                 (N878)? mem[845] : 
                 (N880)? mem[847] : 
                 (N882)? mem[849] : 
                 (N884)? mem[851] : 
                 (N886)? mem[853] : 
                 (N888)? mem[855] : 
                 (N890)? mem[857] : 
                 (N892)? mem[859] : 
                 (N894)? mem[861] : 
                 (N896)? mem[863] : 
                 (N898)? mem[865] : 
                 (N900)? mem[867] : 
                 (N902)? mem[869] : 
                 (N904)? mem[871] : 
                 (N906)? mem[873] : 
                 (N908)? mem[875] : 
                 (N910)? mem[877] : 
                 (N912)? mem[879] : 
                 (N914)? mem[881] : 
                 (N916)? mem[883] : 
                 (N918)? mem[885] : 
                 (N920)? mem[887] : 
                 (N922)? mem[889] : 
                 (N924)? mem[891] : 
                 (N926)? mem[893] : 
                 (N928)? mem[895] : 
                 (N930)? mem[897] : 
                 (N932)? mem[899] : 
                 (N934)? mem[901] : 
                 (N936)? mem[903] : 
                 (N938)? mem[905] : 
                 (N940)? mem[907] : 
                 (N942)? mem[909] : 
                 (N944)? mem[911] : 
                 (N946)? mem[913] : 
                 (N948)? mem[915] : 
                 (N950)? mem[917] : 
                 (N952)? mem[919] : 
                 (N954)? mem[921] : 
                 (N956)? mem[923] : 
                 (N958)? mem[925] : 
                 (N960)? mem[927] : 
                 (N962)? mem[929] : 
                 (N964)? mem[931] : 
                 (N966)? mem[933] : 
                 (N968)? mem[935] : 
                 (N970)? mem[937] : 
                 (N972)? mem[939] : 
                 (N974)? mem[941] : 
                 (N976)? mem[943] : 
                 (N978)? mem[945] : 
                 (N980)? mem[947] : 
                 (N982)? mem[949] : 
                 (N984)? mem[951] : 
                 (N986)? mem[953] : 
                 (N988)? mem[955] : 
                 (N990)? mem[957] : 
                 (N992)? mem[959] : 
                 (N994)? mem[961] : 
                 (N996)? mem[963] : 
                 (N998)? mem[965] : 
                 (N1000)? mem[967] : 
                 (N1002)? mem[969] : 
                 (N1004)? mem[971] : 
                 (N1006)? mem[973] : 
                 (N1008)? mem[975] : 
                 (N1010)? mem[977] : 
                 (N1012)? mem[979] : 
                 (N1014)? mem[981] : 
                 (N1016)? mem[983] : 
                 (N1018)? mem[985] : 
                 (N1020)? mem[987] : 
                 (N1022)? mem[989] : 
                 (N1024)? mem[991] : 
                 (N1026)? mem[993] : 
                 (N1028)? mem[995] : 
                 (N1030)? mem[997] : 
                 (N1032)? mem[999] : 
                 (N1034)? mem[1001] : 
                 (N1036)? mem[1003] : 
                 (N1038)? mem[1005] : 
                 (N1040)? mem[1007] : 
                 (N1042)? mem[1009] : 
                 (N1044)? mem[1011] : 
                 (N1046)? mem[1013] : 
                 (N1048)? mem[1015] : 
                 (N1050)? mem[1017] : 
                 (N1052)? mem[1019] : 
                 (N1054)? mem[1021] : 
                 (N1056)? mem[1023] : 1'b0;
  assign N1896 = (N1416)? mem[1] : 
                 (N1418)? mem[3] : 
                 (N1420)? mem[5] : 
                 (N1422)? mem[7] : 
                 (N1424)? mem[9] : 
                 (N1426)? mem[11] : 
                 (N1428)? mem[13] : 
                 (N1430)? mem[15] : 
                 (N1432)? mem[17] : 
                 (N1434)? mem[19] : 
                 (N1436)? mem[21] : 
                 (N1438)? mem[23] : 
                 (N1440)? mem[25] : 
                 (N1442)? mem[27] : 
                 (N1444)? mem[29] : 
                 (N1446)? mem[31] : 
                 (N1448)? mem[33] : 
                 (N1450)? mem[35] : 
                 (N1452)? mem[37] : 
                 (N1454)? mem[39] : 
                 (N1456)? mem[41] : 
                 (N1458)? mem[43] : 
                 (N1460)? mem[45] : 
                 (N1462)? mem[47] : 
                 (N1464)? mem[49] : 
                 (N1466)? mem[51] : 
                 (N1468)? mem[53] : 
                 (N1470)? mem[55] : 
                 (N1472)? mem[57] : 
                 (N1474)? mem[59] : 
                 (N1476)? mem[61] : 
                 (N1478)? mem[63] : 
                 (N1480)? mem[65] : 
                 (N1482)? mem[67] : 
                 (N1484)? mem[69] : 
                 (N1486)? mem[71] : 
                 (N1488)? mem[73] : 
                 (N1490)? mem[75] : 
                 (N1492)? mem[77] : 
                 (N1494)? mem[79] : 
                 (N1496)? mem[81] : 
                 (N1498)? mem[83] : 
                 (N1500)? mem[85] : 
                 (N1502)? mem[87] : 
                 (N1504)? mem[89] : 
                 (N1506)? mem[91] : 
                 (N1508)? mem[93] : 
                 (N1510)? mem[95] : 
                 (N1512)? mem[97] : 
                 (N1514)? mem[99] : 
                 (N1516)? mem[101] : 
                 (N1518)? mem[103] : 
                 (N1520)? mem[105] : 
                 (N1522)? mem[107] : 
                 (N1524)? mem[109] : 
                 (N1526)? mem[111] : 
                 (N1528)? mem[113] : 
                 (N1530)? mem[115] : 
                 (N1532)? mem[117] : 
                 (N1534)? mem[119] : 
                 (N1536)? mem[121] : 
                 (N1538)? mem[123] : 
                 (N1540)? mem[125] : 
                 (N1542)? mem[127] : 
                 (N1544)? mem[129] : 
                 (N1546)? mem[131] : 
                 (N1548)? mem[133] : 
                 (N1550)? mem[135] : 
                 (N1552)? mem[137] : 
                 (N1554)? mem[139] : 
                 (N1556)? mem[141] : 
                 (N1558)? mem[143] : 
                 (N1560)? mem[145] : 
                 (N1562)? mem[147] : 
                 (N1564)? mem[149] : 
                 (N1566)? mem[151] : 
                 (N1568)? mem[153] : 
                 (N1570)? mem[155] : 
                 (N1572)? mem[157] : 
                 (N1574)? mem[159] : 
                 (N1576)? mem[161] : 
                 (N1578)? mem[163] : 
                 (N1580)? mem[165] : 
                 (N1582)? mem[167] : 
                 (N1584)? mem[169] : 
                 (N1586)? mem[171] : 
                 (N1588)? mem[173] : 
                 (N1590)? mem[175] : 
                 (N1592)? mem[177] : 
                 (N1594)? mem[179] : 
                 (N1596)? mem[181] : 
                 (N1598)? mem[183] : 
                 (N1600)? mem[185] : 
                 (N1602)? mem[187] : 
                 (N1604)? mem[189] : 
                 (N1606)? mem[191] : 
                 (N1608)? mem[193] : 
                 (N1610)? mem[195] : 
                 (N1612)? mem[197] : 
                 (N1614)? mem[199] : 
                 (N1616)? mem[201] : 
                 (N1618)? mem[203] : 
                 (N1620)? mem[205] : 
                 (N1622)? mem[207] : 
                 (N1624)? mem[209] : 
                 (N1626)? mem[211] : 
                 (N1628)? mem[213] : 
                 (N1630)? mem[215] : 
                 (N1632)? mem[217] : 
                 (N1634)? mem[219] : 
                 (N1636)? mem[221] : 
                 (N1638)? mem[223] : 
                 (N1640)? mem[225] : 
                 (N1642)? mem[227] : 
                 (N1644)? mem[229] : 
                 (N1646)? mem[231] : 
                 (N1648)? mem[233] : 
                 (N1650)? mem[235] : 
                 (N1652)? mem[237] : 
                 (N1654)? mem[239] : 
                 (N1656)? mem[241] : 
                 (N1658)? mem[243] : 
                 (N1660)? mem[245] : 
                 (N1662)? mem[247] : 
                 (N1664)? mem[249] : 
                 (N1666)? mem[251] : 
                 (N1668)? mem[253] : 
                 (N1670)? mem[255] : 
                 (N1672)? mem[257] : 
                 (N1674)? mem[259] : 
                 (N1676)? mem[261] : 
                 (N1678)? mem[263] : 
                 (N1680)? mem[265] : 
                 (N1682)? mem[267] : 
                 (N1684)? mem[269] : 
                 (N1686)? mem[271] : 
                 (N1688)? mem[273] : 
                 (N1690)? mem[275] : 
                 (N1692)? mem[277] : 
                 (N1694)? mem[279] : 
                 (N1696)? mem[281] : 
                 (N1698)? mem[283] : 
                 (N1700)? mem[285] : 
                 (N1702)? mem[287] : 
                 (N1704)? mem[289] : 
                 (N1706)? mem[291] : 
                 (N1708)? mem[293] : 
                 (N1710)? mem[295] : 
                 (N1712)? mem[297] : 
                 (N1714)? mem[299] : 
                 (N1716)? mem[301] : 
                 (N1718)? mem[303] : 
                 (N1720)? mem[305] : 
                 (N1722)? mem[307] : 
                 (N1724)? mem[309] : 
                 (N1726)? mem[311] : 
                 (N1728)? mem[313] : 
                 (N1730)? mem[315] : 
                 (N1732)? mem[317] : 
                 (N1734)? mem[319] : 
                 (N1736)? mem[321] : 
                 (N1738)? mem[323] : 
                 (N1740)? mem[325] : 
                 (N1742)? mem[327] : 
                 (N1744)? mem[329] : 
                 (N1746)? mem[331] : 
                 (N1748)? mem[333] : 
                 (N1750)? mem[335] : 
                 (N1752)? mem[337] : 
                 (N1754)? mem[339] : 
                 (N1756)? mem[341] : 
                 (N1758)? mem[343] : 
                 (N1760)? mem[345] : 
                 (N1762)? mem[347] : 
                 (N1764)? mem[349] : 
                 (N1766)? mem[351] : 
                 (N1768)? mem[353] : 
                 (N1770)? mem[355] : 
                 (N1772)? mem[357] : 
                 (N1774)? mem[359] : 
                 (N1776)? mem[361] : 
                 (N1778)? mem[363] : 
                 (N1780)? mem[365] : 
                 (N1782)? mem[367] : 
                 (N1784)? mem[369] : 
                 (N1786)? mem[371] : 
                 (N1788)? mem[373] : 
                 (N1790)? mem[375] : 
                 (N1792)? mem[377] : 
                 (N1794)? mem[379] : 
                 (N1796)? mem[381] : 
                 (N1798)? mem[383] : 
                 (N1800)? mem[385] : 
                 (N1802)? mem[387] : 
                 (N1804)? mem[389] : 
                 (N1806)? mem[391] : 
                 (N1808)? mem[393] : 
                 (N1810)? mem[395] : 
                 (N1812)? mem[397] : 
                 (N1814)? mem[399] : 
                 (N1816)? mem[401] : 
                 (N1818)? mem[403] : 
                 (N1820)? mem[405] : 
                 (N1822)? mem[407] : 
                 (N1824)? mem[409] : 
                 (N1826)? mem[411] : 
                 (N1828)? mem[413] : 
                 (N1830)? mem[415] : 
                 (N1832)? mem[417] : 
                 (N1834)? mem[419] : 
                 (N1836)? mem[421] : 
                 (N1838)? mem[423] : 
                 (N1840)? mem[425] : 
                 (N1842)? mem[427] : 
                 (N1844)? mem[429] : 
                 (N1846)? mem[431] : 
                 (N1848)? mem[433] : 
                 (N1850)? mem[435] : 
                 (N1852)? mem[437] : 
                 (N1854)? mem[439] : 
                 (N1856)? mem[441] : 
                 (N1858)? mem[443] : 
                 (N1860)? mem[445] : 
                 (N1862)? mem[447] : 
                 (N1864)? mem[449] : 
                 (N1865)? mem[451] : 
                 (N1866)? mem[453] : 
                 (N1867)? mem[455] : 
                 (N1868)? mem[457] : 
                 (N1869)? mem[459] : 
                 (N1870)? mem[461] : 
                 (N1871)? mem[463] : 
                 (N1872)? mem[465] : 
                 (N1873)? mem[467] : 
                 (N1874)? mem[469] : 
                 (N1875)? mem[471] : 
                 (N1876)? mem[473] : 
                 (N1877)? mem[475] : 
                 (N1878)? mem[477] : 
                 (N1879)? mem[479] : 
                 (N1880)? mem[481] : 
                 (N1881)? mem[483] : 
                 (N1882)? mem[485] : 
                 (N1883)? mem[487] : 
                 (N1884)? mem[489] : 
                 (N1885)? mem[491] : 
                 (N1886)? mem[493] : 
                 (N1887)? mem[495] : 
                 (N1888)? mem[497] : 
                 (N1889)? mem[499] : 
                 (N1890)? mem[501] : 
                 (N1891)? mem[503] : 
                 (N1892)? mem[505] : 
                 (N1893)? mem[507] : 
                 (N1894)? mem[509] : 
                 (N1895)? mem[511] : 
                 (N1417)? mem[513] : 
                 (N1419)? mem[515] : 
                 (N1421)? mem[517] : 
                 (N1423)? mem[519] : 
                 (N1425)? mem[521] : 
                 (N1427)? mem[523] : 
                 (N1429)? mem[525] : 
                 (N1431)? mem[527] : 
                 (N1433)? mem[529] : 
                 (N1435)? mem[531] : 
                 (N1437)? mem[533] : 
                 (N1439)? mem[535] : 
                 (N1441)? mem[537] : 
                 (N1443)? mem[539] : 
                 (N1445)? mem[541] : 
                 (N1447)? mem[543] : 
                 (N1449)? mem[545] : 
                 (N1451)? mem[547] : 
                 (N1453)? mem[549] : 
                 (N1455)? mem[551] : 
                 (N1457)? mem[553] : 
                 (N1459)? mem[555] : 
                 (N1461)? mem[557] : 
                 (N1463)? mem[559] : 
                 (N1465)? mem[561] : 
                 (N1467)? mem[563] : 
                 (N1469)? mem[565] : 
                 (N1471)? mem[567] : 
                 (N1473)? mem[569] : 
                 (N1475)? mem[571] : 
                 (N1477)? mem[573] : 
                 (N1479)? mem[575] : 
                 (N1481)? mem[577] : 
                 (N1483)? mem[579] : 
                 (N1485)? mem[581] : 
                 (N1487)? mem[583] : 
                 (N1489)? mem[585] : 
                 (N1491)? mem[587] : 
                 (N1493)? mem[589] : 
                 (N1495)? mem[591] : 
                 (N1497)? mem[593] : 
                 (N1499)? mem[595] : 
                 (N1501)? mem[597] : 
                 (N1503)? mem[599] : 
                 (N1505)? mem[601] : 
                 (N1507)? mem[603] : 
                 (N1509)? mem[605] : 
                 (N1511)? mem[607] : 
                 (N1513)? mem[609] : 
                 (N1515)? mem[611] : 
                 (N1517)? mem[613] : 
                 (N1519)? mem[615] : 
                 (N1521)? mem[617] : 
                 (N1523)? mem[619] : 
                 (N1525)? mem[621] : 
                 (N1527)? mem[623] : 
                 (N1529)? mem[625] : 
                 (N1531)? mem[627] : 
                 (N1533)? mem[629] : 
                 (N1535)? mem[631] : 
                 (N1537)? mem[633] : 
                 (N1539)? mem[635] : 
                 (N1541)? mem[637] : 
                 (N1543)? mem[639] : 
                 (N1545)? mem[641] : 
                 (N1547)? mem[643] : 
                 (N1549)? mem[645] : 
                 (N1551)? mem[647] : 
                 (N1553)? mem[649] : 
                 (N1555)? mem[651] : 
                 (N1557)? mem[653] : 
                 (N1559)? mem[655] : 
                 (N1561)? mem[657] : 
                 (N1563)? mem[659] : 
                 (N1565)? mem[661] : 
                 (N1567)? mem[663] : 
                 (N1569)? mem[665] : 
                 (N1571)? mem[667] : 
                 (N1573)? mem[669] : 
                 (N1575)? mem[671] : 
                 (N1577)? mem[673] : 
                 (N1579)? mem[675] : 
                 (N1581)? mem[677] : 
                 (N1583)? mem[679] : 
                 (N1585)? mem[681] : 
                 (N1587)? mem[683] : 
                 (N1589)? mem[685] : 
                 (N1591)? mem[687] : 
                 (N1593)? mem[689] : 
                 (N1595)? mem[691] : 
                 (N1597)? mem[693] : 
                 (N1599)? mem[695] : 
                 (N1601)? mem[697] : 
                 (N1603)? mem[699] : 
                 (N1605)? mem[701] : 
                 (N1607)? mem[703] : 
                 (N1609)? mem[705] : 
                 (N1611)? mem[707] : 
                 (N1613)? mem[709] : 
                 (N1615)? mem[711] : 
                 (N1617)? mem[713] : 
                 (N1619)? mem[715] : 
                 (N1621)? mem[717] : 
                 (N1623)? mem[719] : 
                 (N1625)? mem[721] : 
                 (N1627)? mem[723] : 
                 (N1629)? mem[725] : 
                 (N1631)? mem[727] : 
                 (N1633)? mem[729] : 
                 (N1635)? mem[731] : 
                 (N1637)? mem[733] : 
                 (N1639)? mem[735] : 
                 (N1641)? mem[737] : 
                 (N1643)? mem[739] : 
                 (N1645)? mem[741] : 
                 (N1647)? mem[743] : 
                 (N1649)? mem[745] : 
                 (N1651)? mem[747] : 
                 (N1653)? mem[749] : 
                 (N1655)? mem[751] : 
                 (N1657)? mem[753] : 
                 (N1659)? mem[755] : 
                 (N1661)? mem[757] : 
                 (N1663)? mem[759] : 
                 (N1665)? mem[761] : 
                 (N1667)? mem[763] : 
                 (N1669)? mem[765] : 
                 (N1671)? mem[767] : 
                 (N1673)? mem[769] : 
                 (N1675)? mem[771] : 
                 (N1677)? mem[773] : 
                 (N1679)? mem[775] : 
                 (N1681)? mem[777] : 
                 (N1683)? mem[779] : 
                 (N1685)? mem[781] : 
                 (N1687)? mem[783] : 
                 (N1689)? mem[785] : 
                 (N1691)? mem[787] : 
                 (N1693)? mem[789] : 
                 (N1695)? mem[791] : 
                 (N1697)? mem[793] : 
                 (N1699)? mem[795] : 
                 (N1701)? mem[797] : 
                 (N1703)? mem[799] : 
                 (N1705)? mem[801] : 
                 (N1707)? mem[803] : 
                 (N1709)? mem[805] : 
                 (N1711)? mem[807] : 
                 (N1713)? mem[809] : 
                 (N1715)? mem[811] : 
                 (N1717)? mem[813] : 
                 (N1719)? mem[815] : 
                 (N1721)? mem[817] : 
                 (N1723)? mem[819] : 
                 (N1725)? mem[821] : 
                 (N1727)? mem[823] : 
                 (N1729)? mem[825] : 
                 (N1731)? mem[827] : 
                 (N1733)? mem[829] : 
                 (N1735)? mem[831] : 
                 (N1737)? mem[833] : 
                 (N1739)? mem[835] : 
                 (N1741)? mem[837] : 
                 (N1743)? mem[839] : 
                 (N1745)? mem[841] : 
                 (N1747)? mem[843] : 
                 (N1749)? mem[845] : 
                 (N1751)? mem[847] : 
                 (N1753)? mem[849] : 
                 (N1755)? mem[851] : 
                 (N1757)? mem[853] : 
                 (N1759)? mem[855] : 
                 (N1761)? mem[857] : 
                 (N1763)? mem[859] : 
                 (N1765)? mem[861] : 
                 (N1767)? mem[863] : 
                 (N1769)? mem[865] : 
                 (N1771)? mem[867] : 
                 (N1773)? mem[869] : 
                 (N1775)? mem[871] : 
                 (N1777)? mem[873] : 
                 (N1779)? mem[875] : 
                 (N1781)? mem[877] : 
                 (N1783)? mem[879] : 
                 (N1785)? mem[881] : 
                 (N1787)? mem[883] : 
                 (N1789)? mem[885] : 
                 (N1791)? mem[887] : 
                 (N1793)? mem[889] : 
                 (N1795)? mem[891] : 
                 (N1797)? mem[893] : 
                 (N1799)? mem[895] : 
                 (N1801)? mem[897] : 
                 (N1803)? mem[899] : 
                 (N1805)? mem[901] : 
                 (N1807)? mem[903] : 
                 (N1809)? mem[905] : 
                 (N1811)? mem[907] : 
                 (N1813)? mem[909] : 
                 (N1815)? mem[911] : 
                 (N1817)? mem[913] : 
                 (N1819)? mem[915] : 
                 (N1821)? mem[917] : 
                 (N1823)? mem[919] : 
                 (N1825)? mem[921] : 
                 (N1827)? mem[923] : 
                 (N1829)? mem[925] : 
                 (N1831)? mem[927] : 
                 (N1833)? mem[929] : 
                 (N1835)? mem[931] : 
                 (N1837)? mem[933] : 
                 (N1839)? mem[935] : 
                 (N1841)? mem[937] : 
                 (N1843)? mem[939] : 
                 (N1845)? mem[941] : 
                 (N1847)? mem[943] : 
                 (N1849)? mem[945] : 
                 (N1851)? mem[947] : 
                 (N1853)? mem[949] : 
                 (N1855)? mem[951] : 
                 (N1857)? mem[953] : 
                 (N1859)? mem[955] : 
                 (N1861)? mem[957] : 
                 (N1863)? mem[959] : 
                 (N4517)? mem[961] : 
                 (N4519)? mem[963] : 
                 (N4521)? mem[965] : 
                 (N4523)? mem[967] : 
                 (N4525)? mem[969] : 
                 (N4527)? mem[971] : 
                 (N4529)? mem[973] : 
                 (N4531)? mem[975] : 
                 (N4533)? mem[977] : 
                 (N4535)? mem[979] : 
                 (N4537)? mem[981] : 
                 (N4539)? mem[983] : 
                 (N4541)? mem[985] : 
                 (N4543)? mem[987] : 
                 (N4545)? mem[989] : 
                 (N4547)? mem[991] : 
                 (N3628)? mem[993] : 
                 (N3630)? mem[995] : 
                 (N3632)? mem[997] : 
                 (N3634)? mem[999] : 
                 (N3636)? mem[1001] : 
                 (N3638)? mem[1003] : 
                 (N3640)? mem[1005] : 
                 (N3642)? mem[1007] : 
                 (N12097)? mem[1009] : 
                 (N12099)? mem[1011] : 
                 (N12101)? mem[1013] : 
                 (N12103)? mem[1015] : 
                 (N12105)? mem[1017] : 
                 (N12107)? mem[1019] : 
                 (N12109)? mem[1021] : 
                 (N12111)? mem[1023] : 1'b0;
  assign N2665 = (N2201)? mem[0] : 
                 (N2203)? mem[2] : 
                 (N2205)? mem[4] : 
                 (N2207)? mem[6] : 
                 (N2209)? mem[8] : 
                 (N2211)? mem[10] : 
                 (N2213)? mem[12] : 
                 (N2215)? mem[14] : 
                 (N2217)? mem[16] : 
                 (N2219)? mem[18] : 
                 (N2221)? mem[20] : 
                 (N2223)? mem[22] : 
                 (N2225)? mem[24] : 
                 (N2227)? mem[26] : 
                 (N2229)? mem[28] : 
                 (N2231)? mem[30] : 
                 (N2233)? mem[32] : 
                 (N2235)? mem[34] : 
                 (N2237)? mem[36] : 
                 (N2239)? mem[38] : 
                 (N2241)? mem[40] : 
                 (N2243)? mem[42] : 
                 (N2245)? mem[44] : 
                 (N2247)? mem[46] : 
                 (N2249)? mem[48] : 
                 (N2251)? mem[50] : 
                 (N2253)? mem[52] : 
                 (N2255)? mem[54] : 
                 (N2257)? mem[56] : 
                 (N2259)? mem[58] : 
                 (N2261)? mem[60] : 
                 (N2263)? mem[62] : 
                 (N2265)? mem[64] : 
                 (N2267)? mem[66] : 
                 (N2269)? mem[68] : 
                 (N2271)? mem[70] : 
                 (N2273)? mem[72] : 
                 (N2275)? mem[74] : 
                 (N2277)? mem[76] : 
                 (N2279)? mem[78] : 
                 (N2281)? mem[80] : 
                 (N2283)? mem[82] : 
                 (N2285)? mem[84] : 
                 (N2287)? mem[86] : 
                 (N2289)? mem[88] : 
                 (N2291)? mem[90] : 
                 (N2293)? mem[92] : 
                 (N2295)? mem[94] : 
                 (N2297)? mem[96] : 
                 (N2299)? mem[98] : 
                 (N2301)? mem[100] : 
                 (N2303)? mem[102] : 
                 (N2305)? mem[104] : 
                 (N2307)? mem[106] : 
                 (N2309)? mem[108] : 
                 (N2311)? mem[110] : 
                 (N2313)? mem[112] : 
                 (N2315)? mem[114] : 
                 (N2317)? mem[116] : 
                 (N2319)? mem[118] : 
                 (N2321)? mem[120] : 
                 (N2323)? mem[122] : 
                 (N2325)? mem[124] : 
                 (N2327)? mem[126] : 
                 (N2329)? mem[128] : 
                 (N2331)? mem[130] : 
                 (N2333)? mem[132] : 
                 (N2335)? mem[134] : 
                 (N2337)? mem[136] : 
                 (N2339)? mem[138] : 
                 (N2341)? mem[140] : 
                 (N2343)? mem[142] : 
                 (N2345)? mem[144] : 
                 (N2347)? mem[146] : 
                 (N2349)? mem[148] : 
                 (N2351)? mem[150] : 
                 (N2353)? mem[152] : 
                 (N2355)? mem[154] : 
                 (N2357)? mem[156] : 
                 (N2359)? mem[158] : 
                 (N2361)? mem[160] : 
                 (N2363)? mem[162] : 
                 (N2365)? mem[164] : 
                 (N2367)? mem[166] : 
                 (N2369)? mem[168] : 
                 (N2371)? mem[170] : 
                 (N2373)? mem[172] : 
                 (N2375)? mem[174] : 
                 (N2377)? mem[176] : 
                 (N2379)? mem[178] : 
                 (N2381)? mem[180] : 
                 (N2383)? mem[182] : 
                 (N2385)? mem[184] : 
                 (N2387)? mem[186] : 
                 (N2389)? mem[188] : 
                 (N2391)? mem[190] : 
                 (N2393)? mem[192] : 
                 (N2395)? mem[194] : 
                 (N2397)? mem[196] : 
                 (N2399)? mem[198] : 
                 (N2401)? mem[200] : 
                 (N2403)? mem[202] : 
                 (N2405)? mem[204] : 
                 (N2407)? mem[206] : 
                 (N2409)? mem[208] : 
                 (N2411)? mem[210] : 
                 (N2413)? mem[212] : 
                 (N2415)? mem[214] : 
                 (N2417)? mem[216] : 
                 (N2419)? mem[218] : 
                 (N2421)? mem[220] : 
                 (N2423)? mem[222] : 
                 (N2425)? mem[224] : 
                 (N2427)? mem[226] : 
                 (N2429)? mem[228] : 
                 (N2431)? mem[230] : 
                 (N2433)? mem[232] : 
                 (N2435)? mem[234] : 
                 (N2437)? mem[236] : 
                 (N2439)? mem[238] : 
                 (N2441)? mem[240] : 
                 (N2443)? mem[242] : 
                 (N2445)? mem[244] : 
                 (N2447)? mem[246] : 
                 (N2449)? mem[248] : 
                 (N2451)? mem[250] : 
                 (N2453)? mem[252] : 
                 (N2455)? mem[254] : 
                 (N2457)? mem[256] : 
                 (N2459)? mem[258] : 
                 (N2461)? mem[260] : 
                 (N2463)? mem[262] : 
                 (N2465)? mem[264] : 
                 (N2467)? mem[266] : 
                 (N2469)? mem[268] : 
                 (N2471)? mem[270] : 
                 (N2473)? mem[272] : 
                 (N2475)? mem[274] : 
                 (N2477)? mem[276] : 
                 (N2479)? mem[278] : 
                 (N2481)? mem[280] : 
                 (N2483)? mem[282] : 
                 (N2485)? mem[284] : 
                 (N2487)? mem[286] : 
                 (N2489)? mem[288] : 
                 (N2491)? mem[290] : 
                 (N2493)? mem[292] : 
                 (N2495)? mem[294] : 
                 (N2497)? mem[296] : 
                 (N2499)? mem[298] : 
                 (N2501)? mem[300] : 
                 (N2503)? mem[302] : 
                 (N2505)? mem[304] : 
                 (N2507)? mem[306] : 
                 (N2509)? mem[308] : 
                 (N2511)? mem[310] : 
                 (N2513)? mem[312] : 
                 (N2515)? mem[314] : 
                 (N2517)? mem[316] : 
                 (N2519)? mem[318] : 
                 (N2521)? mem[320] : 
                 (N2523)? mem[322] : 
                 (N2525)? mem[324] : 
                 (N2527)? mem[326] : 
                 (N2529)? mem[328] : 
                 (N2531)? mem[330] : 
                 (N2533)? mem[332] : 
                 (N2535)? mem[334] : 
                 (N2537)? mem[336] : 
                 (N2539)? mem[338] : 
                 (N2541)? mem[340] : 
                 (N2543)? mem[342] : 
                 (N2545)? mem[344] : 
                 (N2547)? mem[346] : 
                 (N2549)? mem[348] : 
                 (N2551)? mem[350] : 
                 (N2553)? mem[352] : 
                 (N2555)? mem[354] : 
                 (N2557)? mem[356] : 
                 (N2559)? mem[358] : 
                 (N2561)? mem[360] : 
                 (N2563)? mem[362] : 
                 (N2565)? mem[364] : 
                 (N2567)? mem[366] : 
                 (N2569)? mem[368] : 
                 (N2571)? mem[370] : 
                 (N2573)? mem[372] : 
                 (N2575)? mem[374] : 
                 (N2577)? mem[376] : 
                 (N2579)? mem[378] : 
                 (N2581)? mem[380] : 
                 (N2583)? mem[382] : 
                 (N2585)? mem[384] : 
                 (N2587)? mem[386] : 
                 (N2589)? mem[388] : 
                 (N2591)? mem[390] : 
                 (N2593)? mem[392] : 
                 (N2595)? mem[394] : 
                 (N2597)? mem[396] : 
                 (N2599)? mem[398] : 
                 (N2601)? mem[400] : 
                 (N2602)? mem[402] : 
                 (N2603)? mem[404] : 
                 (N2604)? mem[406] : 
                 (N2605)? mem[408] : 
                 (N2606)? mem[410] : 
                 (N2607)? mem[412] : 
                 (N2608)? mem[414] : 
                 (N2609)? mem[416] : 
                 (N2611)? mem[418] : 
                 (N2613)? mem[420] : 
                 (N2615)? mem[422] : 
                 (N2617)? mem[424] : 
                 (N2619)? mem[426] : 
                 (N2621)? mem[428] : 
                 (N2623)? mem[430] : 
                 (N2625)? mem[432] : 
                 (N2626)? mem[434] : 
                 (N2627)? mem[436] : 
                 (N2628)? mem[438] : 
                 (N2629)? mem[440] : 
                 (N2630)? mem[442] : 
                 (N2631)? mem[444] : 
                 (N2632)? mem[446] : 
                 (N2633)? mem[448] : 
                 (N2634)? mem[450] : 
                 (N2635)? mem[452] : 
                 (N2636)? mem[454] : 
                 (N2637)? mem[456] : 
                 (N2638)? mem[458] : 
                 (N2639)? mem[460] : 
                 (N2640)? mem[462] : 
                 (N2641)? mem[464] : 
                 (N2642)? mem[466] : 
                 (N2643)? mem[468] : 
                 (N2644)? mem[470] : 
                 (N2645)? mem[472] : 
                 (N2646)? mem[474] : 
                 (N2647)? mem[476] : 
                 (N2648)? mem[478] : 
                 (N2649)? mem[480] : 
                 (N2650)? mem[482] : 
                 (N2651)? mem[484] : 
                 (N2652)? mem[486] : 
                 (N2653)? mem[488] : 
                 (N2654)? mem[490] : 
                 (N2655)? mem[492] : 
                 (N2656)? mem[494] : 
                 (N2657)? mem[496] : 
                 (N2658)? mem[498] : 
                 (N2659)? mem[500] : 
                 (N2660)? mem[502] : 
                 (N2661)? mem[504] : 
                 (N2662)? mem[506] : 
                 (N2663)? mem[508] : 
                 (N2664)? mem[510] : 
                 (N2202)? mem[512] : 
                 (N2204)? mem[514] : 
                 (N2206)? mem[516] : 
                 (N2208)? mem[518] : 
                 (N2210)? mem[520] : 
                 (N2212)? mem[522] : 
                 (N2214)? mem[524] : 
                 (N2216)? mem[526] : 
                 (N2218)? mem[528] : 
                 (N2220)? mem[530] : 
                 (N2222)? mem[532] : 
                 (N2224)? mem[534] : 
                 (N2226)? mem[536] : 
                 (N2228)? mem[538] : 
                 (N2230)? mem[540] : 
                 (N2232)? mem[542] : 
                 (N2234)? mem[544] : 
                 (N2236)? mem[546] : 
                 (N2238)? mem[548] : 
                 (N2240)? mem[550] : 
                 (N2242)? mem[552] : 
                 (N2244)? mem[554] : 
                 (N2246)? mem[556] : 
                 (N2248)? mem[558] : 
                 (N2250)? mem[560] : 
                 (N2252)? mem[562] : 
                 (N2254)? mem[564] : 
                 (N2256)? mem[566] : 
                 (N2258)? mem[568] : 
                 (N2260)? mem[570] : 
                 (N2262)? mem[572] : 
                 (N2264)? mem[574] : 
                 (N2266)? mem[576] : 
                 (N2268)? mem[578] : 
                 (N2270)? mem[580] : 
                 (N2272)? mem[582] : 
                 (N2274)? mem[584] : 
                 (N2276)? mem[586] : 
                 (N2278)? mem[588] : 
                 (N2280)? mem[590] : 
                 (N2282)? mem[592] : 
                 (N2284)? mem[594] : 
                 (N2286)? mem[596] : 
                 (N2288)? mem[598] : 
                 (N2290)? mem[600] : 
                 (N2292)? mem[602] : 
                 (N2294)? mem[604] : 
                 (N2296)? mem[606] : 
                 (N2298)? mem[608] : 
                 (N2300)? mem[610] : 
                 (N2302)? mem[612] : 
                 (N2304)? mem[614] : 
                 (N2306)? mem[616] : 
                 (N2308)? mem[618] : 
                 (N2310)? mem[620] : 
                 (N2312)? mem[622] : 
                 (N2314)? mem[624] : 
                 (N2316)? mem[626] : 
                 (N2318)? mem[628] : 
                 (N2320)? mem[630] : 
                 (N2322)? mem[632] : 
                 (N2324)? mem[634] : 
                 (N2326)? mem[636] : 
                 (N2328)? mem[638] : 
                 (N2330)? mem[640] : 
                 (N2332)? mem[642] : 
                 (N2334)? mem[644] : 
                 (N2336)? mem[646] : 
                 (N2338)? mem[648] : 
                 (N2340)? mem[650] : 
                 (N2342)? mem[652] : 
                 (N2344)? mem[654] : 
                 (N2346)? mem[656] : 
                 (N2348)? mem[658] : 
                 (N2350)? mem[660] : 
                 (N2352)? mem[662] : 
                 (N2354)? mem[664] : 
                 (N2356)? mem[666] : 
                 (N2358)? mem[668] : 
                 (N2360)? mem[670] : 
                 (N2362)? mem[672] : 
                 (N2364)? mem[674] : 
                 (N2366)? mem[676] : 
                 (N2368)? mem[678] : 
                 (N2370)? mem[680] : 
                 (N2372)? mem[682] : 
                 (N2374)? mem[684] : 
                 (N2376)? mem[686] : 
                 (N2378)? mem[688] : 
                 (N2380)? mem[690] : 
                 (N2382)? mem[692] : 
                 (N2384)? mem[694] : 
                 (N2386)? mem[696] : 
                 (N2388)? mem[698] : 
                 (N2390)? mem[700] : 
                 (N2392)? mem[702] : 
                 (N2394)? mem[704] : 
                 (N2396)? mem[706] : 
                 (N2398)? mem[708] : 
                 (N2400)? mem[710] : 
                 (N2402)? mem[712] : 
                 (N2404)? mem[714] : 
                 (N2406)? mem[716] : 
                 (N2408)? mem[718] : 
                 (N2410)? mem[720] : 
                 (N2412)? mem[722] : 
                 (N2414)? mem[724] : 
                 (N2416)? mem[726] : 
                 (N2418)? mem[728] : 
                 (N2420)? mem[730] : 
                 (N2422)? mem[732] : 
                 (N2424)? mem[734] : 
                 (N2426)? mem[736] : 
                 (N2428)? mem[738] : 
                 (N2430)? mem[740] : 
                 (N2432)? mem[742] : 
                 (N2434)? mem[744] : 
                 (N2436)? mem[746] : 
                 (N2438)? mem[748] : 
                 (N2440)? mem[750] : 
                 (N2442)? mem[752] : 
                 (N2444)? mem[754] : 
                 (N2446)? mem[756] : 
                 (N2448)? mem[758] : 
                 (N2450)? mem[760] : 
                 (N2452)? mem[762] : 
                 (N2454)? mem[764] : 
                 (N2456)? mem[766] : 
                 (N2458)? mem[768] : 
                 (N2460)? mem[770] : 
                 (N2462)? mem[772] : 
                 (N2464)? mem[774] : 
                 (N2466)? mem[776] : 
                 (N2468)? mem[778] : 
                 (N2470)? mem[780] : 
                 (N2472)? mem[782] : 
                 (N2474)? mem[784] : 
                 (N2476)? mem[786] : 
                 (N2478)? mem[788] : 
                 (N2480)? mem[790] : 
                 (N2482)? mem[792] : 
                 (N2484)? mem[794] : 
                 (N2486)? mem[796] : 
                 (N2488)? mem[798] : 
                 (N2490)? mem[800] : 
                 (N2492)? mem[802] : 
                 (N2494)? mem[804] : 
                 (N2496)? mem[806] : 
                 (N2498)? mem[808] : 
                 (N2500)? mem[810] : 
                 (N2502)? mem[812] : 
                 (N2504)? mem[814] : 
                 (N2506)? mem[816] : 
                 (N2508)? mem[818] : 
                 (N2510)? mem[820] : 
                 (N2512)? mem[822] : 
                 (N2514)? mem[824] : 
                 (N2516)? mem[826] : 
                 (N2518)? mem[828] : 
                 (N2520)? mem[830] : 
                 (N2522)? mem[832] : 
                 (N2524)? mem[834] : 
                 (N2526)? mem[836] : 
                 (N2528)? mem[838] : 
                 (N2530)? mem[840] : 
                 (N2532)? mem[842] : 
                 (N2534)? mem[844] : 
                 (N2536)? mem[846] : 
                 (N2538)? mem[848] : 
                 (N2540)? mem[850] : 
                 (N2542)? mem[852] : 
                 (N2544)? mem[854] : 
                 (N2546)? mem[856] : 
                 (N2548)? mem[858] : 
                 (N2550)? mem[860] : 
                 (N2552)? mem[862] : 
                 (N2554)? mem[864] : 
                 (N2556)? mem[866] : 
                 (N2558)? mem[868] : 
                 (N2560)? mem[870] : 
                 (N2562)? mem[872] : 
                 (N2564)? mem[874] : 
                 (N2566)? mem[876] : 
                 (N2568)? mem[878] : 
                 (N2570)? mem[880] : 
                 (N2572)? mem[882] : 
                 (N2574)? mem[884] : 
                 (N2576)? mem[886] : 
                 (N2578)? mem[888] : 
                 (N2580)? mem[890] : 
                 (N2582)? mem[892] : 
                 (N2584)? mem[894] : 
                 (N2586)? mem[896] : 
                 (N2588)? mem[898] : 
                 (N2590)? mem[900] : 
                 (N2592)? mem[902] : 
                 (N2594)? mem[904] : 
                 (N2596)? mem[906] : 
                 (N2598)? mem[908] : 
                 (N2600)? mem[910] : 
                 (N5863)? mem[912] : 
                 (N5865)? mem[914] : 
                 (N5867)? mem[916] : 
                 (N5869)? mem[918] : 
                 (N5871)? mem[920] : 
                 (N5873)? mem[922] : 
                 (N5875)? mem[924] : 
                 (N5877)? mem[926] : 
                 (N2610)? mem[928] : 
                 (N2612)? mem[930] : 
                 (N2614)? mem[932] : 
                 (N2616)? mem[934] : 
                 (N2618)? mem[936] : 
                 (N2620)? mem[938] : 
                 (N2622)? mem[940] : 
                 (N2624)? mem[942] : 
                 (N5895)? mem[944] : 
                 (N5897)? mem[946] : 
                 (N5899)? mem[948] : 
                 (N5901)? mem[950] : 
                 (N5903)? mem[952] : 
                 (N5905)? mem[954] : 
                 (N5907)? mem[956] : 
                 (N5909)? mem[958] : 
                 (N4517)? mem[960] : 
                 (N4519)? mem[962] : 
                 (N4521)? mem[964] : 
                 (N4523)? mem[966] : 
                 (N4525)? mem[968] : 
                 (N4527)? mem[970] : 
                 (N4529)? mem[972] : 
                 (N4531)? mem[974] : 
                 (N4533)? mem[976] : 
                 (N4535)? mem[978] : 
                 (N4537)? mem[980] : 
                 (N4539)? mem[982] : 
                 (N4541)? mem[984] : 
                 (N4543)? mem[986] : 
                 (N4545)? mem[988] : 
                 (N4547)? mem[990] : 
                 (N3628)? mem[992] : 
                 (N3630)? mem[994] : 
                 (N3632)? mem[996] : 
                 (N3634)? mem[998] : 
                 (N3636)? mem[1000] : 
                 (N3638)? mem[1002] : 
                 (N3640)? mem[1004] : 
                 (N3642)? mem[1006] : 
                 (N12097)? mem[1008] : 
                 (N12099)? mem[1010] : 
                 (N12101)? mem[1012] : 
                 (N12103)? mem[1014] : 
                 (N12105)? mem[1016] : 
                 (N12107)? mem[1018] : 
                 (N12109)? mem[1020] : 
                 (N12111)? mem[1022] : 1'b0;
  assign N2669 = N2666 & N2667;
  assign N2670 = N2669 & N2668;
  assign N2671 = correct_i | N1896;
  assign N2672 = N2671 | N2668;
  assign N2674 = correct_i | N2667;
  assign N2675 = N2674 | N2665;
  assign N2677 = N2674 | N2668;
  assign N2679 = N2666 | N1896;
  assign N2680 = N2679 | N2665;
  assign N2682 = N2679 | N2668;
  assign N2684 = N2666 | N2667;
  assign N2685 = N2684 | N2665;
  assign N2687 = correct_i & N1896;
  assign N2688 = N2687 & N2665;
  assign N3651 = (N3147)? mem[1] : 
                 (N3149)? mem[3] : 
                 (N3151)? mem[5] : 
                 (N3153)? mem[7] : 
                 (N3155)? mem[9] : 
                 (N3157)? mem[11] : 
                 (N3159)? mem[13] : 
                 (N3161)? mem[15] : 
                 (N3163)? mem[17] : 
                 (N3165)? mem[19] : 
                 (N3167)? mem[21] : 
                 (N3169)? mem[23] : 
                 (N3171)? mem[25] : 
                 (N3173)? mem[27] : 
                 (N3175)? mem[29] : 
                 (N3177)? mem[31] : 
                 (N3179)? mem[33] : 
                 (N3181)? mem[35] : 
                 (N3183)? mem[37] : 
                 (N3185)? mem[39] : 
                 (N3187)? mem[41] : 
                 (N3189)? mem[43] : 
                 (N3191)? mem[45] : 
                 (N3193)? mem[47] : 
                 (N3195)? mem[49] : 
                 (N3197)? mem[51] : 
                 (N3199)? mem[53] : 
                 (N3201)? mem[55] : 
                 (N3203)? mem[57] : 
                 (N3205)? mem[59] : 
                 (N3207)? mem[61] : 
                 (N3209)? mem[63] : 
                 (N3211)? mem[65] : 
                 (N3213)? mem[67] : 
                 (N3215)? mem[69] : 
                 (N3217)? mem[71] : 
                 (N3219)? mem[73] : 
                 (N3221)? mem[75] : 
                 (N3223)? mem[77] : 
                 (N3225)? mem[79] : 
                 (N3227)? mem[81] : 
                 (N3229)? mem[83] : 
                 (N3231)? mem[85] : 
                 (N3233)? mem[87] : 
                 (N3235)? mem[89] : 
                 (N3237)? mem[91] : 
                 (N3239)? mem[93] : 
                 (N3241)? mem[95] : 
                 (N3243)? mem[97] : 
                 (N3245)? mem[99] : 
                 (N3247)? mem[101] : 
                 (N3249)? mem[103] : 
                 (N3251)? mem[105] : 
                 (N3253)? mem[107] : 
                 (N3255)? mem[109] : 
                 (N3257)? mem[111] : 
                 (N3259)? mem[113] : 
                 (N3261)? mem[115] : 
                 (N3263)? mem[117] : 
                 (N3265)? mem[119] : 
                 (N3267)? mem[121] : 
                 (N3269)? mem[123] : 
                 (N3271)? mem[125] : 
                 (N3273)? mem[127] : 
                 (N3275)? mem[129] : 
                 (N3277)? mem[131] : 
                 (N3279)? mem[133] : 
                 (N3281)? mem[135] : 
                 (N3283)? mem[137] : 
                 (N3285)? mem[139] : 
                 (N3287)? mem[141] : 
                 (N3289)? mem[143] : 
                 (N3291)? mem[145] : 
                 (N3293)? mem[147] : 
                 (N3295)? mem[149] : 
                 (N3297)? mem[151] : 
                 (N3299)? mem[153] : 
                 (N3301)? mem[155] : 
                 (N3303)? mem[157] : 
                 (N3305)? mem[159] : 
                 (N3307)? mem[161] : 
                 (N3309)? mem[163] : 
                 (N3311)? mem[165] : 
                 (N3313)? mem[167] : 
                 (N3315)? mem[169] : 
                 (N3317)? mem[171] : 
                 (N3319)? mem[173] : 
                 (N3321)? mem[175] : 
                 (N3323)? mem[177] : 
                 (N3325)? mem[179] : 
                 (N3327)? mem[181] : 
                 (N3329)? mem[183] : 
                 (N3331)? mem[185] : 
                 (N3333)? mem[187] : 
                 (N3335)? mem[189] : 
                 (N3337)? mem[191] : 
                 (N3339)? mem[193] : 
                 (N3341)? mem[195] : 
                 (N3343)? mem[197] : 
                 (N3345)? mem[199] : 
                 (N3347)? mem[201] : 
                 (N3349)? mem[203] : 
                 (N3351)? mem[205] : 
                 (N3353)? mem[207] : 
                 (N3355)? mem[209] : 
                 (N3357)? mem[211] : 
                 (N3359)? mem[213] : 
                 (N3361)? mem[215] : 
                 (N3363)? mem[217] : 
                 (N3365)? mem[219] : 
                 (N3367)? mem[221] : 
                 (N3369)? mem[223] : 
                 (N3371)? mem[225] : 
                 (N3373)? mem[227] : 
                 (N3375)? mem[229] : 
                 (N3377)? mem[231] : 
                 (N3379)? mem[233] : 
                 (N3381)? mem[235] : 
                 (N3383)? mem[237] : 
                 (N3385)? mem[239] : 
                 (N3387)? mem[241] : 
                 (N3389)? mem[243] : 
                 (N3391)? mem[245] : 
                 (N3393)? mem[247] : 
                 (N3395)? mem[249] : 
                 (N3397)? mem[251] : 
                 (N3399)? mem[253] : 
                 (N3401)? mem[255] : 
                 (N3403)? mem[257] : 
                 (N3405)? mem[259] : 
                 (N3407)? mem[261] : 
                 (N3409)? mem[263] : 
                 (N3411)? mem[265] : 
                 (N3413)? mem[267] : 
                 (N3415)? mem[269] : 
                 (N3417)? mem[271] : 
                 (N3419)? mem[273] : 
                 (N3421)? mem[275] : 
                 (N3423)? mem[277] : 
                 (N3425)? mem[279] : 
                 (N3427)? mem[281] : 
                 (N3429)? mem[283] : 
                 (N3431)? mem[285] : 
                 (N3433)? mem[287] : 
                 (N3435)? mem[289] : 
                 (N3437)? mem[291] : 
                 (N3439)? mem[293] : 
                 (N3441)? mem[295] : 
                 (N3443)? mem[297] : 
                 (N3445)? mem[299] : 
                 (N3447)? mem[301] : 
                 (N3449)? mem[303] : 
                 (N3451)? mem[305] : 
                 (N3453)? mem[307] : 
                 (N3455)? mem[309] : 
                 (N3457)? mem[311] : 
                 (N3459)? mem[313] : 
                 (N3461)? mem[315] : 
                 (N3463)? mem[317] : 
                 (N3465)? mem[319] : 
                 (N3467)? mem[321] : 
                 (N3469)? mem[323] : 
                 (N3471)? mem[325] : 
                 (N3473)? mem[327] : 
                 (N3475)? mem[329] : 
                 (N3477)? mem[331] : 
                 (N3479)? mem[333] : 
                 (N3481)? mem[335] : 
                 (N3483)? mem[337] : 
                 (N3485)? mem[339] : 
                 (N3487)? mem[341] : 
                 (N3489)? mem[343] : 
                 (N3491)? mem[345] : 
                 (N3493)? mem[347] : 
                 (N3495)? mem[349] : 
                 (N3497)? mem[351] : 
                 (N3499)? mem[353] : 
                 (N3501)? mem[355] : 
                 (N3503)? mem[357] : 
                 (N3505)? mem[359] : 
                 (N3507)? mem[361] : 
                 (N3509)? mem[363] : 
                 (N3511)? mem[365] : 
                 (N3513)? mem[367] : 
                 (N3515)? mem[369] : 
                 (N3517)? mem[371] : 
                 (N3519)? mem[373] : 
                 (N3521)? mem[375] : 
                 (N3523)? mem[377] : 
                 (N3525)? mem[379] : 
                 (N3527)? mem[381] : 
                 (N3529)? mem[383] : 
                 (N3531)? mem[385] : 
                 (N3533)? mem[387] : 
                 (N3535)? mem[389] : 
                 (N3537)? mem[391] : 
                 (N3539)? mem[393] : 
                 (N3541)? mem[395] : 
                 (N3543)? mem[397] : 
                 (N3545)? mem[399] : 
                 (N3547)? mem[401] : 
                 (N3549)? mem[403] : 
                 (N3551)? mem[405] : 
                 (N3553)? mem[407] : 
                 (N3555)? mem[409] : 
                 (N3557)? mem[411] : 
                 (N3559)? mem[413] : 
                 (N3561)? mem[415] : 
                 (N3563)? mem[417] : 
                 (N3565)? mem[419] : 
                 (N3567)? mem[421] : 
                 (N3569)? mem[423] : 
                 (N3571)? mem[425] : 
                 (N3573)? mem[427] : 
                 (N3575)? mem[429] : 
                 (N3577)? mem[431] : 
                 (N3579)? mem[433] : 
                 (N3581)? mem[435] : 
                 (N3583)? mem[437] : 
                 (N3585)? mem[439] : 
                 (N3587)? mem[441] : 
                 (N3589)? mem[443] : 
                 (N3591)? mem[445] : 
                 (N3593)? mem[447] : 
                 (N3595)? mem[449] : 
                 (N3597)? mem[451] : 
                 (N3599)? mem[453] : 
                 (N3601)? mem[455] : 
                 (N3603)? mem[457] : 
                 (N3605)? mem[459] : 
                 (N3607)? mem[461] : 
                 (N3609)? mem[463] : 
                 (N3611)? mem[465] : 
                 (N3613)? mem[467] : 
                 (N3615)? mem[469] : 
                 (N3617)? mem[471] : 
                 (N3619)? mem[473] : 
                 (N3621)? mem[475] : 
                 (N3623)? mem[477] : 
                 (N3625)? mem[479] : 
                 (N3627)? mem[481] : 
                 (N3629)? mem[483] : 
                 (N3631)? mem[485] : 
                 (N3633)? mem[487] : 
                 (N3635)? mem[489] : 
                 (N3637)? mem[491] : 
                 (N3639)? mem[493] : 
                 (N3641)? mem[495] : 
                 (N3643)? mem[497] : 
                 (N3644)? mem[499] : 
                 (N3645)? mem[501] : 
                 (N3646)? mem[503] : 
                 (N3647)? mem[505] : 
                 (N3648)? mem[507] : 
                 (N3649)? mem[509] : 
                 (N3650)? mem[511] : 
                 (N3148)? mem[513] : 
                 (N3150)? mem[515] : 
                 (N3152)? mem[517] : 
                 (N3154)? mem[519] : 
                 (N3156)? mem[521] : 
                 (N3158)? mem[523] : 
                 (N3160)? mem[525] : 
                 (N3162)? mem[527] : 
                 (N3164)? mem[529] : 
                 (N3166)? mem[531] : 
                 (N3168)? mem[533] : 
                 (N3170)? mem[535] : 
                 (N3172)? mem[537] : 
                 (N3174)? mem[539] : 
                 (N3176)? mem[541] : 
                 (N3178)? mem[543] : 
                 (N3180)? mem[545] : 
                 (N3182)? mem[547] : 
                 (N3184)? mem[549] : 
                 (N3186)? mem[551] : 
                 (N3188)? mem[553] : 
                 (N3190)? mem[555] : 
                 (N3192)? mem[557] : 
                 (N3194)? mem[559] : 
                 (N3196)? mem[561] : 
                 (N3198)? mem[563] : 
                 (N3200)? mem[565] : 
                 (N3202)? mem[567] : 
                 (N3204)? mem[569] : 
                 (N3206)? mem[571] : 
                 (N3208)? mem[573] : 
                 (N3210)? mem[575] : 
                 (N3212)? mem[577] : 
                 (N3214)? mem[579] : 
                 (N3216)? mem[581] : 
                 (N3218)? mem[583] : 
                 (N3220)? mem[585] : 
                 (N3222)? mem[587] : 
                 (N3224)? mem[589] : 
                 (N3226)? mem[591] : 
                 (N3228)? mem[593] : 
                 (N3230)? mem[595] : 
                 (N3232)? mem[597] : 
                 (N3234)? mem[599] : 
                 (N3236)? mem[601] : 
                 (N3238)? mem[603] : 
                 (N3240)? mem[605] : 
                 (N3242)? mem[607] : 
                 (N3244)? mem[609] : 
                 (N3246)? mem[611] : 
                 (N3248)? mem[613] : 
                 (N3250)? mem[615] : 
                 (N3252)? mem[617] : 
                 (N3254)? mem[619] : 
                 (N3256)? mem[621] : 
                 (N3258)? mem[623] : 
                 (N3260)? mem[625] : 
                 (N3262)? mem[627] : 
                 (N3264)? mem[629] : 
                 (N3266)? mem[631] : 
                 (N3268)? mem[633] : 
                 (N3270)? mem[635] : 
                 (N3272)? mem[637] : 
                 (N3274)? mem[639] : 
                 (N3276)? mem[641] : 
                 (N3278)? mem[643] : 
                 (N3280)? mem[645] : 
                 (N3282)? mem[647] : 
                 (N3284)? mem[649] : 
                 (N3286)? mem[651] : 
                 (N3288)? mem[653] : 
                 (N3290)? mem[655] : 
                 (N3292)? mem[657] : 
                 (N3294)? mem[659] : 
                 (N3296)? mem[661] : 
                 (N3298)? mem[663] : 
                 (N3300)? mem[665] : 
                 (N3302)? mem[667] : 
                 (N3304)? mem[669] : 
                 (N3306)? mem[671] : 
                 (N3308)? mem[673] : 
                 (N3310)? mem[675] : 
                 (N3312)? mem[677] : 
                 (N3314)? mem[679] : 
                 (N3316)? mem[681] : 
                 (N3318)? mem[683] : 
                 (N3320)? mem[685] : 
                 (N3322)? mem[687] : 
                 (N3324)? mem[689] : 
                 (N3326)? mem[691] : 
                 (N3328)? mem[693] : 
                 (N3330)? mem[695] : 
                 (N3332)? mem[697] : 
                 (N3334)? mem[699] : 
                 (N3336)? mem[701] : 
                 (N3338)? mem[703] : 
                 (N3340)? mem[705] : 
                 (N3342)? mem[707] : 
                 (N3344)? mem[709] : 
                 (N3346)? mem[711] : 
                 (N3348)? mem[713] : 
                 (N3350)? mem[715] : 
                 (N3352)? mem[717] : 
                 (N3354)? mem[719] : 
                 (N3356)? mem[721] : 
                 (N3358)? mem[723] : 
                 (N3360)? mem[725] : 
                 (N3362)? mem[727] : 
                 (N3364)? mem[729] : 
                 (N3366)? mem[731] : 
                 (N3368)? mem[733] : 
                 (N3370)? mem[735] : 
                 (N3372)? mem[737] : 
                 (N3374)? mem[739] : 
                 (N3376)? mem[741] : 
                 (N3378)? mem[743] : 
                 (N3380)? mem[745] : 
                 (N3382)? mem[747] : 
                 (N3384)? mem[749] : 
                 (N3386)? mem[751] : 
                 (N3388)? mem[753] : 
                 (N3390)? mem[755] : 
                 (N3392)? mem[757] : 
                 (N3394)? mem[759] : 
                 (N3396)? mem[761] : 
                 (N3398)? mem[763] : 
                 (N3400)? mem[765] : 
                 (N3402)? mem[767] : 
                 (N3404)? mem[769] : 
                 (N3406)? mem[771] : 
                 (N3408)? mem[773] : 
                 (N3410)? mem[775] : 
                 (N3412)? mem[777] : 
                 (N3414)? mem[779] : 
                 (N3416)? mem[781] : 
                 (N3418)? mem[783] : 
                 (N3420)? mem[785] : 
                 (N3422)? mem[787] : 
                 (N3424)? mem[789] : 
                 (N3426)? mem[791] : 
                 (N3428)? mem[793] : 
                 (N3430)? mem[795] : 
                 (N3432)? mem[797] : 
                 (N3434)? mem[799] : 
                 (N3436)? mem[801] : 
                 (N3438)? mem[803] : 
                 (N3440)? mem[805] : 
                 (N3442)? mem[807] : 
                 (N3444)? mem[809] : 
                 (N3446)? mem[811] : 
                 (N3448)? mem[813] : 
                 (N3450)? mem[815] : 
                 (N3452)? mem[817] : 
                 (N3454)? mem[819] : 
                 (N3456)? mem[821] : 
                 (N3458)? mem[823] : 
                 (N3460)? mem[825] : 
                 (N3462)? mem[827] : 
                 (N3464)? mem[829] : 
                 (N3466)? mem[831] : 
                 (N3468)? mem[833] : 
                 (N3470)? mem[835] : 
                 (N3472)? mem[837] : 
                 (N3474)? mem[839] : 
                 (N3476)? mem[841] : 
                 (N3478)? mem[843] : 
                 (N3480)? mem[845] : 
                 (N3482)? mem[847] : 
                 (N3484)? mem[849] : 
                 (N3486)? mem[851] : 
                 (N3488)? mem[853] : 
                 (N3490)? mem[855] : 
                 (N3492)? mem[857] : 
                 (N3494)? mem[859] : 
                 (N3496)? mem[861] : 
                 (N3498)? mem[863] : 
                 (N3500)? mem[865] : 
                 (N3502)? mem[867] : 
                 (N3504)? mem[869] : 
                 (N3506)? mem[871] : 
                 (N3508)? mem[873] : 
                 (N3510)? mem[875] : 
                 (N3512)? mem[877] : 
                 (N3514)? mem[879] : 
                 (N3516)? mem[881] : 
                 (N3518)? mem[883] : 
                 (N3520)? mem[885] : 
                 (N3522)? mem[887] : 
                 (N3524)? mem[889] : 
                 (N3526)? mem[891] : 
                 (N3528)? mem[893] : 
                 (N3530)? mem[895] : 
                 (N3532)? mem[897] : 
                 (N3534)? mem[899] : 
                 (N3536)? mem[901] : 
                 (N3538)? mem[903] : 
                 (N3540)? mem[905] : 
                 (N3542)? mem[907] : 
                 (N3544)? mem[909] : 
                 (N3546)? mem[911] : 
                 (N3548)? mem[913] : 
                 (N3550)? mem[915] : 
                 (N3552)? mem[917] : 
                 (N3554)? mem[919] : 
                 (N3556)? mem[921] : 
                 (N3558)? mem[923] : 
                 (N3560)? mem[925] : 
                 (N3562)? mem[927] : 
                 (N3564)? mem[929] : 
                 (N3566)? mem[931] : 
                 (N3568)? mem[933] : 
                 (N3570)? mem[935] : 
                 (N3572)? mem[937] : 
                 (N3574)? mem[939] : 
                 (N3576)? mem[941] : 
                 (N3578)? mem[943] : 
                 (N3580)? mem[945] : 
                 (N3582)? mem[947] : 
                 (N3584)? mem[949] : 
                 (N3586)? mem[951] : 
                 (N3588)? mem[953] : 
                 (N3590)? mem[955] : 
                 (N3592)? mem[957] : 
                 (N3594)? mem[959] : 
                 (N3596)? mem[961] : 
                 (N3598)? mem[963] : 
                 (N3600)? mem[965] : 
                 (N3602)? mem[967] : 
                 (N3604)? mem[969] : 
                 (N3606)? mem[971] : 
                 (N3608)? mem[973] : 
                 (N3610)? mem[975] : 
                 (N3612)? mem[977] : 
                 (N3614)? mem[979] : 
                 (N3616)? mem[981] : 
                 (N3618)? mem[983] : 
                 (N3620)? mem[985] : 
                 (N3622)? mem[987] : 
                 (N3624)? mem[989] : 
                 (N3626)? mem[991] : 
                 (N3628)? mem[993] : 
                 (N3630)? mem[995] : 
                 (N3632)? mem[997] : 
                 (N3634)? mem[999] : 
                 (N3636)? mem[1001] : 
                 (N3638)? mem[1003] : 
                 (N3640)? mem[1005] : 
                 (N3642)? mem[1007] : 
                 (N12097)? mem[1009] : 
                 (N12099)? mem[1011] : 
                 (N12101)? mem[1013] : 
                 (N12103)? mem[1015] : 
                 (N12105)? mem[1017] : 
                 (N12107)? mem[1019] : 
                 (N12109)? mem[1021] : 
                 (N12111)? mem[1023] : 1'b0;
  assign N4564 = (N4068)? mem[0] : 
                 (N4070)? mem[2] : 
                 (N4072)? mem[4] : 
                 (N4074)? mem[6] : 
                 (N4076)? mem[8] : 
                 (N4078)? mem[10] : 
                 (N4080)? mem[12] : 
                 (N4082)? mem[14] : 
                 (N4084)? mem[16] : 
                 (N4086)? mem[18] : 
                 (N4088)? mem[20] : 
                 (N4090)? mem[22] : 
                 (N4092)? mem[24] : 
                 (N4094)? mem[26] : 
                 (N4096)? mem[28] : 
                 (N4098)? mem[30] : 
                 (N4100)? mem[32] : 
                 (N4102)? mem[34] : 
                 (N4104)? mem[36] : 
                 (N4106)? mem[38] : 
                 (N4108)? mem[40] : 
                 (N4110)? mem[42] : 
                 (N4112)? mem[44] : 
                 (N4114)? mem[46] : 
                 (N4116)? mem[48] : 
                 (N4118)? mem[50] : 
                 (N4120)? mem[52] : 
                 (N4122)? mem[54] : 
                 (N4124)? mem[56] : 
                 (N4126)? mem[58] : 
                 (N4128)? mem[60] : 
                 (N4130)? mem[62] : 
                 (N4132)? mem[64] : 
                 (N4134)? mem[66] : 
                 (N4136)? mem[68] : 
                 (N4138)? mem[70] : 
                 (N4140)? mem[72] : 
                 (N4142)? mem[74] : 
                 (N4144)? mem[76] : 
                 (N4146)? mem[78] : 
                 (N4148)? mem[80] : 
                 (N4150)? mem[82] : 
                 (N4152)? mem[84] : 
                 (N4154)? mem[86] : 
                 (N4156)? mem[88] : 
                 (N4158)? mem[90] : 
                 (N4160)? mem[92] : 
                 (N4162)? mem[94] : 
                 (N4164)? mem[96] : 
                 (N4166)? mem[98] : 
                 (N4168)? mem[100] : 
                 (N4170)? mem[102] : 
                 (N4172)? mem[104] : 
                 (N4174)? mem[106] : 
                 (N4176)? mem[108] : 
                 (N4178)? mem[110] : 
                 (N4180)? mem[112] : 
                 (N4182)? mem[114] : 
                 (N4184)? mem[116] : 
                 (N4186)? mem[118] : 
                 (N4188)? mem[120] : 
                 (N4190)? mem[122] : 
                 (N4192)? mem[124] : 
                 (N4194)? mem[126] : 
                 (N4196)? mem[128] : 
                 (N4198)? mem[130] : 
                 (N4200)? mem[132] : 
                 (N4202)? mem[134] : 
                 (N4204)? mem[136] : 
                 (N4206)? mem[138] : 
                 (N4208)? mem[140] : 
                 (N4210)? mem[142] : 
                 (N4212)? mem[144] : 
                 (N4214)? mem[146] : 
                 (N4216)? mem[148] : 
                 (N4218)? mem[150] : 
                 (N4220)? mem[152] : 
                 (N4222)? mem[154] : 
                 (N4224)? mem[156] : 
                 (N4226)? mem[158] : 
                 (N4228)? mem[160] : 
                 (N4230)? mem[162] : 
                 (N4232)? mem[164] : 
                 (N4234)? mem[166] : 
                 (N4236)? mem[168] : 
                 (N4238)? mem[170] : 
                 (N4240)? mem[172] : 
                 (N4242)? mem[174] : 
                 (N4244)? mem[176] : 
                 (N4246)? mem[178] : 
                 (N4248)? mem[180] : 
                 (N4250)? mem[182] : 
                 (N4252)? mem[184] : 
                 (N4254)? mem[186] : 
                 (N4256)? mem[188] : 
                 (N4258)? mem[190] : 
                 (N4260)? mem[192] : 
                 (N4262)? mem[194] : 
                 (N4264)? mem[196] : 
                 (N4266)? mem[198] : 
                 (N4268)? mem[200] : 
                 (N4270)? mem[202] : 
                 (N4272)? mem[204] : 
                 (N4274)? mem[206] : 
                 (N4276)? mem[208] : 
                 (N4278)? mem[210] : 
                 (N4280)? mem[212] : 
                 (N4282)? mem[214] : 
                 (N4284)? mem[216] : 
                 (N4286)? mem[218] : 
                 (N4288)? mem[220] : 
                 (N4290)? mem[222] : 
                 (N4292)? mem[224] : 
                 (N4294)? mem[226] : 
                 (N4296)? mem[228] : 
                 (N4298)? mem[230] : 
                 (N4300)? mem[232] : 
                 (N4302)? mem[234] : 
                 (N4304)? mem[236] : 
                 (N4306)? mem[238] : 
                 (N4308)? mem[240] : 
                 (N4310)? mem[242] : 
                 (N4312)? mem[244] : 
                 (N4314)? mem[246] : 
                 (N4316)? mem[248] : 
                 (N4318)? mem[250] : 
                 (N4320)? mem[252] : 
                 (N4322)? mem[254] : 
                 (N4324)? mem[256] : 
                 (N4326)? mem[258] : 
                 (N4328)? mem[260] : 
                 (N4330)? mem[262] : 
                 (N4332)? mem[264] : 
                 (N4334)? mem[266] : 
                 (N4336)? mem[268] : 
                 (N4338)? mem[270] : 
                 (N4340)? mem[272] : 
                 (N4342)? mem[274] : 
                 (N4344)? mem[276] : 
                 (N4346)? mem[278] : 
                 (N4348)? mem[280] : 
                 (N4350)? mem[282] : 
                 (N4352)? mem[284] : 
                 (N4354)? mem[286] : 
                 (N4356)? mem[288] : 
                 (N4358)? mem[290] : 
                 (N4360)? mem[292] : 
                 (N4362)? mem[294] : 
                 (N4364)? mem[296] : 
                 (N4366)? mem[298] : 
                 (N4368)? mem[300] : 
                 (N4370)? mem[302] : 
                 (N4372)? mem[304] : 
                 (N4374)? mem[306] : 
                 (N4376)? mem[308] : 
                 (N4378)? mem[310] : 
                 (N4380)? mem[312] : 
                 (N4382)? mem[314] : 
                 (N4384)? mem[316] : 
                 (N4386)? mem[318] : 
                 (N4388)? mem[320] : 
                 (N4390)? mem[322] : 
                 (N4392)? mem[324] : 
                 (N4394)? mem[326] : 
                 (N4396)? mem[328] : 
                 (N4398)? mem[330] : 
                 (N4400)? mem[332] : 
                 (N4402)? mem[334] : 
                 (N4404)? mem[336] : 
                 (N4406)? mem[338] : 
                 (N4408)? mem[340] : 
                 (N4410)? mem[342] : 
                 (N4412)? mem[344] : 
                 (N4414)? mem[346] : 
                 (N4416)? mem[348] : 
                 (N4418)? mem[350] : 
                 (N4420)? mem[352] : 
                 (N4422)? mem[354] : 
                 (N4424)? mem[356] : 
                 (N4426)? mem[358] : 
                 (N4428)? mem[360] : 
                 (N4430)? mem[362] : 
                 (N4432)? mem[364] : 
                 (N4434)? mem[366] : 
                 (N4436)? mem[368] : 
                 (N4438)? mem[370] : 
                 (N4440)? mem[372] : 
                 (N4442)? mem[374] : 
                 (N4444)? mem[376] : 
                 (N4446)? mem[378] : 
                 (N4448)? mem[380] : 
                 (N4450)? mem[382] : 
                 (N4452)? mem[384] : 
                 (N4454)? mem[386] : 
                 (N4456)? mem[388] : 
                 (N4458)? mem[390] : 
                 (N4460)? mem[392] : 
                 (N4462)? mem[394] : 
                 (N4464)? mem[396] : 
                 (N4466)? mem[398] : 
                 (N4468)? mem[400] : 
                 (N4470)? mem[402] : 
                 (N4472)? mem[404] : 
                 (N4474)? mem[406] : 
                 (N4476)? mem[408] : 
                 (N4478)? mem[410] : 
                 (N4480)? mem[412] : 
                 (N4482)? mem[414] : 
                 (N4484)? mem[416] : 
                 (N4486)? mem[418] : 
                 (N4488)? mem[420] : 
                 (N4490)? mem[422] : 
                 (N4492)? mem[424] : 
                 (N4494)? mem[426] : 
                 (N4496)? mem[428] : 
                 (N4498)? mem[430] : 
                 (N4500)? mem[432] : 
                 (N4502)? mem[434] : 
                 (N4504)? mem[436] : 
                 (N4506)? mem[438] : 
                 (N4508)? mem[440] : 
                 (N4510)? mem[442] : 
                 (N4512)? mem[444] : 
                 (N4514)? mem[446] : 
                 (N4516)? mem[448] : 
                 (N4518)? mem[450] : 
                 (N4520)? mem[452] : 
                 (N4522)? mem[454] : 
                 (N4524)? mem[456] : 
                 (N4526)? mem[458] : 
                 (N4528)? mem[460] : 
                 (N4530)? mem[462] : 
                 (N4532)? mem[464] : 
                 (N4534)? mem[466] : 
                 (N4536)? mem[468] : 
                 (N4538)? mem[470] : 
                 (N4540)? mem[472] : 
                 (N4542)? mem[474] : 
                 (N4544)? mem[476] : 
                 (N4546)? mem[478] : 
                 (N4548)? mem[480] : 
                 (N4549)? mem[482] : 
                 (N4550)? mem[484] : 
                 (N4551)? mem[486] : 
                 (N4552)? mem[488] : 
                 (N4553)? mem[490] : 
                 (N4554)? mem[492] : 
                 (N4555)? mem[494] : 
                 (N4556)? mem[496] : 
                 (N4557)? mem[498] : 
                 (N4558)? mem[500] : 
                 (N4559)? mem[502] : 
                 (N4560)? mem[504] : 
                 (N4561)? mem[506] : 
                 (N4562)? mem[508] : 
                 (N4563)? mem[510] : 
                 (N4069)? mem[512] : 
                 (N4071)? mem[514] : 
                 (N4073)? mem[516] : 
                 (N4075)? mem[518] : 
                 (N4077)? mem[520] : 
                 (N4079)? mem[522] : 
                 (N4081)? mem[524] : 
                 (N4083)? mem[526] : 
                 (N4085)? mem[528] : 
                 (N4087)? mem[530] : 
                 (N4089)? mem[532] : 
                 (N4091)? mem[534] : 
                 (N4093)? mem[536] : 
                 (N4095)? mem[538] : 
                 (N4097)? mem[540] : 
                 (N4099)? mem[542] : 
                 (N4101)? mem[544] : 
                 (N4103)? mem[546] : 
                 (N4105)? mem[548] : 
                 (N4107)? mem[550] : 
                 (N4109)? mem[552] : 
                 (N4111)? mem[554] : 
                 (N4113)? mem[556] : 
                 (N4115)? mem[558] : 
                 (N4117)? mem[560] : 
                 (N4119)? mem[562] : 
                 (N4121)? mem[564] : 
                 (N4123)? mem[566] : 
                 (N4125)? mem[568] : 
                 (N4127)? mem[570] : 
                 (N4129)? mem[572] : 
                 (N4131)? mem[574] : 
                 (N4133)? mem[576] : 
                 (N4135)? mem[578] : 
                 (N4137)? mem[580] : 
                 (N4139)? mem[582] : 
                 (N4141)? mem[584] : 
                 (N4143)? mem[586] : 
                 (N4145)? mem[588] : 
                 (N4147)? mem[590] : 
                 (N4149)? mem[592] : 
                 (N4151)? mem[594] : 
                 (N4153)? mem[596] : 
                 (N4155)? mem[598] : 
                 (N4157)? mem[600] : 
                 (N4159)? mem[602] : 
                 (N4161)? mem[604] : 
                 (N4163)? mem[606] : 
                 (N4165)? mem[608] : 
                 (N4167)? mem[610] : 
                 (N4169)? mem[612] : 
                 (N4171)? mem[614] : 
                 (N4173)? mem[616] : 
                 (N4175)? mem[618] : 
                 (N4177)? mem[620] : 
                 (N4179)? mem[622] : 
                 (N4181)? mem[624] : 
                 (N4183)? mem[626] : 
                 (N4185)? mem[628] : 
                 (N4187)? mem[630] : 
                 (N4189)? mem[632] : 
                 (N4191)? mem[634] : 
                 (N4193)? mem[636] : 
                 (N4195)? mem[638] : 
                 (N4197)? mem[640] : 
                 (N4199)? mem[642] : 
                 (N4201)? mem[644] : 
                 (N4203)? mem[646] : 
                 (N4205)? mem[648] : 
                 (N4207)? mem[650] : 
                 (N4209)? mem[652] : 
                 (N4211)? mem[654] : 
                 (N4213)? mem[656] : 
                 (N4215)? mem[658] : 
                 (N4217)? mem[660] : 
                 (N4219)? mem[662] : 
                 (N4221)? mem[664] : 
                 (N4223)? mem[666] : 
                 (N4225)? mem[668] : 
                 (N4227)? mem[670] : 
                 (N4229)? mem[672] : 
                 (N4231)? mem[674] : 
                 (N4233)? mem[676] : 
                 (N4235)? mem[678] : 
                 (N4237)? mem[680] : 
                 (N4239)? mem[682] : 
                 (N4241)? mem[684] : 
                 (N4243)? mem[686] : 
                 (N4245)? mem[688] : 
                 (N4247)? mem[690] : 
                 (N4249)? mem[692] : 
                 (N4251)? mem[694] : 
                 (N4253)? mem[696] : 
                 (N4255)? mem[698] : 
                 (N4257)? mem[700] : 
                 (N4259)? mem[702] : 
                 (N4261)? mem[704] : 
                 (N4263)? mem[706] : 
                 (N4265)? mem[708] : 
                 (N4267)? mem[710] : 
                 (N4269)? mem[712] : 
                 (N4271)? mem[714] : 
                 (N4273)? mem[716] : 
                 (N4275)? mem[718] : 
                 (N4277)? mem[720] : 
                 (N4279)? mem[722] : 
                 (N4281)? mem[724] : 
                 (N4283)? mem[726] : 
                 (N4285)? mem[728] : 
                 (N4287)? mem[730] : 
                 (N4289)? mem[732] : 
                 (N4291)? mem[734] : 
                 (N4293)? mem[736] : 
                 (N4295)? mem[738] : 
                 (N4297)? mem[740] : 
                 (N4299)? mem[742] : 
                 (N4301)? mem[744] : 
                 (N4303)? mem[746] : 
                 (N4305)? mem[748] : 
                 (N4307)? mem[750] : 
                 (N4309)? mem[752] : 
                 (N4311)? mem[754] : 
                 (N4313)? mem[756] : 
                 (N4315)? mem[758] : 
                 (N4317)? mem[760] : 
                 (N4319)? mem[762] : 
                 (N4321)? mem[764] : 
                 (N4323)? mem[766] : 
                 (N4325)? mem[768] : 
                 (N4327)? mem[770] : 
                 (N4329)? mem[772] : 
                 (N4331)? mem[774] : 
                 (N4333)? mem[776] : 
                 (N4335)? mem[778] : 
                 (N4337)? mem[780] : 
                 (N4339)? mem[782] : 
                 (N4341)? mem[784] : 
                 (N4343)? mem[786] : 
                 (N4345)? mem[788] : 
                 (N4347)? mem[790] : 
                 (N4349)? mem[792] : 
                 (N4351)? mem[794] : 
                 (N4353)? mem[796] : 
                 (N4355)? mem[798] : 
                 (N4357)? mem[800] : 
                 (N4359)? mem[802] : 
                 (N4361)? mem[804] : 
                 (N4363)? mem[806] : 
                 (N4365)? mem[808] : 
                 (N4367)? mem[810] : 
                 (N4369)? mem[812] : 
                 (N4371)? mem[814] : 
                 (N4373)? mem[816] : 
                 (N4375)? mem[818] : 
                 (N4377)? mem[820] : 
                 (N4379)? mem[822] : 
                 (N4381)? mem[824] : 
                 (N4383)? mem[826] : 
                 (N4385)? mem[828] : 
                 (N4387)? mem[830] : 
                 (N4389)? mem[832] : 
                 (N4391)? mem[834] : 
                 (N4393)? mem[836] : 
                 (N4395)? mem[838] : 
                 (N4397)? mem[840] : 
                 (N4399)? mem[842] : 
                 (N4401)? mem[844] : 
                 (N4403)? mem[846] : 
                 (N4405)? mem[848] : 
                 (N4407)? mem[850] : 
                 (N4409)? mem[852] : 
                 (N4411)? mem[854] : 
                 (N4413)? mem[856] : 
                 (N4415)? mem[858] : 
                 (N4417)? mem[860] : 
                 (N4419)? mem[862] : 
                 (N4421)? mem[864] : 
                 (N4423)? mem[866] : 
                 (N4425)? mem[868] : 
                 (N4427)? mem[870] : 
                 (N4429)? mem[872] : 
                 (N4431)? mem[874] : 
                 (N4433)? mem[876] : 
                 (N4435)? mem[878] : 
                 (N4437)? mem[880] : 
                 (N4439)? mem[882] : 
                 (N4441)? mem[884] : 
                 (N4443)? mem[886] : 
                 (N4445)? mem[888] : 
                 (N4447)? mem[890] : 
                 (N4449)? mem[892] : 
                 (N4451)? mem[894] : 
                 (N4453)? mem[896] : 
                 (N4455)? mem[898] : 
                 (N4457)? mem[900] : 
                 (N4459)? mem[902] : 
                 (N4461)? mem[904] : 
                 (N4463)? mem[906] : 
                 (N4465)? mem[908] : 
                 (N4467)? mem[910] : 
                 (N4469)? mem[912] : 
                 (N4471)? mem[914] : 
                 (N4473)? mem[916] : 
                 (N4475)? mem[918] : 
                 (N4477)? mem[920] : 
                 (N4479)? mem[922] : 
                 (N4481)? mem[924] : 
                 (N4483)? mem[926] : 
                 (N4485)? mem[928] : 
                 (N4487)? mem[930] : 
                 (N4489)? mem[932] : 
                 (N4491)? mem[934] : 
                 (N4493)? mem[936] : 
                 (N4495)? mem[938] : 
                 (N4497)? mem[940] : 
                 (N4499)? mem[942] : 
                 (N4501)? mem[944] : 
                 (N4503)? mem[946] : 
                 (N4505)? mem[948] : 
                 (N4507)? mem[950] : 
                 (N4509)? mem[952] : 
                 (N4511)? mem[954] : 
                 (N4513)? mem[956] : 
                 (N4515)? mem[958] : 
                 (N4517)? mem[960] : 
                 (N4519)? mem[962] : 
                 (N4521)? mem[964] : 
                 (N4523)? mem[966] : 
                 (N4525)? mem[968] : 
                 (N4527)? mem[970] : 
                 (N4529)? mem[972] : 
                 (N4531)? mem[974] : 
                 (N4533)? mem[976] : 
                 (N4535)? mem[978] : 
                 (N4537)? mem[980] : 
                 (N4539)? mem[982] : 
                 (N4541)? mem[984] : 
                 (N4543)? mem[986] : 
                 (N4545)? mem[988] : 
                 (N4547)? mem[990] : 
                 (N3628)? mem[992] : 
                 (N3630)? mem[994] : 
                 (N3632)? mem[996] : 
                 (N3634)? mem[998] : 
                 (N3636)? mem[1000] : 
                 (N3638)? mem[1002] : 
                 (N3640)? mem[1004] : 
                 (N3642)? mem[1006] : 
                 (N12097)? mem[1008] : 
                 (N12099)? mem[1010] : 
                 (N12101)? mem[1012] : 
                 (N12103)? mem[1014] : 
                 (N12105)? mem[1016] : 
                 (N12107)? mem[1018] : 
                 (N12109)? mem[1020] : 
                 (N12111)? mem[1022] : 1'b0;
  assign N5950 = (N5462)? mem[1] : 
                 (N5464)? mem[3] : 
                 (N5466)? mem[5] : 
                 (N5468)? mem[7] : 
                 (N5470)? mem[9] : 
                 (N5472)? mem[11] : 
                 (N5474)? mem[13] : 
                 (N5476)? mem[15] : 
                 (N5478)? mem[17] : 
                 (N5480)? mem[19] : 
                 (N5482)? mem[21] : 
                 (N5484)? mem[23] : 
                 (N5486)? mem[25] : 
                 (N5488)? mem[27] : 
                 (N5490)? mem[29] : 
                 (N5492)? mem[31] : 
                 (N5494)? mem[33] : 
                 (N5496)? mem[35] : 
                 (N5498)? mem[37] : 
                 (N5500)? mem[39] : 
                 (N5502)? mem[41] : 
                 (N5504)? mem[43] : 
                 (N5506)? mem[45] : 
                 (N5508)? mem[47] : 
                 (N5510)? mem[49] : 
                 (N5512)? mem[51] : 
                 (N5514)? mem[53] : 
                 (N5516)? mem[55] : 
                 (N5518)? mem[57] : 
                 (N5520)? mem[59] : 
                 (N5522)? mem[61] : 
                 (N5524)? mem[63] : 
                 (N5526)? mem[65] : 
                 (N5528)? mem[67] : 
                 (N5530)? mem[69] : 
                 (N5532)? mem[71] : 
                 (N5534)? mem[73] : 
                 (N5536)? mem[75] : 
                 (N5538)? mem[77] : 
                 (N5540)? mem[79] : 
                 (N5542)? mem[81] : 
                 (N5544)? mem[83] : 
                 (N5546)? mem[85] : 
                 (N5548)? mem[87] : 
                 (N5550)? mem[89] : 
                 (N5552)? mem[91] : 
                 (N5554)? mem[93] : 
                 (N5556)? mem[95] : 
                 (N5558)? mem[97] : 
                 (N5560)? mem[99] : 
                 (N5562)? mem[101] : 
                 (N5564)? mem[103] : 
                 (N5566)? mem[105] : 
                 (N5568)? mem[107] : 
                 (N5570)? mem[109] : 
                 (N5572)? mem[111] : 
                 (N5574)? mem[113] : 
                 (N5576)? mem[115] : 
                 (N5578)? mem[117] : 
                 (N5580)? mem[119] : 
                 (N5582)? mem[121] : 
                 (N5584)? mem[123] : 
                 (N5586)? mem[125] : 
                 (N5588)? mem[127] : 
                 (N5590)? mem[129] : 
                 (N5592)? mem[131] : 
                 (N5594)? mem[133] : 
                 (N5596)? mem[135] : 
                 (N5598)? mem[137] : 
                 (N5600)? mem[139] : 
                 (N5602)? mem[141] : 
                 (N5604)? mem[143] : 
                 (N5606)? mem[145] : 
                 (N5608)? mem[147] : 
                 (N5610)? mem[149] : 
                 (N5612)? mem[151] : 
                 (N5614)? mem[153] : 
                 (N5616)? mem[155] : 
                 (N5618)? mem[157] : 
                 (N5620)? mem[159] : 
                 (N5622)? mem[161] : 
                 (N5624)? mem[163] : 
                 (N5626)? mem[165] : 
                 (N5628)? mem[167] : 
                 (N5630)? mem[169] : 
                 (N5632)? mem[171] : 
                 (N5634)? mem[173] : 
                 (N5636)? mem[175] : 
                 (N5638)? mem[177] : 
                 (N5640)? mem[179] : 
                 (N5642)? mem[181] : 
                 (N5644)? mem[183] : 
                 (N5646)? mem[185] : 
                 (N5648)? mem[187] : 
                 (N5650)? mem[189] : 
                 (N5652)? mem[191] : 
                 (N5654)? mem[193] : 
                 (N5656)? mem[195] : 
                 (N5658)? mem[197] : 
                 (N5660)? mem[199] : 
                 (N5662)? mem[201] : 
                 (N5664)? mem[203] : 
                 (N5666)? mem[205] : 
                 (N5668)? mem[207] : 
                 (N5670)? mem[209] : 
                 (N5672)? mem[211] : 
                 (N5674)? mem[213] : 
                 (N5676)? mem[215] : 
                 (N5678)? mem[217] : 
                 (N5680)? mem[219] : 
                 (N5682)? mem[221] : 
                 (N5684)? mem[223] : 
                 (N5686)? mem[225] : 
                 (N5688)? mem[227] : 
                 (N5690)? mem[229] : 
                 (N5692)? mem[231] : 
                 (N5694)? mem[233] : 
                 (N5696)? mem[235] : 
                 (N5698)? mem[237] : 
                 (N5700)? mem[239] : 
                 (N5702)? mem[241] : 
                 (N5704)? mem[243] : 
                 (N5706)? mem[245] : 
                 (N5708)? mem[247] : 
                 (N5710)? mem[249] : 
                 (N5712)? mem[251] : 
                 (N5714)? mem[253] : 
                 (N5716)? mem[255] : 
                 (N5718)? mem[257] : 
                 (N5720)? mem[259] : 
                 (N5722)? mem[261] : 
                 (N5724)? mem[263] : 
                 (N5726)? mem[265] : 
                 (N5728)? mem[267] : 
                 (N5730)? mem[269] : 
                 (N5732)? mem[271] : 
                 (N5734)? mem[273] : 
                 (N5736)? mem[275] : 
                 (N5738)? mem[277] : 
                 (N5740)? mem[279] : 
                 (N5742)? mem[281] : 
                 (N5744)? mem[283] : 
                 (N5746)? mem[285] : 
                 (N5748)? mem[287] : 
                 (N5750)? mem[289] : 
                 (N5752)? mem[291] : 
                 (N5754)? mem[293] : 
                 (N5756)? mem[295] : 
                 (N5758)? mem[297] : 
                 (N5760)? mem[299] : 
                 (N5762)? mem[301] : 
                 (N5764)? mem[303] : 
                 (N5766)? mem[305] : 
                 (N5768)? mem[307] : 
                 (N5770)? mem[309] : 
                 (N5772)? mem[311] : 
                 (N5774)? mem[313] : 
                 (N5776)? mem[315] : 
                 (N5778)? mem[317] : 
                 (N5780)? mem[319] : 
                 (N5782)? mem[321] : 
                 (N5784)? mem[323] : 
                 (N5786)? mem[325] : 
                 (N5788)? mem[327] : 
                 (N5790)? mem[329] : 
                 (N5792)? mem[331] : 
                 (N5794)? mem[333] : 
                 (N5796)? mem[335] : 
                 (N5798)? mem[337] : 
                 (N5800)? mem[339] : 
                 (N5802)? mem[341] : 
                 (N5804)? mem[343] : 
                 (N5806)? mem[345] : 
                 (N5808)? mem[347] : 
                 (N5810)? mem[349] : 
                 (N5812)? mem[351] : 
                 (N5814)? mem[353] : 
                 (N5816)? mem[355] : 
                 (N5818)? mem[357] : 
                 (N5820)? mem[359] : 
                 (N5822)? mem[361] : 
                 (N5824)? mem[363] : 
                 (N5826)? mem[365] : 
                 (N5828)? mem[367] : 
                 (N5830)? mem[369] : 
                 (N5832)? mem[371] : 
                 (N5834)? mem[373] : 
                 (N5836)? mem[375] : 
                 (N5838)? mem[377] : 
                 (N5840)? mem[379] : 
                 (N5842)? mem[381] : 
                 (N5844)? mem[383] : 
                 (N5846)? mem[385] : 
                 (N5848)? mem[387] : 
                 (N5850)? mem[389] : 
                 (N5852)? mem[391] : 
                 (N5854)? mem[393] : 
                 (N5856)? mem[395] : 
                 (N5858)? mem[397] : 
                 (N5860)? mem[399] : 
                 (N5862)? mem[401] : 
                 (N5864)? mem[403] : 
                 (N5866)? mem[405] : 
                 (N5868)? mem[407] : 
                 (N5870)? mem[409] : 
                 (N5872)? mem[411] : 
                 (N5874)? mem[413] : 
                 (N5876)? mem[415] : 
                 (N5878)? mem[417] : 
                 (N5880)? mem[419] : 
                 (N5882)? mem[421] : 
                 (N5884)? mem[423] : 
                 (N5886)? mem[425] : 
                 (N5888)? mem[427] : 
                 (N5890)? mem[429] : 
                 (N5892)? mem[431] : 
                 (N5894)? mem[433] : 
                 (N5896)? mem[435] : 
                 (N5898)? mem[437] : 
                 (N5900)? mem[439] : 
                 (N5902)? mem[441] : 
                 (N5904)? mem[443] : 
                 (N5906)? mem[445] : 
                 (N5908)? mem[447] : 
                 (N5910)? mem[449] : 
                 (N5912)? mem[451] : 
                 (N5914)? mem[453] : 
                 (N5916)? mem[455] : 
                 (N5918)? mem[457] : 
                 (N5920)? mem[459] : 
                 (N5922)? mem[461] : 
                 (N5924)? mem[463] : 
                 (N5926)? mem[465] : 
                 (N5927)? mem[467] : 
                 (N5928)? mem[469] : 
                 (N5929)? mem[471] : 
                 (N5930)? mem[473] : 
                 (N5931)? mem[475] : 
                 (N5932)? mem[477] : 
                 (N5933)? mem[479] : 
                 (N5934)? mem[481] : 
                 (N5935)? mem[483] : 
                 (N5936)? mem[485] : 
                 (N5937)? mem[487] : 
                 (N5938)? mem[489] : 
                 (N5939)? mem[491] : 
                 (N5940)? mem[493] : 
                 (N5941)? mem[495] : 
                 (N5942)? mem[497] : 
                 (N5943)? mem[499] : 
                 (N5944)? mem[501] : 
                 (N5945)? mem[503] : 
                 (N5946)? mem[505] : 
                 (N5947)? mem[507] : 
                 (N5948)? mem[509] : 
                 (N5949)? mem[511] : 
                 (N5463)? mem[513] : 
                 (N5465)? mem[515] : 
                 (N5467)? mem[517] : 
                 (N5469)? mem[519] : 
                 (N5471)? mem[521] : 
                 (N5473)? mem[523] : 
                 (N5475)? mem[525] : 
                 (N5477)? mem[527] : 
                 (N5479)? mem[529] : 
                 (N5481)? mem[531] : 
                 (N5483)? mem[533] : 
                 (N5485)? mem[535] : 
                 (N5487)? mem[537] : 
                 (N5489)? mem[539] : 
                 (N5491)? mem[541] : 
                 (N5493)? mem[543] : 
                 (N5495)? mem[545] : 
                 (N5497)? mem[547] : 
                 (N5499)? mem[549] : 
                 (N5501)? mem[551] : 
                 (N5503)? mem[553] : 
                 (N5505)? mem[555] : 
                 (N5507)? mem[557] : 
                 (N5509)? mem[559] : 
                 (N5511)? mem[561] : 
                 (N5513)? mem[563] : 
                 (N5515)? mem[565] : 
                 (N5517)? mem[567] : 
                 (N5519)? mem[569] : 
                 (N5521)? mem[571] : 
                 (N5523)? mem[573] : 
                 (N5525)? mem[575] : 
                 (N5527)? mem[577] : 
                 (N5529)? mem[579] : 
                 (N5531)? mem[581] : 
                 (N5533)? mem[583] : 
                 (N5535)? mem[585] : 
                 (N5537)? mem[587] : 
                 (N5539)? mem[589] : 
                 (N5541)? mem[591] : 
                 (N5543)? mem[593] : 
                 (N5545)? mem[595] : 
                 (N5547)? mem[597] : 
                 (N5549)? mem[599] : 
                 (N5551)? mem[601] : 
                 (N5553)? mem[603] : 
                 (N5555)? mem[605] : 
                 (N5557)? mem[607] : 
                 (N5559)? mem[609] : 
                 (N5561)? mem[611] : 
                 (N5563)? mem[613] : 
                 (N5565)? mem[615] : 
                 (N5567)? mem[617] : 
                 (N5569)? mem[619] : 
                 (N5571)? mem[621] : 
                 (N5573)? mem[623] : 
                 (N5575)? mem[625] : 
                 (N5577)? mem[627] : 
                 (N5579)? mem[629] : 
                 (N5581)? mem[631] : 
                 (N5583)? mem[633] : 
                 (N5585)? mem[635] : 
                 (N5587)? mem[637] : 
                 (N5589)? mem[639] : 
                 (N5591)? mem[641] : 
                 (N5593)? mem[643] : 
                 (N5595)? mem[645] : 
                 (N5597)? mem[647] : 
                 (N5599)? mem[649] : 
                 (N5601)? mem[651] : 
                 (N5603)? mem[653] : 
                 (N5605)? mem[655] : 
                 (N5607)? mem[657] : 
                 (N5609)? mem[659] : 
                 (N5611)? mem[661] : 
                 (N5613)? mem[663] : 
                 (N5615)? mem[665] : 
                 (N5617)? mem[667] : 
                 (N5619)? mem[669] : 
                 (N5621)? mem[671] : 
                 (N5623)? mem[673] : 
                 (N5625)? mem[675] : 
                 (N5627)? mem[677] : 
                 (N5629)? mem[679] : 
                 (N5631)? mem[681] : 
                 (N5633)? mem[683] : 
                 (N5635)? mem[685] : 
                 (N5637)? mem[687] : 
                 (N5639)? mem[689] : 
                 (N5641)? mem[691] : 
                 (N5643)? mem[693] : 
                 (N5645)? mem[695] : 
                 (N5647)? mem[697] : 
                 (N5649)? mem[699] : 
                 (N5651)? mem[701] : 
                 (N5653)? mem[703] : 
                 (N5655)? mem[705] : 
                 (N5657)? mem[707] : 
                 (N5659)? mem[709] : 
                 (N5661)? mem[711] : 
                 (N5663)? mem[713] : 
                 (N5665)? mem[715] : 
                 (N5667)? mem[717] : 
                 (N5669)? mem[719] : 
                 (N5671)? mem[721] : 
                 (N5673)? mem[723] : 
                 (N5675)? mem[725] : 
                 (N5677)? mem[727] : 
                 (N5679)? mem[729] : 
                 (N5681)? mem[731] : 
                 (N5683)? mem[733] : 
                 (N5685)? mem[735] : 
                 (N5687)? mem[737] : 
                 (N5689)? mem[739] : 
                 (N5691)? mem[741] : 
                 (N5693)? mem[743] : 
                 (N5695)? mem[745] : 
                 (N5697)? mem[747] : 
                 (N5699)? mem[749] : 
                 (N5701)? mem[751] : 
                 (N5703)? mem[753] : 
                 (N5705)? mem[755] : 
                 (N5707)? mem[757] : 
                 (N5709)? mem[759] : 
                 (N5711)? mem[761] : 
                 (N5713)? mem[763] : 
                 (N5715)? mem[765] : 
                 (N5717)? mem[767] : 
                 (N5719)? mem[769] : 
                 (N5721)? mem[771] : 
                 (N5723)? mem[773] : 
                 (N5725)? mem[775] : 
                 (N5727)? mem[777] : 
                 (N5729)? mem[779] : 
                 (N5731)? mem[781] : 
                 (N5733)? mem[783] : 
                 (N5735)? mem[785] : 
                 (N5737)? mem[787] : 
                 (N5739)? mem[789] : 
                 (N5741)? mem[791] : 
                 (N5743)? mem[793] : 
                 (N5745)? mem[795] : 
                 (N5747)? mem[797] : 
                 (N5749)? mem[799] : 
                 (N5751)? mem[801] : 
                 (N5753)? mem[803] : 
                 (N5755)? mem[805] : 
                 (N5757)? mem[807] : 
                 (N5759)? mem[809] : 
                 (N5761)? mem[811] : 
                 (N5763)? mem[813] : 
                 (N5765)? mem[815] : 
                 (N5767)? mem[817] : 
                 (N5769)? mem[819] : 
                 (N5771)? mem[821] : 
                 (N5773)? mem[823] : 
                 (N5775)? mem[825] : 
                 (N5777)? mem[827] : 
                 (N5779)? mem[829] : 
                 (N5781)? mem[831] : 
                 (N5783)? mem[833] : 
                 (N5785)? mem[835] : 
                 (N5787)? mem[837] : 
                 (N5789)? mem[839] : 
                 (N5791)? mem[841] : 
                 (N5793)? mem[843] : 
                 (N5795)? mem[845] : 
                 (N5797)? mem[847] : 
                 (N5799)? mem[849] : 
                 (N5801)? mem[851] : 
                 (N5803)? mem[853] : 
                 (N5805)? mem[855] : 
                 (N5807)? mem[857] : 
                 (N5809)? mem[859] : 
                 (N5811)? mem[861] : 
                 (N5813)? mem[863] : 
                 (N5815)? mem[865] : 
                 (N5817)? mem[867] : 
                 (N5819)? mem[869] : 
                 (N5821)? mem[871] : 
                 (N5823)? mem[873] : 
                 (N5825)? mem[875] : 
                 (N5827)? mem[877] : 
                 (N5829)? mem[879] : 
                 (N5831)? mem[881] : 
                 (N5833)? mem[883] : 
                 (N5835)? mem[885] : 
                 (N5837)? mem[887] : 
                 (N5839)? mem[889] : 
                 (N5841)? mem[891] : 
                 (N5843)? mem[893] : 
                 (N5845)? mem[895] : 
                 (N5847)? mem[897] : 
                 (N5849)? mem[899] : 
                 (N5851)? mem[901] : 
                 (N5853)? mem[903] : 
                 (N5855)? mem[905] : 
                 (N5857)? mem[907] : 
                 (N5859)? mem[909] : 
                 (N5861)? mem[911] : 
                 (N5863)? mem[913] : 
                 (N5865)? mem[915] : 
                 (N5867)? mem[917] : 
                 (N5869)? mem[919] : 
                 (N5871)? mem[921] : 
                 (N5873)? mem[923] : 
                 (N5875)? mem[925] : 
                 (N5877)? mem[927] : 
                 (N5879)? mem[929] : 
                 (N5881)? mem[931] : 
                 (N5883)? mem[933] : 
                 (N5885)? mem[935] : 
                 (N5887)? mem[937] : 
                 (N5889)? mem[939] : 
                 (N5891)? mem[941] : 
                 (N5893)? mem[943] : 
                 (N5895)? mem[945] : 
                 (N5897)? mem[947] : 
                 (N5899)? mem[949] : 
                 (N5901)? mem[951] : 
                 (N5903)? mem[953] : 
                 (N5905)? mem[955] : 
                 (N5907)? mem[957] : 
                 (N5909)? mem[959] : 
                 (N5911)? mem[961] : 
                 (N5913)? mem[963] : 
                 (N5915)? mem[965] : 
                 (N5917)? mem[967] : 
                 (N5919)? mem[969] : 
                 (N5921)? mem[971] : 
                 (N5923)? mem[973] : 
                 (N5925)? mem[975] : 
                 (N4533)? mem[977] : 
                 (N4535)? mem[979] : 
                 (N4537)? mem[981] : 
                 (N4539)? mem[983] : 
                 (N4541)? mem[985] : 
                 (N4543)? mem[987] : 
                 (N4545)? mem[989] : 
                 (N4547)? mem[991] : 
                 (N12081)? mem[993] : 
                 (N12083)? mem[995] : 
                 (N12085)? mem[997] : 
                 (N12087)? mem[999] : 
                 (N12089)? mem[1001] : 
                 (N12091)? mem[1003] : 
                 (N12093)? mem[1005] : 
                 (N12095)? mem[1007] : 
                 (N12097)? mem[1009] : 
                 (N12099)? mem[1011] : 
                 (N12101)? mem[1013] : 
                 (N12103)? mem[1015] : 
                 (N12105)? mem[1017] : 
                 (N12107)? mem[1019] : 
                 (N12109)? mem[1021] : 
                 (N12111)? mem[1023] : 1'b0;
  assign N6759 = (N6287)? mem[0] : 
                 (N6289)? mem[2] : 
                 (N6291)? mem[4] : 
                 (N6293)? mem[6] : 
                 (N6295)? mem[8] : 
                 (N6297)? mem[10] : 
                 (N6299)? mem[12] : 
                 (N6301)? mem[14] : 
                 (N6303)? mem[16] : 
                 (N6305)? mem[18] : 
                 (N6307)? mem[20] : 
                 (N6309)? mem[22] : 
                 (N6311)? mem[24] : 
                 (N6313)? mem[26] : 
                 (N6315)? mem[28] : 
                 (N6317)? mem[30] : 
                 (N6319)? mem[32] : 
                 (N6321)? mem[34] : 
                 (N6323)? mem[36] : 
                 (N6325)? mem[38] : 
                 (N6327)? mem[40] : 
                 (N6329)? mem[42] : 
                 (N6331)? mem[44] : 
                 (N6333)? mem[46] : 
                 (N6335)? mem[48] : 
                 (N6337)? mem[50] : 
                 (N6339)? mem[52] : 
                 (N6341)? mem[54] : 
                 (N6343)? mem[56] : 
                 (N6345)? mem[58] : 
                 (N6347)? mem[60] : 
                 (N6349)? mem[62] : 
                 (N6351)? mem[64] : 
                 (N6353)? mem[66] : 
                 (N6355)? mem[68] : 
                 (N6357)? mem[70] : 
                 (N6359)? mem[72] : 
                 (N6361)? mem[74] : 
                 (N6363)? mem[76] : 
                 (N6365)? mem[78] : 
                 (N6367)? mem[80] : 
                 (N6369)? mem[82] : 
                 (N6371)? mem[84] : 
                 (N6373)? mem[86] : 
                 (N6375)? mem[88] : 
                 (N6377)? mem[90] : 
                 (N6379)? mem[92] : 
                 (N6381)? mem[94] : 
                 (N6383)? mem[96] : 
                 (N6385)? mem[98] : 
                 (N6387)? mem[100] : 
                 (N6389)? mem[102] : 
                 (N6391)? mem[104] : 
                 (N6393)? mem[106] : 
                 (N6395)? mem[108] : 
                 (N6397)? mem[110] : 
                 (N6399)? mem[112] : 
                 (N6401)? mem[114] : 
                 (N6403)? mem[116] : 
                 (N6405)? mem[118] : 
                 (N6407)? mem[120] : 
                 (N6409)? mem[122] : 
                 (N6411)? mem[124] : 
                 (N6413)? mem[126] : 
                 (N6415)? mem[128] : 
                 (N6417)? mem[130] : 
                 (N6419)? mem[132] : 
                 (N6421)? mem[134] : 
                 (N6423)? mem[136] : 
                 (N6425)? mem[138] : 
                 (N6427)? mem[140] : 
                 (N6429)? mem[142] : 
                 (N6431)? mem[144] : 
                 (N6433)? mem[146] : 
                 (N6435)? mem[148] : 
                 (N6437)? mem[150] : 
                 (N6439)? mem[152] : 
                 (N6441)? mem[154] : 
                 (N6443)? mem[156] : 
                 (N6445)? mem[158] : 
                 (N6447)? mem[160] : 
                 (N6449)? mem[162] : 
                 (N6451)? mem[164] : 
                 (N6453)? mem[166] : 
                 (N6455)? mem[168] : 
                 (N6457)? mem[170] : 
                 (N6459)? mem[172] : 
                 (N6461)? mem[174] : 
                 (N6463)? mem[176] : 
                 (N6465)? mem[178] : 
                 (N6467)? mem[180] : 
                 (N6469)? mem[182] : 
                 (N6471)? mem[184] : 
                 (N6473)? mem[186] : 
                 (N6475)? mem[188] : 
                 (N6477)? mem[190] : 
                 (N6479)? mem[192] : 
                 (N6481)? mem[194] : 
                 (N6483)? mem[196] : 
                 (N6485)? mem[198] : 
                 (N6487)? mem[200] : 
                 (N6489)? mem[202] : 
                 (N6491)? mem[204] : 
                 (N6493)? mem[206] : 
                 (N6495)? mem[208] : 
                 (N6497)? mem[210] : 
                 (N6499)? mem[212] : 
                 (N6501)? mem[214] : 
                 (N6503)? mem[216] : 
                 (N6505)? mem[218] : 
                 (N6507)? mem[220] : 
                 (N6509)? mem[222] : 
                 (N6511)? mem[224] : 
                 (N6513)? mem[226] : 
                 (N6515)? mem[228] : 
                 (N6517)? mem[230] : 
                 (N6519)? mem[232] : 
                 (N6521)? mem[234] : 
                 (N6523)? mem[236] : 
                 (N6525)? mem[238] : 
                 (N6527)? mem[240] : 
                 (N6529)? mem[242] : 
                 (N6531)? mem[244] : 
                 (N6533)? mem[246] : 
                 (N6535)? mem[248] : 
                 (N6537)? mem[250] : 
                 (N6539)? mem[252] : 
                 (N6541)? mem[254] : 
                 (N6543)? mem[256] : 
                 (N6545)? mem[258] : 
                 (N6547)? mem[260] : 
                 (N6549)? mem[262] : 
                 (N6551)? mem[264] : 
                 (N6553)? mem[266] : 
                 (N6555)? mem[268] : 
                 (N6557)? mem[270] : 
                 (N6559)? mem[272] : 
                 (N6561)? mem[274] : 
                 (N6563)? mem[276] : 
                 (N6565)? mem[278] : 
                 (N6567)? mem[280] : 
                 (N6569)? mem[282] : 
                 (N6571)? mem[284] : 
                 (N6573)? mem[286] : 
                 (N6575)? mem[288] : 
                 (N6577)? mem[290] : 
                 (N6579)? mem[292] : 
                 (N6581)? mem[294] : 
                 (N6583)? mem[296] : 
                 (N6585)? mem[298] : 
                 (N6587)? mem[300] : 
                 (N6589)? mem[302] : 
                 (N6591)? mem[304] : 
                 (N6593)? mem[306] : 
                 (N6595)? mem[308] : 
                 (N6597)? mem[310] : 
                 (N6599)? mem[312] : 
                 (N6601)? mem[314] : 
                 (N6603)? mem[316] : 
                 (N6605)? mem[318] : 
                 (N6607)? mem[320] : 
                 (N6609)? mem[322] : 
                 (N6611)? mem[324] : 
                 (N6613)? mem[326] : 
                 (N6615)? mem[328] : 
                 (N6617)? mem[330] : 
                 (N6619)? mem[332] : 
                 (N6621)? mem[334] : 
                 (N6623)? mem[336] : 
                 (N6625)? mem[338] : 
                 (N6627)? mem[340] : 
                 (N6629)? mem[342] : 
                 (N6631)? mem[344] : 
                 (N6633)? mem[346] : 
                 (N6635)? mem[348] : 
                 (N6637)? mem[350] : 
                 (N6639)? mem[352] : 
                 (N6641)? mem[354] : 
                 (N6643)? mem[356] : 
                 (N6645)? mem[358] : 
                 (N6647)? mem[360] : 
                 (N6649)? mem[362] : 
                 (N6651)? mem[364] : 
                 (N6653)? mem[366] : 
                 (N6655)? mem[368] : 
                 (N6657)? mem[370] : 
                 (N6659)? mem[372] : 
                 (N6661)? mem[374] : 
                 (N6663)? mem[376] : 
                 (N6665)? mem[378] : 
                 (N6667)? mem[380] : 
                 (N6669)? mem[382] : 
                 (N6671)? mem[384] : 
                 (N6673)? mem[386] : 
                 (N6675)? mem[388] : 
                 (N6677)? mem[390] : 
                 (N6679)? mem[392] : 
                 (N6681)? mem[394] : 
                 (N6683)? mem[396] : 
                 (N6685)? mem[398] : 
                 (N6687)? mem[400] : 
                 (N6689)? mem[402] : 
                 (N6691)? mem[404] : 
                 (N6693)? mem[406] : 
                 (N6695)? mem[408] : 
                 (N6697)? mem[410] : 
                 (N6699)? mem[412] : 
                 (N6701)? mem[414] : 
                 (N6703)? mem[416] : 
                 (N6704)? mem[418] : 
                 (N6705)? mem[420] : 
                 (N6706)? mem[422] : 
                 (N6707)? mem[424] : 
                 (N6708)? mem[426] : 
                 (N6709)? mem[428] : 
                 (N6710)? mem[430] : 
                 (N6711)? mem[432] : 
                 (N6712)? mem[434] : 
                 (N6713)? mem[436] : 
                 (N6714)? mem[438] : 
                 (N6715)? mem[440] : 
                 (N6716)? mem[442] : 
                 (N6717)? mem[444] : 
                 (N6718)? mem[446] : 
                 (N6719)? mem[448] : 
                 (N6721)? mem[450] : 
                 (N6723)? mem[452] : 
                 (N6725)? mem[454] : 
                 (N6727)? mem[456] : 
                 (N6729)? mem[458] : 
                 (N6731)? mem[460] : 
                 (N6733)? mem[462] : 
                 (N6735)? mem[464] : 
                 (N6736)? mem[466] : 
                 (N6737)? mem[468] : 
                 (N6738)? mem[470] : 
                 (N6739)? mem[472] : 
                 (N6740)? mem[474] : 
                 (N6741)? mem[476] : 
                 (N6742)? mem[478] : 
                 (N6743)? mem[480] : 
                 (N6744)? mem[482] : 
                 (N6745)? mem[484] : 
                 (N6746)? mem[486] : 
                 (N6747)? mem[488] : 
                 (N6748)? mem[490] : 
                 (N6749)? mem[492] : 
                 (N6750)? mem[494] : 
                 (N6751)? mem[496] : 
                 (N6752)? mem[498] : 
                 (N6753)? mem[500] : 
                 (N6754)? mem[502] : 
                 (N6755)? mem[504] : 
                 (N6756)? mem[506] : 
                 (N6757)? mem[508] : 
                 (N6758)? mem[510] : 
                 (N6288)? mem[512] : 
                 (N6290)? mem[514] : 
                 (N6292)? mem[516] : 
                 (N6294)? mem[518] : 
                 (N6296)? mem[520] : 
                 (N6298)? mem[522] : 
                 (N6300)? mem[524] : 
                 (N6302)? mem[526] : 
                 (N6304)? mem[528] : 
                 (N6306)? mem[530] : 
                 (N6308)? mem[532] : 
                 (N6310)? mem[534] : 
                 (N6312)? mem[536] : 
                 (N6314)? mem[538] : 
                 (N6316)? mem[540] : 
                 (N6318)? mem[542] : 
                 (N6320)? mem[544] : 
                 (N6322)? mem[546] : 
                 (N6324)? mem[548] : 
                 (N6326)? mem[550] : 
                 (N6328)? mem[552] : 
                 (N6330)? mem[554] : 
                 (N6332)? mem[556] : 
                 (N6334)? mem[558] : 
                 (N6336)? mem[560] : 
                 (N6338)? mem[562] : 
                 (N6340)? mem[564] : 
                 (N6342)? mem[566] : 
                 (N6344)? mem[568] : 
                 (N6346)? mem[570] : 
                 (N6348)? mem[572] : 
                 (N6350)? mem[574] : 
                 (N6352)? mem[576] : 
                 (N6354)? mem[578] : 
                 (N6356)? mem[580] : 
                 (N6358)? mem[582] : 
                 (N6360)? mem[584] : 
                 (N6362)? mem[586] : 
                 (N6364)? mem[588] : 
                 (N6366)? mem[590] : 
                 (N6368)? mem[592] : 
                 (N6370)? mem[594] : 
                 (N6372)? mem[596] : 
                 (N6374)? mem[598] : 
                 (N6376)? mem[600] : 
                 (N6378)? mem[602] : 
                 (N6380)? mem[604] : 
                 (N6382)? mem[606] : 
                 (N6384)? mem[608] : 
                 (N6386)? mem[610] : 
                 (N6388)? mem[612] : 
                 (N6390)? mem[614] : 
                 (N6392)? mem[616] : 
                 (N6394)? mem[618] : 
                 (N6396)? mem[620] : 
                 (N6398)? mem[622] : 
                 (N6400)? mem[624] : 
                 (N6402)? mem[626] : 
                 (N6404)? mem[628] : 
                 (N6406)? mem[630] : 
                 (N6408)? mem[632] : 
                 (N6410)? mem[634] : 
                 (N6412)? mem[636] : 
                 (N6414)? mem[638] : 
                 (N6416)? mem[640] : 
                 (N6418)? mem[642] : 
                 (N6420)? mem[644] : 
                 (N6422)? mem[646] : 
                 (N6424)? mem[648] : 
                 (N6426)? mem[650] : 
                 (N6428)? mem[652] : 
                 (N6430)? mem[654] : 
                 (N6432)? mem[656] : 
                 (N6434)? mem[658] : 
                 (N6436)? mem[660] : 
                 (N6438)? mem[662] : 
                 (N6440)? mem[664] : 
                 (N6442)? mem[666] : 
                 (N6444)? mem[668] : 
                 (N6446)? mem[670] : 
                 (N6448)? mem[672] : 
                 (N6450)? mem[674] : 
                 (N6452)? mem[676] : 
                 (N6454)? mem[678] : 
                 (N6456)? mem[680] : 
                 (N6458)? mem[682] : 
                 (N6460)? mem[684] : 
                 (N6462)? mem[686] : 
                 (N6464)? mem[688] : 
                 (N6466)? mem[690] : 
                 (N6468)? mem[692] : 
                 (N6470)? mem[694] : 
                 (N6472)? mem[696] : 
                 (N6474)? mem[698] : 
                 (N6476)? mem[700] : 
                 (N6478)? mem[702] : 
                 (N6480)? mem[704] : 
                 (N6482)? mem[706] : 
                 (N6484)? mem[708] : 
                 (N6486)? mem[710] : 
                 (N6488)? mem[712] : 
                 (N6490)? mem[714] : 
                 (N6492)? mem[716] : 
                 (N6494)? mem[718] : 
                 (N6496)? mem[720] : 
                 (N6498)? mem[722] : 
                 (N6500)? mem[724] : 
                 (N6502)? mem[726] : 
                 (N6504)? mem[728] : 
                 (N6506)? mem[730] : 
                 (N6508)? mem[732] : 
                 (N6510)? mem[734] : 
                 (N6512)? mem[736] : 
                 (N6514)? mem[738] : 
                 (N6516)? mem[740] : 
                 (N6518)? mem[742] : 
                 (N6520)? mem[744] : 
                 (N6522)? mem[746] : 
                 (N6524)? mem[748] : 
                 (N6526)? mem[750] : 
                 (N6528)? mem[752] : 
                 (N6530)? mem[754] : 
                 (N6532)? mem[756] : 
                 (N6534)? mem[758] : 
                 (N6536)? mem[760] : 
                 (N6538)? mem[762] : 
                 (N6540)? mem[764] : 
                 (N6542)? mem[766] : 
                 (N6544)? mem[768] : 
                 (N6546)? mem[770] : 
                 (N6548)? mem[772] : 
                 (N6550)? mem[774] : 
                 (N6552)? mem[776] : 
                 (N6554)? mem[778] : 
                 (N6556)? mem[780] : 
                 (N6558)? mem[782] : 
                 (N6560)? mem[784] : 
                 (N6562)? mem[786] : 
                 (N6564)? mem[788] : 
                 (N6566)? mem[790] : 
                 (N6568)? mem[792] : 
                 (N6570)? mem[794] : 
                 (N6572)? mem[796] : 
                 (N6574)? mem[798] : 
                 (N6576)? mem[800] : 
                 (N6578)? mem[802] : 
                 (N6580)? mem[804] : 
                 (N6582)? mem[806] : 
                 (N6584)? mem[808] : 
                 (N6586)? mem[810] : 
                 (N6588)? mem[812] : 
                 (N6590)? mem[814] : 
                 (N6592)? mem[816] : 
                 (N6594)? mem[818] : 
                 (N6596)? mem[820] : 
                 (N6598)? mem[822] : 
                 (N6600)? mem[824] : 
                 (N6602)? mem[826] : 
                 (N6604)? mem[828] : 
                 (N6606)? mem[830] : 
                 (N6608)? mem[832] : 
                 (N6610)? mem[834] : 
                 (N6612)? mem[836] : 
                 (N6614)? mem[838] : 
                 (N6616)? mem[840] : 
                 (N6618)? mem[842] : 
                 (N6620)? mem[844] : 
                 (N6622)? mem[846] : 
                 (N6624)? mem[848] : 
                 (N6626)? mem[850] : 
                 (N6628)? mem[852] : 
                 (N6630)? mem[854] : 
                 (N6632)? mem[856] : 
                 (N6634)? mem[858] : 
                 (N6636)? mem[860] : 
                 (N6638)? mem[862] : 
                 (N6640)? mem[864] : 
                 (N6642)? mem[866] : 
                 (N6644)? mem[868] : 
                 (N6646)? mem[870] : 
                 (N6648)? mem[872] : 
                 (N6650)? mem[874] : 
                 (N6652)? mem[876] : 
                 (N6654)? mem[878] : 
                 (N6656)? mem[880] : 
                 (N6658)? mem[882] : 
                 (N6660)? mem[884] : 
                 (N6662)? mem[886] : 
                 (N6664)? mem[888] : 
                 (N6666)? mem[890] : 
                 (N6668)? mem[892] : 
                 (N6670)? mem[894] : 
                 (N6672)? mem[896] : 
                 (N6674)? mem[898] : 
                 (N6676)? mem[900] : 
                 (N6678)? mem[902] : 
                 (N6680)? mem[904] : 
                 (N6682)? mem[906] : 
                 (N6684)? mem[908] : 
                 (N6686)? mem[910] : 
                 (N6688)? mem[912] : 
                 (N6690)? mem[914] : 
                 (N6692)? mem[916] : 
                 (N6694)? mem[918] : 
                 (N6696)? mem[920] : 
                 (N6698)? mem[922] : 
                 (N6700)? mem[924] : 
                 (N6702)? mem[926] : 
                 (N5879)? mem[928] : 
                 (N5881)? mem[930] : 
                 (N5883)? mem[932] : 
                 (N5885)? mem[934] : 
                 (N5887)? mem[936] : 
                 (N5889)? mem[938] : 
                 (N5891)? mem[940] : 
                 (N5893)? mem[942] : 
                 (N5895)? mem[944] : 
                 (N5897)? mem[946] : 
                 (N5899)? mem[948] : 
                 (N5901)? mem[950] : 
                 (N5903)? mem[952] : 
                 (N5905)? mem[954] : 
                 (N5907)? mem[956] : 
                 (N5909)? mem[958] : 
                 (N6720)? mem[960] : 
                 (N6722)? mem[962] : 
                 (N6724)? mem[964] : 
                 (N6726)? mem[966] : 
                 (N6728)? mem[968] : 
                 (N6730)? mem[970] : 
                 (N6732)? mem[972] : 
                 (N6734)? mem[974] : 
                 (N3612)? mem[976] : 
                 (N3614)? mem[978] : 
                 (N3616)? mem[980] : 
                 (N3618)? mem[982] : 
                 (N3620)? mem[984] : 
                 (N3622)? mem[986] : 
                 (N3624)? mem[988] : 
                 (N3626)? mem[990] : 
                 (N12081)? mem[992] : 
                 (N12083)? mem[994] : 
                 (N12085)? mem[996] : 
                 (N12087)? mem[998] : 
                 (N12089)? mem[1000] : 
                 (N12091)? mem[1002] : 
                 (N12093)? mem[1004] : 
                 (N12095)? mem[1006] : 
                 (N12097)? mem[1008] : 
                 (N12099)? mem[1010] : 
                 (N12101)? mem[1012] : 
                 (N12103)? mem[1014] : 
                 (N12105)? mem[1016] : 
                 (N12107)? mem[1018] : 
                 (N12109)? mem[1020] : 
                 (N12111)? mem[1022] : 1'b0;
  assign N7561 = (N7089)? mem[1] : 
                 (N7091)? mem[3] : 
                 (N7093)? mem[5] : 
                 (N7095)? mem[7] : 
                 (N7097)? mem[9] : 
                 (N7099)? mem[11] : 
                 (N7101)? mem[13] : 
                 (N7103)? mem[15] : 
                 (N7105)? mem[17] : 
                 (N7107)? mem[19] : 
                 (N7109)? mem[21] : 
                 (N7111)? mem[23] : 
                 (N7113)? mem[25] : 
                 (N7115)? mem[27] : 
                 (N7117)? mem[29] : 
                 (N7119)? mem[31] : 
                 (N7121)? mem[33] : 
                 (N7123)? mem[35] : 
                 (N7125)? mem[37] : 
                 (N7127)? mem[39] : 
                 (N7129)? mem[41] : 
                 (N7131)? mem[43] : 
                 (N7133)? mem[45] : 
                 (N7135)? mem[47] : 
                 (N7137)? mem[49] : 
                 (N7139)? mem[51] : 
                 (N7141)? mem[53] : 
                 (N7143)? mem[55] : 
                 (N7145)? mem[57] : 
                 (N7147)? mem[59] : 
                 (N7149)? mem[61] : 
                 (N7151)? mem[63] : 
                 (N7153)? mem[65] : 
                 (N7155)? mem[67] : 
                 (N7157)? mem[69] : 
                 (N7159)? mem[71] : 
                 (N7161)? mem[73] : 
                 (N7163)? mem[75] : 
                 (N7165)? mem[77] : 
                 (N7167)? mem[79] : 
                 (N7169)? mem[81] : 
                 (N7171)? mem[83] : 
                 (N7173)? mem[85] : 
                 (N7175)? mem[87] : 
                 (N7177)? mem[89] : 
                 (N7179)? mem[91] : 
                 (N7181)? mem[93] : 
                 (N7183)? mem[95] : 
                 (N7185)? mem[97] : 
                 (N7187)? mem[99] : 
                 (N7189)? mem[101] : 
                 (N7191)? mem[103] : 
                 (N7193)? mem[105] : 
                 (N7195)? mem[107] : 
                 (N7197)? mem[109] : 
                 (N7199)? mem[111] : 
                 (N7201)? mem[113] : 
                 (N7203)? mem[115] : 
                 (N7205)? mem[117] : 
                 (N7207)? mem[119] : 
                 (N7209)? mem[121] : 
                 (N7211)? mem[123] : 
                 (N7213)? mem[125] : 
                 (N7215)? mem[127] : 
                 (N7217)? mem[129] : 
                 (N7219)? mem[131] : 
                 (N7221)? mem[133] : 
                 (N7223)? mem[135] : 
                 (N7225)? mem[137] : 
                 (N7227)? mem[139] : 
                 (N7229)? mem[141] : 
                 (N7231)? mem[143] : 
                 (N7233)? mem[145] : 
                 (N7235)? mem[147] : 
                 (N7237)? mem[149] : 
                 (N7239)? mem[151] : 
                 (N7241)? mem[153] : 
                 (N7243)? mem[155] : 
                 (N7245)? mem[157] : 
                 (N7247)? mem[159] : 
                 (N7249)? mem[161] : 
                 (N7251)? mem[163] : 
                 (N7253)? mem[165] : 
                 (N7255)? mem[167] : 
                 (N7257)? mem[169] : 
                 (N7259)? mem[171] : 
                 (N7261)? mem[173] : 
                 (N7263)? mem[175] : 
                 (N7265)? mem[177] : 
                 (N7267)? mem[179] : 
                 (N7269)? mem[181] : 
                 (N7271)? mem[183] : 
                 (N7273)? mem[185] : 
                 (N7275)? mem[187] : 
                 (N7277)? mem[189] : 
                 (N7279)? mem[191] : 
                 (N7281)? mem[193] : 
                 (N7283)? mem[195] : 
                 (N7285)? mem[197] : 
                 (N7287)? mem[199] : 
                 (N7289)? mem[201] : 
                 (N7291)? mem[203] : 
                 (N7293)? mem[205] : 
                 (N7295)? mem[207] : 
                 (N7297)? mem[209] : 
                 (N7299)? mem[211] : 
                 (N7301)? mem[213] : 
                 (N7303)? mem[215] : 
                 (N7305)? mem[217] : 
                 (N7307)? mem[219] : 
                 (N7309)? mem[221] : 
                 (N7311)? mem[223] : 
                 (N7313)? mem[225] : 
                 (N7315)? mem[227] : 
                 (N7317)? mem[229] : 
                 (N7319)? mem[231] : 
                 (N7321)? mem[233] : 
                 (N7323)? mem[235] : 
                 (N7325)? mem[237] : 
                 (N7327)? mem[239] : 
                 (N7329)? mem[241] : 
                 (N7331)? mem[243] : 
                 (N7333)? mem[245] : 
                 (N7335)? mem[247] : 
                 (N7337)? mem[249] : 
                 (N7339)? mem[251] : 
                 (N7341)? mem[253] : 
                 (N7343)? mem[255] : 
                 (N7345)? mem[257] : 
                 (N7347)? mem[259] : 
                 (N7349)? mem[261] : 
                 (N7351)? mem[263] : 
                 (N7353)? mem[265] : 
                 (N7355)? mem[267] : 
                 (N7357)? mem[269] : 
                 (N7359)? mem[271] : 
                 (N7361)? mem[273] : 
                 (N7363)? mem[275] : 
                 (N7365)? mem[277] : 
                 (N7367)? mem[279] : 
                 (N7369)? mem[281] : 
                 (N7371)? mem[283] : 
                 (N7373)? mem[285] : 
                 (N7375)? mem[287] : 
                 (N7377)? mem[289] : 
                 (N7379)? mem[291] : 
                 (N7381)? mem[293] : 
                 (N7383)? mem[295] : 
                 (N7385)? mem[297] : 
                 (N7387)? mem[299] : 
                 (N7389)? mem[301] : 
                 (N7391)? mem[303] : 
                 (N7393)? mem[305] : 
                 (N7395)? mem[307] : 
                 (N7397)? mem[309] : 
                 (N7399)? mem[311] : 
                 (N7401)? mem[313] : 
                 (N7403)? mem[315] : 
                 (N7405)? mem[317] : 
                 (N7407)? mem[319] : 
                 (N7409)? mem[321] : 
                 (N7411)? mem[323] : 
                 (N7413)? mem[325] : 
                 (N7415)? mem[327] : 
                 (N7417)? mem[329] : 
                 (N7419)? mem[331] : 
                 (N7421)? mem[333] : 
                 (N7423)? mem[335] : 
                 (N7425)? mem[337] : 
                 (N7427)? mem[339] : 
                 (N7429)? mem[341] : 
                 (N7431)? mem[343] : 
                 (N7433)? mem[345] : 
                 (N7435)? mem[347] : 
                 (N7437)? mem[349] : 
                 (N7439)? mem[351] : 
                 (N7441)? mem[353] : 
                 (N7443)? mem[355] : 
                 (N7445)? mem[357] : 
                 (N7447)? mem[359] : 
                 (N7449)? mem[361] : 
                 (N7451)? mem[363] : 
                 (N7453)? mem[365] : 
                 (N7455)? mem[367] : 
                 (N7457)? mem[369] : 
                 (N7459)? mem[371] : 
                 (N7461)? mem[373] : 
                 (N7463)? mem[375] : 
                 (N7465)? mem[377] : 
                 (N7467)? mem[379] : 
                 (N7469)? mem[381] : 
                 (N7471)? mem[383] : 
                 (N7473)? mem[385] : 
                 (N7475)? mem[387] : 
                 (N7477)? mem[389] : 
                 (N7479)? mem[391] : 
                 (N7481)? mem[393] : 
                 (N7483)? mem[395] : 
                 (N7485)? mem[397] : 
                 (N7487)? mem[399] : 
                 (N7489)? mem[401] : 
                 (N7491)? mem[403] : 
                 (N7493)? mem[405] : 
                 (N7495)? mem[407] : 
                 (N7497)? mem[409] : 
                 (N7499)? mem[411] : 
                 (N7501)? mem[413] : 
                 (N7503)? mem[415] : 
                 (N7505)? mem[417] : 
                 (N7507)? mem[419] : 
                 (N7509)? mem[421] : 
                 (N7511)? mem[423] : 
                 (N7513)? mem[425] : 
                 (N7515)? mem[427] : 
                 (N7517)? mem[429] : 
                 (N7519)? mem[431] : 
                 (N7521)? mem[433] : 
                 (N7522)? mem[435] : 
                 (N7523)? mem[437] : 
                 (N7524)? mem[439] : 
                 (N7525)? mem[441] : 
                 (N7526)? mem[443] : 
                 (N7527)? mem[445] : 
                 (N7528)? mem[447] : 
                 (N7529)? mem[449] : 
                 (N7530)? mem[451] : 
                 (N7531)? mem[453] : 
                 (N7532)? mem[455] : 
                 (N7533)? mem[457] : 
                 (N7534)? mem[459] : 
                 (N7535)? mem[461] : 
                 (N7536)? mem[463] : 
                 (N7537)? mem[465] : 
                 (N7538)? mem[467] : 
                 (N7539)? mem[469] : 
                 (N7540)? mem[471] : 
                 (N7541)? mem[473] : 
                 (N7542)? mem[475] : 
                 (N7543)? mem[477] : 
                 (N7544)? mem[479] : 
                 (N7545)? mem[481] : 
                 (N7546)? mem[483] : 
                 (N7547)? mem[485] : 
                 (N7548)? mem[487] : 
                 (N7549)? mem[489] : 
                 (N7550)? mem[491] : 
                 (N7551)? mem[493] : 
                 (N7552)? mem[495] : 
                 (N7553)? mem[497] : 
                 (N7554)? mem[499] : 
                 (N7555)? mem[501] : 
                 (N7556)? mem[503] : 
                 (N7557)? mem[505] : 
                 (N7558)? mem[507] : 
                 (N7559)? mem[509] : 
                 (N7560)? mem[511] : 
                 (N7090)? mem[513] : 
                 (N7092)? mem[515] : 
                 (N7094)? mem[517] : 
                 (N7096)? mem[519] : 
                 (N7098)? mem[521] : 
                 (N7100)? mem[523] : 
                 (N7102)? mem[525] : 
                 (N7104)? mem[527] : 
                 (N7106)? mem[529] : 
                 (N7108)? mem[531] : 
                 (N7110)? mem[533] : 
                 (N7112)? mem[535] : 
                 (N7114)? mem[537] : 
                 (N7116)? mem[539] : 
                 (N7118)? mem[541] : 
                 (N7120)? mem[543] : 
                 (N7122)? mem[545] : 
                 (N7124)? mem[547] : 
                 (N7126)? mem[549] : 
                 (N7128)? mem[551] : 
                 (N7130)? mem[553] : 
                 (N7132)? mem[555] : 
                 (N7134)? mem[557] : 
                 (N7136)? mem[559] : 
                 (N7138)? mem[561] : 
                 (N7140)? mem[563] : 
                 (N7142)? mem[565] : 
                 (N7144)? mem[567] : 
                 (N7146)? mem[569] : 
                 (N7148)? mem[571] : 
                 (N7150)? mem[573] : 
                 (N7152)? mem[575] : 
                 (N7154)? mem[577] : 
                 (N7156)? mem[579] : 
                 (N7158)? mem[581] : 
                 (N7160)? mem[583] : 
                 (N7162)? mem[585] : 
                 (N7164)? mem[587] : 
                 (N7166)? mem[589] : 
                 (N7168)? mem[591] : 
                 (N7170)? mem[593] : 
                 (N7172)? mem[595] : 
                 (N7174)? mem[597] : 
                 (N7176)? mem[599] : 
                 (N7178)? mem[601] : 
                 (N7180)? mem[603] : 
                 (N7182)? mem[605] : 
                 (N7184)? mem[607] : 
                 (N7186)? mem[609] : 
                 (N7188)? mem[611] : 
                 (N7190)? mem[613] : 
                 (N7192)? mem[615] : 
                 (N7194)? mem[617] : 
                 (N7196)? mem[619] : 
                 (N7198)? mem[621] : 
                 (N7200)? mem[623] : 
                 (N7202)? mem[625] : 
                 (N7204)? mem[627] : 
                 (N7206)? mem[629] : 
                 (N7208)? mem[631] : 
                 (N7210)? mem[633] : 
                 (N7212)? mem[635] : 
                 (N7214)? mem[637] : 
                 (N7216)? mem[639] : 
                 (N7218)? mem[641] : 
                 (N7220)? mem[643] : 
                 (N7222)? mem[645] : 
                 (N7224)? mem[647] : 
                 (N7226)? mem[649] : 
                 (N7228)? mem[651] : 
                 (N7230)? mem[653] : 
                 (N7232)? mem[655] : 
                 (N7234)? mem[657] : 
                 (N7236)? mem[659] : 
                 (N7238)? mem[661] : 
                 (N7240)? mem[663] : 
                 (N7242)? mem[665] : 
                 (N7244)? mem[667] : 
                 (N7246)? mem[669] : 
                 (N7248)? mem[671] : 
                 (N7250)? mem[673] : 
                 (N7252)? mem[675] : 
                 (N7254)? mem[677] : 
                 (N7256)? mem[679] : 
                 (N7258)? mem[681] : 
                 (N7260)? mem[683] : 
                 (N7262)? mem[685] : 
                 (N7264)? mem[687] : 
                 (N7266)? mem[689] : 
                 (N7268)? mem[691] : 
                 (N7270)? mem[693] : 
                 (N7272)? mem[695] : 
                 (N7274)? mem[697] : 
                 (N7276)? mem[699] : 
                 (N7278)? mem[701] : 
                 (N7280)? mem[703] : 
                 (N7282)? mem[705] : 
                 (N7284)? mem[707] : 
                 (N7286)? mem[709] : 
                 (N7288)? mem[711] : 
                 (N7290)? mem[713] : 
                 (N7292)? mem[715] : 
                 (N7294)? mem[717] : 
                 (N7296)? mem[719] : 
                 (N7298)? mem[721] : 
                 (N7300)? mem[723] : 
                 (N7302)? mem[725] : 
                 (N7304)? mem[727] : 
                 (N7306)? mem[729] : 
                 (N7308)? mem[731] : 
                 (N7310)? mem[733] : 
                 (N7312)? mem[735] : 
                 (N7314)? mem[737] : 
                 (N7316)? mem[739] : 
                 (N7318)? mem[741] : 
                 (N7320)? mem[743] : 
                 (N7322)? mem[745] : 
                 (N7324)? mem[747] : 
                 (N7326)? mem[749] : 
                 (N7328)? mem[751] : 
                 (N7330)? mem[753] : 
                 (N7332)? mem[755] : 
                 (N7334)? mem[757] : 
                 (N7336)? mem[759] : 
                 (N7338)? mem[761] : 
                 (N7340)? mem[763] : 
                 (N7342)? mem[765] : 
                 (N7344)? mem[767] : 
                 (N7346)? mem[769] : 
                 (N7348)? mem[771] : 
                 (N7350)? mem[773] : 
                 (N7352)? mem[775] : 
                 (N7354)? mem[777] : 
                 (N7356)? mem[779] : 
                 (N7358)? mem[781] : 
                 (N7360)? mem[783] : 
                 (N7362)? mem[785] : 
                 (N7364)? mem[787] : 
                 (N7366)? mem[789] : 
                 (N7368)? mem[791] : 
                 (N7370)? mem[793] : 
                 (N7372)? mem[795] : 
                 (N7374)? mem[797] : 
                 (N7376)? mem[799] : 
                 (N7378)? mem[801] : 
                 (N7380)? mem[803] : 
                 (N7382)? mem[805] : 
                 (N7384)? mem[807] : 
                 (N7386)? mem[809] : 
                 (N7388)? mem[811] : 
                 (N7390)? mem[813] : 
                 (N7392)? mem[815] : 
                 (N7394)? mem[817] : 
                 (N7396)? mem[819] : 
                 (N7398)? mem[821] : 
                 (N7400)? mem[823] : 
                 (N7402)? mem[825] : 
                 (N7404)? mem[827] : 
                 (N7406)? mem[829] : 
                 (N7408)? mem[831] : 
                 (N7410)? mem[833] : 
                 (N7412)? mem[835] : 
                 (N7414)? mem[837] : 
                 (N7416)? mem[839] : 
                 (N7418)? mem[841] : 
                 (N7420)? mem[843] : 
                 (N7422)? mem[845] : 
                 (N7424)? mem[847] : 
                 (N7426)? mem[849] : 
                 (N7428)? mem[851] : 
                 (N7430)? mem[853] : 
                 (N7432)? mem[855] : 
                 (N7434)? mem[857] : 
                 (N7436)? mem[859] : 
                 (N7438)? mem[861] : 
                 (N7440)? mem[863] : 
                 (N7442)? mem[865] : 
                 (N7444)? mem[867] : 
                 (N7446)? mem[869] : 
                 (N7448)? mem[871] : 
                 (N7450)? mem[873] : 
                 (N7452)? mem[875] : 
                 (N7454)? mem[877] : 
                 (N7456)? mem[879] : 
                 (N7458)? mem[881] : 
                 (N7460)? mem[883] : 
                 (N7462)? mem[885] : 
                 (N7464)? mem[887] : 
                 (N7466)? mem[889] : 
                 (N7468)? mem[891] : 
                 (N7470)? mem[893] : 
                 (N7472)? mem[895] : 
                 (N7474)? mem[897] : 
                 (N7476)? mem[899] : 
                 (N7478)? mem[901] : 
                 (N7480)? mem[903] : 
                 (N7482)? mem[905] : 
                 (N7484)? mem[907] : 
                 (N7486)? mem[909] : 
                 (N7488)? mem[911] : 
                 (N7490)? mem[913] : 
                 (N7492)? mem[915] : 
                 (N7494)? mem[917] : 
                 (N7496)? mem[919] : 
                 (N7498)? mem[921] : 
                 (N7500)? mem[923] : 
                 (N7502)? mem[925] : 
                 (N7504)? mem[927] : 
                 (N7506)? mem[929] : 
                 (N7508)? mem[931] : 
                 (N7510)? mem[933] : 
                 (N7512)? mem[935] : 
                 (N7514)? mem[937] : 
                 (N7516)? mem[939] : 
                 (N7518)? mem[941] : 
                 (N7520)? mem[943] : 
                 (N4501)? mem[945] : 
                 (N4503)? mem[947] : 
                 (N4505)? mem[949] : 
                 (N4507)? mem[951] : 
                 (N4509)? mem[953] : 
                 (N4511)? mem[955] : 
                 (N4513)? mem[957] : 
                 (N4515)? mem[959] : 
                 (N6720)? mem[961] : 
                 (N6722)? mem[963] : 
                 (N6724)? mem[965] : 
                 (N6726)? mem[967] : 
                 (N6728)? mem[969] : 
                 (N6730)? mem[971] : 
                 (N6732)? mem[973] : 
                 (N6734)? mem[975] : 
                 (N3612)? mem[977] : 
                 (N3614)? mem[979] : 
                 (N3616)? mem[981] : 
                 (N3618)? mem[983] : 
                 (N3620)? mem[985] : 
                 (N3622)? mem[987] : 
                 (N3624)? mem[989] : 
                 (N3626)? mem[991] : 
                 (N12081)? mem[993] : 
                 (N12083)? mem[995] : 
                 (N12085)? mem[997] : 
                 (N12087)? mem[999] : 
                 (N12089)? mem[1001] : 
                 (N12091)? mem[1003] : 
                 (N12093)? mem[1005] : 
                 (N12095)? mem[1007] : 
                 (N12097)? mem[1009] : 
                 (N12099)? mem[1011] : 
                 (N12101)? mem[1013] : 
                 (N12103)? mem[1015] : 
                 (N12105)? mem[1017] : 
                 (N12107)? mem[1019] : 
                 (N12109)? mem[1021] : 
                 (N12111)? mem[1023] : 1'b0;
  assign N8266 = (N7818)? mem[0] : 
                 (N7820)? mem[2] : 
                 (N7822)? mem[4] : 
                 (N7824)? mem[6] : 
                 (N7826)? mem[8] : 
                 (N7828)? mem[10] : 
                 (N7830)? mem[12] : 
                 (N7832)? mem[14] : 
                 (N7834)? mem[16] : 
                 (N7836)? mem[18] : 
                 (N7838)? mem[20] : 
                 (N7840)? mem[22] : 
                 (N7842)? mem[24] : 
                 (N7844)? mem[26] : 
                 (N7846)? mem[28] : 
                 (N7848)? mem[30] : 
                 (N7850)? mem[32] : 
                 (N7852)? mem[34] : 
                 (N7854)? mem[36] : 
                 (N7856)? mem[38] : 
                 (N7858)? mem[40] : 
                 (N7860)? mem[42] : 
                 (N7862)? mem[44] : 
                 (N7864)? mem[46] : 
                 (N7866)? mem[48] : 
                 (N7868)? mem[50] : 
                 (N7870)? mem[52] : 
                 (N7872)? mem[54] : 
                 (N7874)? mem[56] : 
                 (N7876)? mem[58] : 
                 (N7878)? mem[60] : 
                 (N7880)? mem[62] : 
                 (N7882)? mem[64] : 
                 (N7884)? mem[66] : 
                 (N7886)? mem[68] : 
                 (N7888)? mem[70] : 
                 (N7890)? mem[72] : 
                 (N7892)? mem[74] : 
                 (N7894)? mem[76] : 
                 (N7896)? mem[78] : 
                 (N7898)? mem[80] : 
                 (N7900)? mem[82] : 
                 (N7902)? mem[84] : 
                 (N7904)? mem[86] : 
                 (N7906)? mem[88] : 
                 (N7908)? mem[90] : 
                 (N7910)? mem[92] : 
                 (N7912)? mem[94] : 
                 (N7914)? mem[96] : 
                 (N7916)? mem[98] : 
                 (N7918)? mem[100] : 
                 (N7920)? mem[102] : 
                 (N7922)? mem[104] : 
                 (N7924)? mem[106] : 
                 (N7926)? mem[108] : 
                 (N7928)? mem[110] : 
                 (N7930)? mem[112] : 
                 (N7932)? mem[114] : 
                 (N7934)? mem[116] : 
                 (N7936)? mem[118] : 
                 (N7938)? mem[120] : 
                 (N7940)? mem[122] : 
                 (N7942)? mem[124] : 
                 (N7944)? mem[126] : 
                 (N7946)? mem[128] : 
                 (N7948)? mem[130] : 
                 (N7950)? mem[132] : 
                 (N7952)? mem[134] : 
                 (N7954)? mem[136] : 
                 (N7956)? mem[138] : 
                 (N7958)? mem[140] : 
                 (N7960)? mem[142] : 
                 (N7962)? mem[144] : 
                 (N7964)? mem[146] : 
                 (N7966)? mem[148] : 
                 (N7968)? mem[150] : 
                 (N7970)? mem[152] : 
                 (N7972)? mem[154] : 
                 (N7974)? mem[156] : 
                 (N7976)? mem[158] : 
                 (N7978)? mem[160] : 
                 (N7980)? mem[162] : 
                 (N7982)? mem[164] : 
                 (N7984)? mem[166] : 
                 (N7986)? mem[168] : 
                 (N7988)? mem[170] : 
                 (N7990)? mem[172] : 
                 (N7992)? mem[174] : 
                 (N7994)? mem[176] : 
                 (N7996)? mem[178] : 
                 (N7998)? mem[180] : 
                 (N8000)? mem[182] : 
                 (N8002)? mem[184] : 
                 (N8004)? mem[186] : 
                 (N8006)? mem[188] : 
                 (N8008)? mem[190] : 
                 (N8010)? mem[192] : 
                 (N8012)? mem[194] : 
                 (N8014)? mem[196] : 
                 (N8016)? mem[198] : 
                 (N8018)? mem[200] : 
                 (N8020)? mem[202] : 
                 (N8022)? mem[204] : 
                 (N8024)? mem[206] : 
                 (N8026)? mem[208] : 
                 (N8028)? mem[210] : 
                 (N8030)? mem[212] : 
                 (N8032)? mem[214] : 
                 (N8034)? mem[216] : 
                 (N8036)? mem[218] : 
                 (N8038)? mem[220] : 
                 (N8040)? mem[222] : 
                 (N8042)? mem[224] : 
                 (N8044)? mem[226] : 
                 (N8046)? mem[228] : 
                 (N8048)? mem[230] : 
                 (N8050)? mem[232] : 
                 (N8052)? mem[234] : 
                 (N8054)? mem[236] : 
                 (N8056)? mem[238] : 
                 (N8058)? mem[240] : 
                 (N8060)? mem[242] : 
                 (N8062)? mem[244] : 
                 (N8064)? mem[246] : 
                 (N8066)? mem[248] : 
                 (N8068)? mem[250] : 
                 (N8070)? mem[252] : 
                 (N8072)? mem[254] : 
                 (N8074)? mem[256] : 
                 (N8076)? mem[258] : 
                 (N8078)? mem[260] : 
                 (N8080)? mem[262] : 
                 (N8082)? mem[264] : 
                 (N8084)? mem[266] : 
                 (N8086)? mem[268] : 
                 (N8088)? mem[270] : 
                 (N8090)? mem[272] : 
                 (N8092)? mem[274] : 
                 (N8094)? mem[276] : 
                 (N8096)? mem[278] : 
                 (N8098)? mem[280] : 
                 (N8100)? mem[282] : 
                 (N8102)? mem[284] : 
                 (N8104)? mem[286] : 
                 (N8106)? mem[288] : 
                 (N8108)? mem[290] : 
                 (N8110)? mem[292] : 
                 (N8112)? mem[294] : 
                 (N8114)? mem[296] : 
                 (N8116)? mem[298] : 
                 (N8118)? mem[300] : 
                 (N8120)? mem[302] : 
                 (N8122)? mem[304] : 
                 (N8124)? mem[306] : 
                 (N8126)? mem[308] : 
                 (N8128)? mem[310] : 
                 (N8130)? mem[312] : 
                 (N8132)? mem[314] : 
                 (N8134)? mem[316] : 
                 (N8136)? mem[318] : 
                 (N8138)? mem[320] : 
                 (N8140)? mem[322] : 
                 (N8142)? mem[324] : 
                 (N8144)? mem[326] : 
                 (N8146)? mem[328] : 
                 (N8148)? mem[330] : 
                 (N8150)? mem[332] : 
                 (N8152)? mem[334] : 
                 (N8154)? mem[336] : 
                 (N8156)? mem[338] : 
                 (N8158)? mem[340] : 
                 (N8160)? mem[342] : 
                 (N8162)? mem[344] : 
                 (N8164)? mem[346] : 
                 (N8166)? mem[348] : 
                 (N8168)? mem[350] : 
                 (N8170)? mem[352] : 
                 (N8172)? mem[354] : 
                 (N8174)? mem[356] : 
                 (N8176)? mem[358] : 
                 (N8178)? mem[360] : 
                 (N8180)? mem[362] : 
                 (N8182)? mem[364] : 
                 (N8184)? mem[366] : 
                 (N8186)? mem[368] : 
                 (N8188)? mem[370] : 
                 (N8190)? mem[372] : 
                 (N8192)? mem[374] : 
                 (N8194)? mem[376] : 
                 (N8196)? mem[378] : 
                 (N8198)? mem[380] : 
                 (N8200)? mem[382] : 
                 (N8202)? mem[384] : 
                 (N8203)? mem[386] : 
                 (N8204)? mem[388] : 
                 (N8205)? mem[390] : 
                 (N8206)? mem[392] : 
                 (N8207)? mem[394] : 
                 (N8208)? mem[396] : 
                 (N8209)? mem[398] : 
                 (N8210)? mem[400] : 
                 (N8211)? mem[402] : 
                 (N8212)? mem[404] : 
                 (N8213)? mem[406] : 
                 (N8214)? mem[408] : 
                 (N8215)? mem[410] : 
                 (N8216)? mem[412] : 
                 (N8217)? mem[414] : 
                 (N8218)? mem[416] : 
                 (N8219)? mem[418] : 
                 (N8220)? mem[420] : 
                 (N8221)? mem[422] : 
                 (N8222)? mem[424] : 
                 (N8223)? mem[426] : 
                 (N8224)? mem[428] : 
                 (N8225)? mem[430] : 
                 (N8226)? mem[432] : 
                 (N8227)? mem[434] : 
                 (N8228)? mem[436] : 
                 (N8229)? mem[438] : 
                 (N8230)? mem[440] : 
                 (N8231)? mem[442] : 
                 (N8232)? mem[444] : 
                 (N8233)? mem[446] : 
                 (N8234)? mem[448] : 
                 (N8235)? mem[450] : 
                 (N8236)? mem[452] : 
                 (N8237)? mem[454] : 
                 (N8238)? mem[456] : 
                 (N8239)? mem[458] : 
                 (N8240)? mem[460] : 
                 (N8241)? mem[462] : 
                 (N8242)? mem[464] : 
                 (N8243)? mem[466] : 
                 (N8244)? mem[468] : 
                 (N8245)? mem[470] : 
                 (N8246)? mem[472] : 
                 (N8247)? mem[474] : 
                 (N8248)? mem[476] : 
                 (N8249)? mem[478] : 
                 (N8250)? mem[480] : 
                 (N8251)? mem[482] : 
                 (N8252)? mem[484] : 
                 (N8253)? mem[486] : 
                 (N8254)? mem[488] : 
                 (N8255)? mem[490] : 
                 (N8256)? mem[492] : 
                 (N8257)? mem[494] : 
                 (N8258)? mem[496] : 
                 (N8259)? mem[498] : 
                 (N8260)? mem[500] : 
                 (N8261)? mem[502] : 
                 (N8262)? mem[504] : 
                 (N8263)? mem[506] : 
                 (N8264)? mem[508] : 
                 (N8265)? mem[510] : 
                 (N7819)? mem[512] : 
                 (N7821)? mem[514] : 
                 (N7823)? mem[516] : 
                 (N7825)? mem[518] : 
                 (N7827)? mem[520] : 
                 (N7829)? mem[522] : 
                 (N7831)? mem[524] : 
                 (N7833)? mem[526] : 
                 (N7835)? mem[528] : 
                 (N7837)? mem[530] : 
                 (N7839)? mem[532] : 
                 (N7841)? mem[534] : 
                 (N7843)? mem[536] : 
                 (N7845)? mem[538] : 
                 (N7847)? mem[540] : 
                 (N7849)? mem[542] : 
                 (N7851)? mem[544] : 
                 (N7853)? mem[546] : 
                 (N7855)? mem[548] : 
                 (N7857)? mem[550] : 
                 (N7859)? mem[552] : 
                 (N7861)? mem[554] : 
                 (N7863)? mem[556] : 
                 (N7865)? mem[558] : 
                 (N7867)? mem[560] : 
                 (N7869)? mem[562] : 
                 (N7871)? mem[564] : 
                 (N7873)? mem[566] : 
                 (N7875)? mem[568] : 
                 (N7877)? mem[570] : 
                 (N7879)? mem[572] : 
                 (N7881)? mem[574] : 
                 (N7883)? mem[576] : 
                 (N7885)? mem[578] : 
                 (N7887)? mem[580] : 
                 (N7889)? mem[582] : 
                 (N7891)? mem[584] : 
                 (N7893)? mem[586] : 
                 (N7895)? mem[588] : 
                 (N7897)? mem[590] : 
                 (N7899)? mem[592] : 
                 (N7901)? mem[594] : 
                 (N7903)? mem[596] : 
                 (N7905)? mem[598] : 
                 (N7907)? mem[600] : 
                 (N7909)? mem[602] : 
                 (N7911)? mem[604] : 
                 (N7913)? mem[606] : 
                 (N7915)? mem[608] : 
                 (N7917)? mem[610] : 
                 (N7919)? mem[612] : 
                 (N7921)? mem[614] : 
                 (N7923)? mem[616] : 
                 (N7925)? mem[618] : 
                 (N7927)? mem[620] : 
                 (N7929)? mem[622] : 
                 (N7931)? mem[624] : 
                 (N7933)? mem[626] : 
                 (N7935)? mem[628] : 
                 (N7937)? mem[630] : 
                 (N7939)? mem[632] : 
                 (N7941)? mem[634] : 
                 (N7943)? mem[636] : 
                 (N7945)? mem[638] : 
                 (N7947)? mem[640] : 
                 (N7949)? mem[642] : 
                 (N7951)? mem[644] : 
                 (N7953)? mem[646] : 
                 (N7955)? mem[648] : 
                 (N7957)? mem[650] : 
                 (N7959)? mem[652] : 
                 (N7961)? mem[654] : 
                 (N7963)? mem[656] : 
                 (N7965)? mem[658] : 
                 (N7967)? mem[660] : 
                 (N7969)? mem[662] : 
                 (N7971)? mem[664] : 
                 (N7973)? mem[666] : 
                 (N7975)? mem[668] : 
                 (N7977)? mem[670] : 
                 (N7979)? mem[672] : 
                 (N7981)? mem[674] : 
                 (N7983)? mem[676] : 
                 (N7985)? mem[678] : 
                 (N7987)? mem[680] : 
                 (N7989)? mem[682] : 
                 (N7991)? mem[684] : 
                 (N7993)? mem[686] : 
                 (N7995)? mem[688] : 
                 (N7997)? mem[690] : 
                 (N7999)? mem[692] : 
                 (N8001)? mem[694] : 
                 (N8003)? mem[696] : 
                 (N8005)? mem[698] : 
                 (N8007)? mem[700] : 
                 (N8009)? mem[702] : 
                 (N8011)? mem[704] : 
                 (N8013)? mem[706] : 
                 (N8015)? mem[708] : 
                 (N8017)? mem[710] : 
                 (N8019)? mem[712] : 
                 (N8021)? mem[714] : 
                 (N8023)? mem[716] : 
                 (N8025)? mem[718] : 
                 (N8027)? mem[720] : 
                 (N8029)? mem[722] : 
                 (N8031)? mem[724] : 
                 (N8033)? mem[726] : 
                 (N8035)? mem[728] : 
                 (N8037)? mem[730] : 
                 (N8039)? mem[732] : 
                 (N8041)? mem[734] : 
                 (N8043)? mem[736] : 
                 (N8045)? mem[738] : 
                 (N8047)? mem[740] : 
                 (N8049)? mem[742] : 
                 (N8051)? mem[744] : 
                 (N8053)? mem[746] : 
                 (N8055)? mem[748] : 
                 (N8057)? mem[750] : 
                 (N8059)? mem[752] : 
                 (N8061)? mem[754] : 
                 (N8063)? mem[756] : 
                 (N8065)? mem[758] : 
                 (N8067)? mem[760] : 
                 (N8069)? mem[762] : 
                 (N8071)? mem[764] : 
                 (N8073)? mem[766] : 
                 (N8075)? mem[768] : 
                 (N8077)? mem[770] : 
                 (N8079)? mem[772] : 
                 (N8081)? mem[774] : 
                 (N8083)? mem[776] : 
                 (N8085)? mem[778] : 
                 (N8087)? mem[780] : 
                 (N8089)? mem[782] : 
                 (N8091)? mem[784] : 
                 (N8093)? mem[786] : 
                 (N8095)? mem[788] : 
                 (N8097)? mem[790] : 
                 (N8099)? mem[792] : 
                 (N8101)? mem[794] : 
                 (N8103)? mem[796] : 
                 (N8105)? mem[798] : 
                 (N8107)? mem[800] : 
                 (N8109)? mem[802] : 
                 (N8111)? mem[804] : 
                 (N8113)? mem[806] : 
                 (N8115)? mem[808] : 
                 (N8117)? mem[810] : 
                 (N8119)? mem[812] : 
                 (N8121)? mem[814] : 
                 (N8123)? mem[816] : 
                 (N8125)? mem[818] : 
                 (N8127)? mem[820] : 
                 (N8129)? mem[822] : 
                 (N8131)? mem[824] : 
                 (N8133)? mem[826] : 
                 (N8135)? mem[828] : 
                 (N8137)? mem[830] : 
                 (N8139)? mem[832] : 
                 (N8141)? mem[834] : 
                 (N8143)? mem[836] : 
                 (N8145)? mem[838] : 
                 (N8147)? mem[840] : 
                 (N8149)? mem[842] : 
                 (N8151)? mem[844] : 
                 (N8153)? mem[846] : 
                 (N8155)? mem[848] : 
                 (N8157)? mem[850] : 
                 (N8159)? mem[852] : 
                 (N8161)? mem[854] : 
                 (N8163)? mem[856] : 
                 (N8165)? mem[858] : 
                 (N8167)? mem[860] : 
                 (N8169)? mem[862] : 
                 (N8171)? mem[864] : 
                 (N8173)? mem[866] : 
                 (N8175)? mem[868] : 
                 (N8177)? mem[870] : 
                 (N8179)? mem[872] : 
                 (N8181)? mem[874] : 
                 (N8183)? mem[876] : 
                 (N8185)? mem[878] : 
                 (N8187)? mem[880] : 
                 (N8189)? mem[882] : 
                 (N8191)? mem[884] : 
                 (N8193)? mem[886] : 
                 (N8195)? mem[888] : 
                 (N8197)? mem[890] : 
                 (N8199)? mem[892] : 
                 (N8201)? mem[894] : 
                 (N7474)? mem[896] : 
                 (N7476)? mem[898] : 
                 (N7478)? mem[900] : 
                 (N7480)? mem[902] : 
                 (N7482)? mem[904] : 
                 (N7484)? mem[906] : 
                 (N7486)? mem[908] : 
                 (N7488)? mem[910] : 
                 (N7490)? mem[912] : 
                 (N7492)? mem[914] : 
                 (N7494)? mem[916] : 
                 (N7496)? mem[918] : 
                 (N7498)? mem[920] : 
                 (N7500)? mem[922] : 
                 (N7502)? mem[924] : 
                 (N7504)? mem[926] : 
                 (N7506)? mem[928] : 
                 (N7508)? mem[930] : 
                 (N7510)? mem[932] : 
                 (N7512)? mem[934] : 
                 (N7514)? mem[936] : 
                 (N7516)? mem[938] : 
                 (N7518)? mem[940] : 
                 (N7520)? mem[942] : 
                 (N4501)? mem[944] : 
                 (N4503)? mem[946] : 
                 (N4505)? mem[948] : 
                 (N4507)? mem[950] : 
                 (N4509)? mem[952] : 
                 (N4511)? mem[954] : 
                 (N4513)? mem[956] : 
                 (N4515)? mem[958] : 
                 (N6720)? mem[960] : 
                 (N6722)? mem[962] : 
                 (N6724)? mem[964] : 
                 (N6726)? mem[966] : 
                 (N6728)? mem[968] : 
                 (N6730)? mem[970] : 
                 (N6732)? mem[972] : 
                 (N6734)? mem[974] : 
                 (N3612)? mem[976] : 
                 (N3614)? mem[978] : 
                 (N3616)? mem[980] : 
                 (N3618)? mem[982] : 
                 (N3620)? mem[984] : 
                 (N3622)? mem[986] : 
                 (N3624)? mem[988] : 
                 (N3626)? mem[990] : 
                 (N12081)? mem[992] : 
                 (N12083)? mem[994] : 
                 (N12085)? mem[996] : 
                 (N12087)? mem[998] : 
                 (N12089)? mem[1000] : 
                 (N12091)? mem[1002] : 
                 (N12093)? mem[1004] : 
                 (N12095)? mem[1006] : 
                 (N12097)? mem[1008] : 
                 (N12099)? mem[1010] : 
                 (N12101)? mem[1012] : 
                 (N12103)? mem[1014] : 
                 (N12105)? mem[1016] : 
                 (N12107)? mem[1018] : 
                 (N12109)? mem[1020] : 
                 (N12111)? mem[1022] : 1'b0;
  assign N9036 = (N8572)? mem[1] : 
                 (N8574)? mem[3] : 
                 (N8576)? mem[5] : 
                 (N8578)? mem[7] : 
                 (N8580)? mem[9] : 
                 (N8582)? mem[11] : 
                 (N8584)? mem[13] : 
                 (N8586)? mem[15] : 
                 (N8588)? mem[17] : 
                 (N8590)? mem[19] : 
                 (N8592)? mem[21] : 
                 (N8594)? mem[23] : 
                 (N8596)? mem[25] : 
                 (N8598)? mem[27] : 
                 (N8600)? mem[29] : 
                 (N8602)? mem[31] : 
                 (N8604)? mem[33] : 
                 (N8606)? mem[35] : 
                 (N8608)? mem[37] : 
                 (N8610)? mem[39] : 
                 (N8612)? mem[41] : 
                 (N8614)? mem[43] : 
                 (N8616)? mem[45] : 
                 (N8618)? mem[47] : 
                 (N8620)? mem[49] : 
                 (N8622)? mem[51] : 
                 (N8624)? mem[53] : 
                 (N8626)? mem[55] : 
                 (N8628)? mem[57] : 
                 (N8630)? mem[59] : 
                 (N8632)? mem[61] : 
                 (N8634)? mem[63] : 
                 (N8636)? mem[65] : 
                 (N8638)? mem[67] : 
                 (N8640)? mem[69] : 
                 (N8642)? mem[71] : 
                 (N8644)? mem[73] : 
                 (N8646)? mem[75] : 
                 (N8648)? mem[77] : 
                 (N8650)? mem[79] : 
                 (N8652)? mem[81] : 
                 (N8654)? mem[83] : 
                 (N8656)? mem[85] : 
                 (N8658)? mem[87] : 
                 (N8660)? mem[89] : 
                 (N8662)? mem[91] : 
                 (N8664)? mem[93] : 
                 (N8666)? mem[95] : 
                 (N8668)? mem[97] : 
                 (N8670)? mem[99] : 
                 (N8672)? mem[101] : 
                 (N8674)? mem[103] : 
                 (N8676)? mem[105] : 
                 (N8678)? mem[107] : 
                 (N8680)? mem[109] : 
                 (N8682)? mem[111] : 
                 (N8684)? mem[113] : 
                 (N8686)? mem[115] : 
                 (N8688)? mem[117] : 
                 (N8690)? mem[119] : 
                 (N8692)? mem[121] : 
                 (N8694)? mem[123] : 
                 (N8696)? mem[125] : 
                 (N8698)? mem[127] : 
                 (N8700)? mem[129] : 
                 (N8702)? mem[131] : 
                 (N8704)? mem[133] : 
                 (N8706)? mem[135] : 
                 (N8708)? mem[137] : 
                 (N8710)? mem[139] : 
                 (N8712)? mem[141] : 
                 (N8714)? mem[143] : 
                 (N8716)? mem[145] : 
                 (N8718)? mem[147] : 
                 (N8720)? mem[149] : 
                 (N8722)? mem[151] : 
                 (N8724)? mem[153] : 
                 (N8726)? mem[155] : 
                 (N8728)? mem[157] : 
                 (N8730)? mem[159] : 
                 (N8732)? mem[161] : 
                 (N8734)? mem[163] : 
                 (N8736)? mem[165] : 
                 (N8738)? mem[167] : 
                 (N8740)? mem[169] : 
                 (N8742)? mem[171] : 
                 (N8744)? mem[173] : 
                 (N8746)? mem[175] : 
                 (N8748)? mem[177] : 
                 (N8750)? mem[179] : 
                 (N8752)? mem[181] : 
                 (N8754)? mem[183] : 
                 (N8756)? mem[185] : 
                 (N8758)? mem[187] : 
                 (N8760)? mem[189] : 
                 (N8762)? mem[191] : 
                 (N8764)? mem[193] : 
                 (N8766)? mem[195] : 
                 (N8768)? mem[197] : 
                 (N8770)? mem[199] : 
                 (N8772)? mem[201] : 
                 (N8774)? mem[203] : 
                 (N8776)? mem[205] : 
                 (N8778)? mem[207] : 
                 (N8780)? mem[209] : 
                 (N8782)? mem[211] : 
                 (N8784)? mem[213] : 
                 (N8786)? mem[215] : 
                 (N8788)? mem[217] : 
                 (N8790)? mem[219] : 
                 (N8792)? mem[221] : 
                 (N8794)? mem[223] : 
                 (N8796)? mem[225] : 
                 (N8798)? mem[227] : 
                 (N8800)? mem[229] : 
                 (N8802)? mem[231] : 
                 (N8804)? mem[233] : 
                 (N8806)? mem[235] : 
                 (N8808)? mem[237] : 
                 (N8810)? mem[239] : 
                 (N8812)? mem[241] : 
                 (N8814)? mem[243] : 
                 (N8816)? mem[245] : 
                 (N8818)? mem[247] : 
                 (N8820)? mem[249] : 
                 (N8822)? mem[251] : 
                 (N8824)? mem[253] : 
                 (N8826)? mem[255] : 
                 (N8828)? mem[257] : 
                 (N8830)? mem[259] : 
                 (N8832)? mem[261] : 
                 (N8834)? mem[263] : 
                 (N8836)? mem[265] : 
                 (N8838)? mem[267] : 
                 (N8840)? mem[269] : 
                 (N8842)? mem[271] : 
                 (N8844)? mem[273] : 
                 (N8846)? mem[275] : 
                 (N8848)? mem[277] : 
                 (N8850)? mem[279] : 
                 (N8852)? mem[281] : 
                 (N8854)? mem[283] : 
                 (N8856)? mem[285] : 
                 (N8858)? mem[287] : 
                 (N8860)? mem[289] : 
                 (N8862)? mem[291] : 
                 (N8864)? mem[293] : 
                 (N8866)? mem[295] : 
                 (N8868)? mem[297] : 
                 (N8870)? mem[299] : 
                 (N8872)? mem[301] : 
                 (N8874)? mem[303] : 
                 (N8876)? mem[305] : 
                 (N8878)? mem[307] : 
                 (N8880)? mem[309] : 
                 (N8882)? mem[311] : 
                 (N8884)? mem[313] : 
                 (N8886)? mem[315] : 
                 (N8888)? mem[317] : 
                 (N8890)? mem[319] : 
                 (N8892)? mem[321] : 
                 (N8894)? mem[323] : 
                 (N8896)? mem[325] : 
                 (N8898)? mem[327] : 
                 (N8900)? mem[329] : 
                 (N8902)? mem[331] : 
                 (N8904)? mem[333] : 
                 (N8906)? mem[335] : 
                 (N8908)? mem[337] : 
                 (N8910)? mem[339] : 
                 (N8912)? mem[341] : 
                 (N8914)? mem[343] : 
                 (N8916)? mem[345] : 
                 (N8918)? mem[347] : 
                 (N8920)? mem[349] : 
                 (N8922)? mem[351] : 
                 (N8924)? mem[353] : 
                 (N8926)? mem[355] : 
                 (N8928)? mem[357] : 
                 (N8930)? mem[359] : 
                 (N8932)? mem[361] : 
                 (N8934)? mem[363] : 
                 (N8936)? mem[365] : 
                 (N8938)? mem[367] : 
                 (N8940)? mem[369] : 
                 (N8942)? mem[371] : 
                 (N8944)? mem[373] : 
                 (N8946)? mem[375] : 
                 (N8948)? mem[377] : 
                 (N8950)? mem[379] : 
                 (N8952)? mem[381] : 
                 (N8954)? mem[383] : 
                 (N8956)? mem[385] : 
                 (N8958)? mem[387] : 
                 (N8960)? mem[389] : 
                 (N8962)? mem[391] : 
                 (N8964)? mem[393] : 
                 (N8966)? mem[395] : 
                 (N8968)? mem[397] : 
                 (N8970)? mem[399] : 
                 (N8972)? mem[401] : 
                 (N8973)? mem[403] : 
                 (N8974)? mem[405] : 
                 (N8975)? mem[407] : 
                 (N8976)? mem[409] : 
                 (N8977)? mem[411] : 
                 (N8978)? mem[413] : 
                 (N8979)? mem[415] : 
                 (N8980)? mem[417] : 
                 (N8982)? mem[419] : 
                 (N8984)? mem[421] : 
                 (N8986)? mem[423] : 
                 (N8988)? mem[425] : 
                 (N8990)? mem[427] : 
                 (N8992)? mem[429] : 
                 (N8994)? mem[431] : 
                 (N8996)? mem[433] : 
                 (N8997)? mem[435] : 
                 (N8998)? mem[437] : 
                 (N8999)? mem[439] : 
                 (N9000)? mem[441] : 
                 (N9001)? mem[443] : 
                 (N9002)? mem[445] : 
                 (N9003)? mem[447] : 
                 (N9004)? mem[449] : 
                 (N9005)? mem[451] : 
                 (N9006)? mem[453] : 
                 (N9007)? mem[455] : 
                 (N9008)? mem[457] : 
                 (N9009)? mem[459] : 
                 (N9010)? mem[461] : 
                 (N9011)? mem[463] : 
                 (N9012)? mem[465] : 
                 (N9013)? mem[467] : 
                 (N9014)? mem[469] : 
                 (N9015)? mem[471] : 
                 (N9016)? mem[473] : 
                 (N9017)? mem[475] : 
                 (N9018)? mem[477] : 
                 (N9019)? mem[479] : 
                 (N9020)? mem[481] : 
                 (N9021)? mem[483] : 
                 (N9022)? mem[485] : 
                 (N9023)? mem[487] : 
                 (N9024)? mem[489] : 
                 (N9025)? mem[491] : 
                 (N9026)? mem[493] : 
                 (N9027)? mem[495] : 
                 (N9028)? mem[497] : 
                 (N9029)? mem[499] : 
                 (N9030)? mem[501] : 
                 (N9031)? mem[503] : 
                 (N9032)? mem[505] : 
                 (N9033)? mem[507] : 
                 (N9034)? mem[509] : 
                 (N9035)? mem[511] : 
                 (N8573)? mem[513] : 
                 (N8575)? mem[515] : 
                 (N8577)? mem[517] : 
                 (N8579)? mem[519] : 
                 (N8581)? mem[521] : 
                 (N8583)? mem[523] : 
                 (N8585)? mem[525] : 
                 (N8587)? mem[527] : 
                 (N8589)? mem[529] : 
                 (N8591)? mem[531] : 
                 (N8593)? mem[533] : 
                 (N8595)? mem[535] : 
                 (N8597)? mem[537] : 
                 (N8599)? mem[539] : 
                 (N8601)? mem[541] : 
                 (N8603)? mem[543] : 
                 (N8605)? mem[545] : 
                 (N8607)? mem[547] : 
                 (N8609)? mem[549] : 
                 (N8611)? mem[551] : 
                 (N8613)? mem[553] : 
                 (N8615)? mem[555] : 
                 (N8617)? mem[557] : 
                 (N8619)? mem[559] : 
                 (N8621)? mem[561] : 
                 (N8623)? mem[563] : 
                 (N8625)? mem[565] : 
                 (N8627)? mem[567] : 
                 (N8629)? mem[569] : 
                 (N8631)? mem[571] : 
                 (N8633)? mem[573] : 
                 (N8635)? mem[575] : 
                 (N8637)? mem[577] : 
                 (N8639)? mem[579] : 
                 (N8641)? mem[581] : 
                 (N8643)? mem[583] : 
                 (N8645)? mem[585] : 
                 (N8647)? mem[587] : 
                 (N8649)? mem[589] : 
                 (N8651)? mem[591] : 
                 (N8653)? mem[593] : 
                 (N8655)? mem[595] : 
                 (N8657)? mem[597] : 
                 (N8659)? mem[599] : 
                 (N8661)? mem[601] : 
                 (N8663)? mem[603] : 
                 (N8665)? mem[605] : 
                 (N8667)? mem[607] : 
                 (N8669)? mem[609] : 
                 (N8671)? mem[611] : 
                 (N8673)? mem[613] : 
                 (N8675)? mem[615] : 
                 (N8677)? mem[617] : 
                 (N8679)? mem[619] : 
                 (N8681)? mem[621] : 
                 (N8683)? mem[623] : 
                 (N8685)? mem[625] : 
                 (N8687)? mem[627] : 
                 (N8689)? mem[629] : 
                 (N8691)? mem[631] : 
                 (N8693)? mem[633] : 
                 (N8695)? mem[635] : 
                 (N8697)? mem[637] : 
                 (N8699)? mem[639] : 
                 (N8701)? mem[641] : 
                 (N8703)? mem[643] : 
                 (N8705)? mem[645] : 
                 (N8707)? mem[647] : 
                 (N8709)? mem[649] : 
                 (N8711)? mem[651] : 
                 (N8713)? mem[653] : 
                 (N8715)? mem[655] : 
                 (N8717)? mem[657] : 
                 (N8719)? mem[659] : 
                 (N8721)? mem[661] : 
                 (N8723)? mem[663] : 
                 (N8725)? mem[665] : 
                 (N8727)? mem[667] : 
                 (N8729)? mem[669] : 
                 (N8731)? mem[671] : 
                 (N8733)? mem[673] : 
                 (N8735)? mem[675] : 
                 (N8737)? mem[677] : 
                 (N8739)? mem[679] : 
                 (N8741)? mem[681] : 
                 (N8743)? mem[683] : 
                 (N8745)? mem[685] : 
                 (N8747)? mem[687] : 
                 (N8749)? mem[689] : 
                 (N8751)? mem[691] : 
                 (N8753)? mem[693] : 
                 (N8755)? mem[695] : 
                 (N8757)? mem[697] : 
                 (N8759)? mem[699] : 
                 (N8761)? mem[701] : 
                 (N8763)? mem[703] : 
                 (N8765)? mem[705] : 
                 (N8767)? mem[707] : 
                 (N8769)? mem[709] : 
                 (N8771)? mem[711] : 
                 (N8773)? mem[713] : 
                 (N8775)? mem[715] : 
                 (N8777)? mem[717] : 
                 (N8779)? mem[719] : 
                 (N8781)? mem[721] : 
                 (N8783)? mem[723] : 
                 (N8785)? mem[725] : 
                 (N8787)? mem[727] : 
                 (N8789)? mem[729] : 
                 (N8791)? mem[731] : 
                 (N8793)? mem[733] : 
                 (N8795)? mem[735] : 
                 (N8797)? mem[737] : 
                 (N8799)? mem[739] : 
                 (N8801)? mem[741] : 
                 (N8803)? mem[743] : 
                 (N8805)? mem[745] : 
                 (N8807)? mem[747] : 
                 (N8809)? mem[749] : 
                 (N8811)? mem[751] : 
                 (N8813)? mem[753] : 
                 (N8815)? mem[755] : 
                 (N8817)? mem[757] : 
                 (N8819)? mem[759] : 
                 (N8821)? mem[761] : 
                 (N8823)? mem[763] : 
                 (N8825)? mem[765] : 
                 (N8827)? mem[767] : 
                 (N8829)? mem[769] : 
                 (N8831)? mem[771] : 
                 (N8833)? mem[773] : 
                 (N8835)? mem[775] : 
                 (N8837)? mem[777] : 
                 (N8839)? mem[779] : 
                 (N8841)? mem[781] : 
                 (N8843)? mem[783] : 
                 (N8845)? mem[785] : 
                 (N8847)? mem[787] : 
                 (N8849)? mem[789] : 
                 (N8851)? mem[791] : 
                 (N8853)? mem[793] : 
                 (N8855)? mem[795] : 
                 (N8857)? mem[797] : 
                 (N8859)? mem[799] : 
                 (N8861)? mem[801] : 
                 (N8863)? mem[803] : 
                 (N8865)? mem[805] : 
                 (N8867)? mem[807] : 
                 (N8869)? mem[809] : 
                 (N8871)? mem[811] : 
                 (N8873)? mem[813] : 
                 (N8875)? mem[815] : 
                 (N8877)? mem[817] : 
                 (N8879)? mem[819] : 
                 (N8881)? mem[821] : 
                 (N8883)? mem[823] : 
                 (N8885)? mem[825] : 
                 (N8887)? mem[827] : 
                 (N8889)? mem[829] : 
                 (N8891)? mem[831] : 
                 (N8893)? mem[833] : 
                 (N8895)? mem[835] : 
                 (N8897)? mem[837] : 
                 (N8899)? mem[839] : 
                 (N8901)? mem[841] : 
                 (N8903)? mem[843] : 
                 (N8905)? mem[845] : 
                 (N8907)? mem[847] : 
                 (N8909)? mem[849] : 
                 (N8911)? mem[851] : 
                 (N8913)? mem[853] : 
                 (N8915)? mem[855] : 
                 (N8917)? mem[857] : 
                 (N8919)? mem[859] : 
                 (N8921)? mem[861] : 
                 (N8923)? mem[863] : 
                 (N8925)? mem[865] : 
                 (N8927)? mem[867] : 
                 (N8929)? mem[869] : 
                 (N8931)? mem[871] : 
                 (N8933)? mem[873] : 
                 (N8935)? mem[875] : 
                 (N8937)? mem[877] : 
                 (N8939)? mem[879] : 
                 (N8941)? mem[881] : 
                 (N8943)? mem[883] : 
                 (N8945)? mem[885] : 
                 (N8947)? mem[887] : 
                 (N8949)? mem[889] : 
                 (N8951)? mem[891] : 
                 (N8953)? mem[893] : 
                 (N8955)? mem[895] : 
                 (N8957)? mem[897] : 
                 (N8959)? mem[899] : 
                 (N8961)? mem[901] : 
                 (N8963)? mem[903] : 
                 (N8965)? mem[905] : 
                 (N8967)? mem[907] : 
                 (N8969)? mem[909] : 
                 (N8971)? mem[911] : 
                 (N3548)? mem[913] : 
                 (N3550)? mem[915] : 
                 (N3552)? mem[917] : 
                 (N3554)? mem[919] : 
                 (N3556)? mem[921] : 
                 (N3558)? mem[923] : 
                 (N3560)? mem[925] : 
                 (N3562)? mem[927] : 
                 (N8981)? mem[929] : 
                 (N8983)? mem[931] : 
                 (N8985)? mem[933] : 
                 (N8987)? mem[935] : 
                 (N8989)? mem[937] : 
                 (N8991)? mem[939] : 
                 (N8993)? mem[941] : 
                 (N8995)? mem[943] : 
                 (N3580)? mem[945] : 
                 (N3582)? mem[947] : 
                 (N3584)? mem[949] : 
                 (N3586)? mem[951] : 
                 (N3588)? mem[953] : 
                 (N3590)? mem[955] : 
                 (N3592)? mem[957] : 
                 (N3594)? mem[959] : 
                 (N6720)? mem[961] : 
                 (N6722)? mem[963] : 
                 (N6724)? mem[965] : 
                 (N6726)? mem[967] : 
                 (N6728)? mem[969] : 
                 (N6730)? mem[971] : 
                 (N6732)? mem[973] : 
                 (N6734)? mem[975] : 
                 (N3612)? mem[977] : 
                 (N3614)? mem[979] : 
                 (N3616)? mem[981] : 
                 (N3618)? mem[983] : 
                 (N3620)? mem[985] : 
                 (N3622)? mem[987] : 
                 (N3624)? mem[989] : 
                 (N3626)? mem[991] : 
                 (N12081)? mem[993] : 
                 (N12083)? mem[995] : 
                 (N12085)? mem[997] : 
                 (N12087)? mem[999] : 
                 (N12089)? mem[1001] : 
                 (N12091)? mem[1003] : 
                 (N12093)? mem[1005] : 
                 (N12095)? mem[1007] : 
                 (N12097)? mem[1009] : 
                 (N12099)? mem[1011] : 
                 (N12101)? mem[1013] : 
                 (N12103)? mem[1015] : 
                 (N12105)? mem[1017] : 
                 (N12107)? mem[1019] : 
                 (N12109)? mem[1021] : 
                 (N12111)? mem[1023] : 1'b0;
  assign N9741 = (N9293)? mem[0] : 
                 (N9295)? mem[2] : 
                 (N9297)? mem[4] : 
                 (N9299)? mem[6] : 
                 (N9301)? mem[8] : 
                 (N9303)? mem[10] : 
                 (N9305)? mem[12] : 
                 (N9307)? mem[14] : 
                 (N9309)? mem[16] : 
                 (N9311)? mem[18] : 
                 (N9313)? mem[20] : 
                 (N9315)? mem[22] : 
                 (N9317)? mem[24] : 
                 (N9319)? mem[26] : 
                 (N9321)? mem[28] : 
                 (N9323)? mem[30] : 
                 (N9325)? mem[32] : 
                 (N9327)? mem[34] : 
                 (N9329)? mem[36] : 
                 (N9331)? mem[38] : 
                 (N9333)? mem[40] : 
                 (N9335)? mem[42] : 
                 (N9337)? mem[44] : 
                 (N9339)? mem[46] : 
                 (N9341)? mem[48] : 
                 (N9343)? mem[50] : 
                 (N9345)? mem[52] : 
                 (N9347)? mem[54] : 
                 (N9349)? mem[56] : 
                 (N9351)? mem[58] : 
                 (N9353)? mem[60] : 
                 (N9355)? mem[62] : 
                 (N9357)? mem[64] : 
                 (N9359)? mem[66] : 
                 (N9361)? mem[68] : 
                 (N9363)? mem[70] : 
                 (N9365)? mem[72] : 
                 (N9367)? mem[74] : 
                 (N9369)? mem[76] : 
                 (N9371)? mem[78] : 
                 (N9373)? mem[80] : 
                 (N9375)? mem[82] : 
                 (N9377)? mem[84] : 
                 (N9379)? mem[86] : 
                 (N9381)? mem[88] : 
                 (N9383)? mem[90] : 
                 (N9385)? mem[92] : 
                 (N9387)? mem[94] : 
                 (N9389)? mem[96] : 
                 (N9391)? mem[98] : 
                 (N9393)? mem[100] : 
                 (N9395)? mem[102] : 
                 (N9397)? mem[104] : 
                 (N9399)? mem[106] : 
                 (N9401)? mem[108] : 
                 (N9403)? mem[110] : 
                 (N9405)? mem[112] : 
                 (N9407)? mem[114] : 
                 (N9409)? mem[116] : 
                 (N9411)? mem[118] : 
                 (N9413)? mem[120] : 
                 (N9415)? mem[122] : 
                 (N9417)? mem[124] : 
                 (N9419)? mem[126] : 
                 (N9421)? mem[128] : 
                 (N9423)? mem[130] : 
                 (N9425)? mem[132] : 
                 (N9427)? mem[134] : 
                 (N9429)? mem[136] : 
                 (N9431)? mem[138] : 
                 (N9433)? mem[140] : 
                 (N9435)? mem[142] : 
                 (N9437)? mem[144] : 
                 (N9439)? mem[146] : 
                 (N9441)? mem[148] : 
                 (N9443)? mem[150] : 
                 (N9445)? mem[152] : 
                 (N9447)? mem[154] : 
                 (N9449)? mem[156] : 
                 (N9451)? mem[158] : 
                 (N9453)? mem[160] : 
                 (N9455)? mem[162] : 
                 (N9457)? mem[164] : 
                 (N9459)? mem[166] : 
                 (N9461)? mem[168] : 
                 (N9463)? mem[170] : 
                 (N9465)? mem[172] : 
                 (N9467)? mem[174] : 
                 (N9469)? mem[176] : 
                 (N9471)? mem[178] : 
                 (N9473)? mem[180] : 
                 (N9475)? mem[182] : 
                 (N9477)? mem[184] : 
                 (N9479)? mem[186] : 
                 (N9481)? mem[188] : 
                 (N9483)? mem[190] : 
                 (N9485)? mem[192] : 
                 (N9487)? mem[194] : 
                 (N9489)? mem[196] : 
                 (N9491)? mem[198] : 
                 (N9493)? mem[200] : 
                 (N9495)? mem[202] : 
                 (N9497)? mem[204] : 
                 (N9499)? mem[206] : 
                 (N9501)? mem[208] : 
                 (N9503)? mem[210] : 
                 (N9505)? mem[212] : 
                 (N9507)? mem[214] : 
                 (N9509)? mem[216] : 
                 (N9511)? mem[218] : 
                 (N9513)? mem[220] : 
                 (N9515)? mem[222] : 
                 (N9517)? mem[224] : 
                 (N9519)? mem[226] : 
                 (N9521)? mem[228] : 
                 (N9523)? mem[230] : 
                 (N9525)? mem[232] : 
                 (N9527)? mem[234] : 
                 (N9529)? mem[236] : 
                 (N9531)? mem[238] : 
                 (N9533)? mem[240] : 
                 (N9535)? mem[242] : 
                 (N9537)? mem[244] : 
                 (N9539)? mem[246] : 
                 (N9541)? mem[248] : 
                 (N9543)? mem[250] : 
                 (N9545)? mem[252] : 
                 (N9547)? mem[254] : 
                 (N9549)? mem[256] : 
                 (N9551)? mem[258] : 
                 (N9553)? mem[260] : 
                 (N9555)? mem[262] : 
                 (N9557)? mem[264] : 
                 (N9559)? mem[266] : 
                 (N9561)? mem[268] : 
                 (N9563)? mem[270] : 
                 (N9565)? mem[272] : 
                 (N9567)? mem[274] : 
                 (N9569)? mem[276] : 
                 (N9571)? mem[278] : 
                 (N9573)? mem[280] : 
                 (N9575)? mem[282] : 
                 (N9577)? mem[284] : 
                 (N9579)? mem[286] : 
                 (N9581)? mem[288] : 
                 (N9583)? mem[290] : 
                 (N9585)? mem[292] : 
                 (N9587)? mem[294] : 
                 (N9589)? mem[296] : 
                 (N9591)? mem[298] : 
                 (N9593)? mem[300] : 
                 (N9595)? mem[302] : 
                 (N9597)? mem[304] : 
                 (N9599)? mem[306] : 
                 (N9601)? mem[308] : 
                 (N9603)? mem[310] : 
                 (N9605)? mem[312] : 
                 (N9607)? mem[314] : 
                 (N9609)? mem[316] : 
                 (N9611)? mem[318] : 
                 (N9613)? mem[320] : 
                 (N9615)? mem[322] : 
                 (N9617)? mem[324] : 
                 (N9619)? mem[326] : 
                 (N9621)? mem[328] : 
                 (N9623)? mem[330] : 
                 (N9625)? mem[332] : 
                 (N9627)? mem[334] : 
                 (N9629)? mem[336] : 
                 (N9631)? mem[338] : 
                 (N9633)? mem[340] : 
                 (N9635)? mem[342] : 
                 (N9637)? mem[344] : 
                 (N9639)? mem[346] : 
                 (N9641)? mem[348] : 
                 (N9643)? mem[350] : 
                 (N9645)? mem[352] : 
                 (N9647)? mem[354] : 
                 (N9649)? mem[356] : 
                 (N9651)? mem[358] : 
                 (N9653)? mem[360] : 
                 (N9655)? mem[362] : 
                 (N9657)? mem[364] : 
                 (N9659)? mem[366] : 
                 (N9661)? mem[368] : 
                 (N9663)? mem[370] : 
                 (N9665)? mem[372] : 
                 (N9667)? mem[374] : 
                 (N9669)? mem[376] : 
                 (N9671)? mem[378] : 
                 (N9673)? mem[380] : 
                 (N9675)? mem[382] : 
                 (N9677)? mem[384] : 
                 (N9678)? mem[386] : 
                 (N9679)? mem[388] : 
                 (N9680)? mem[390] : 
                 (N9681)? mem[392] : 
                 (N9682)? mem[394] : 
                 (N9683)? mem[396] : 
                 (N9684)? mem[398] : 
                 (N9685)? mem[400] : 
                 (N9686)? mem[402] : 
                 (N9687)? mem[404] : 
                 (N9688)? mem[406] : 
                 (N9689)? mem[408] : 
                 (N9690)? mem[410] : 
                 (N9691)? mem[412] : 
                 (N9692)? mem[414] : 
                 (N9693)? mem[416] : 
                 (N9694)? mem[418] : 
                 (N9695)? mem[420] : 
                 (N9696)? mem[422] : 
                 (N9697)? mem[424] : 
                 (N9698)? mem[426] : 
                 (N9699)? mem[428] : 
                 (N9700)? mem[430] : 
                 (N9701)? mem[432] : 
                 (N9702)? mem[434] : 
                 (N9703)? mem[436] : 
                 (N9704)? mem[438] : 
                 (N9705)? mem[440] : 
                 (N9706)? mem[442] : 
                 (N9707)? mem[444] : 
                 (N9708)? mem[446] : 
                 (N9709)? mem[448] : 
                 (N9710)? mem[450] : 
                 (N9711)? mem[452] : 
                 (N9712)? mem[454] : 
                 (N9713)? mem[456] : 
                 (N9714)? mem[458] : 
                 (N9715)? mem[460] : 
                 (N9716)? mem[462] : 
                 (N9717)? mem[464] : 
                 (N9718)? mem[466] : 
                 (N9719)? mem[468] : 
                 (N9720)? mem[470] : 
                 (N9721)? mem[472] : 
                 (N9722)? mem[474] : 
                 (N9723)? mem[476] : 
                 (N9724)? mem[478] : 
                 (N9725)? mem[480] : 
                 (N9726)? mem[482] : 
                 (N9727)? mem[484] : 
                 (N9728)? mem[486] : 
                 (N9729)? mem[488] : 
                 (N9730)? mem[490] : 
                 (N9731)? mem[492] : 
                 (N9732)? mem[494] : 
                 (N9733)? mem[496] : 
                 (N9734)? mem[498] : 
                 (N9735)? mem[500] : 
                 (N9736)? mem[502] : 
                 (N9737)? mem[504] : 
                 (N9738)? mem[506] : 
                 (N9739)? mem[508] : 
                 (N9740)? mem[510] : 
                 (N9294)? mem[512] : 
                 (N9296)? mem[514] : 
                 (N9298)? mem[516] : 
                 (N9300)? mem[518] : 
                 (N9302)? mem[520] : 
                 (N9304)? mem[522] : 
                 (N9306)? mem[524] : 
                 (N9308)? mem[526] : 
                 (N9310)? mem[528] : 
                 (N9312)? mem[530] : 
                 (N9314)? mem[532] : 
                 (N9316)? mem[534] : 
                 (N9318)? mem[536] : 
                 (N9320)? mem[538] : 
                 (N9322)? mem[540] : 
                 (N9324)? mem[542] : 
                 (N9326)? mem[544] : 
                 (N9328)? mem[546] : 
                 (N9330)? mem[548] : 
                 (N9332)? mem[550] : 
                 (N9334)? mem[552] : 
                 (N9336)? mem[554] : 
                 (N9338)? mem[556] : 
                 (N9340)? mem[558] : 
                 (N9342)? mem[560] : 
                 (N9344)? mem[562] : 
                 (N9346)? mem[564] : 
                 (N9348)? mem[566] : 
                 (N9350)? mem[568] : 
                 (N9352)? mem[570] : 
                 (N9354)? mem[572] : 
                 (N9356)? mem[574] : 
                 (N9358)? mem[576] : 
                 (N9360)? mem[578] : 
                 (N9362)? mem[580] : 
                 (N9364)? mem[582] : 
                 (N9366)? mem[584] : 
                 (N9368)? mem[586] : 
                 (N9370)? mem[588] : 
                 (N9372)? mem[590] : 
                 (N9374)? mem[592] : 
                 (N9376)? mem[594] : 
                 (N9378)? mem[596] : 
                 (N9380)? mem[598] : 
                 (N9382)? mem[600] : 
                 (N9384)? mem[602] : 
                 (N9386)? mem[604] : 
                 (N9388)? mem[606] : 
                 (N9390)? mem[608] : 
                 (N9392)? mem[610] : 
                 (N9394)? mem[612] : 
                 (N9396)? mem[614] : 
                 (N9398)? mem[616] : 
                 (N9400)? mem[618] : 
                 (N9402)? mem[620] : 
                 (N9404)? mem[622] : 
                 (N9406)? mem[624] : 
                 (N9408)? mem[626] : 
                 (N9410)? mem[628] : 
                 (N9412)? mem[630] : 
                 (N9414)? mem[632] : 
                 (N9416)? mem[634] : 
                 (N9418)? mem[636] : 
                 (N9420)? mem[638] : 
                 (N9422)? mem[640] : 
                 (N9424)? mem[642] : 
                 (N9426)? mem[644] : 
                 (N9428)? mem[646] : 
                 (N9430)? mem[648] : 
                 (N9432)? mem[650] : 
                 (N9434)? mem[652] : 
                 (N9436)? mem[654] : 
                 (N9438)? mem[656] : 
                 (N9440)? mem[658] : 
                 (N9442)? mem[660] : 
                 (N9444)? mem[662] : 
                 (N9446)? mem[664] : 
                 (N9448)? mem[666] : 
                 (N9450)? mem[668] : 
                 (N9452)? mem[670] : 
                 (N9454)? mem[672] : 
                 (N9456)? mem[674] : 
                 (N9458)? mem[676] : 
                 (N9460)? mem[678] : 
                 (N9462)? mem[680] : 
                 (N9464)? mem[682] : 
                 (N9466)? mem[684] : 
                 (N9468)? mem[686] : 
                 (N9470)? mem[688] : 
                 (N9472)? mem[690] : 
                 (N9474)? mem[692] : 
                 (N9476)? mem[694] : 
                 (N9478)? mem[696] : 
                 (N9480)? mem[698] : 
                 (N9482)? mem[700] : 
                 (N9484)? mem[702] : 
                 (N9486)? mem[704] : 
                 (N9488)? mem[706] : 
                 (N9490)? mem[708] : 
                 (N9492)? mem[710] : 
                 (N9494)? mem[712] : 
                 (N9496)? mem[714] : 
                 (N9498)? mem[716] : 
                 (N9500)? mem[718] : 
                 (N9502)? mem[720] : 
                 (N9504)? mem[722] : 
                 (N9506)? mem[724] : 
                 (N9508)? mem[726] : 
                 (N9510)? mem[728] : 
                 (N9512)? mem[730] : 
                 (N9514)? mem[732] : 
                 (N9516)? mem[734] : 
                 (N9518)? mem[736] : 
                 (N9520)? mem[738] : 
                 (N9522)? mem[740] : 
                 (N9524)? mem[742] : 
                 (N9526)? mem[744] : 
                 (N9528)? mem[746] : 
                 (N9530)? mem[748] : 
                 (N9532)? mem[750] : 
                 (N9534)? mem[752] : 
                 (N9536)? mem[754] : 
                 (N9538)? mem[756] : 
                 (N9540)? mem[758] : 
                 (N9542)? mem[760] : 
                 (N9544)? mem[762] : 
                 (N9546)? mem[764] : 
                 (N9548)? mem[766] : 
                 (N9550)? mem[768] : 
                 (N9552)? mem[770] : 
                 (N9554)? mem[772] : 
                 (N9556)? mem[774] : 
                 (N9558)? mem[776] : 
                 (N9560)? mem[778] : 
                 (N9562)? mem[780] : 
                 (N9564)? mem[782] : 
                 (N9566)? mem[784] : 
                 (N9568)? mem[786] : 
                 (N9570)? mem[788] : 
                 (N9572)? mem[790] : 
                 (N9574)? mem[792] : 
                 (N9576)? mem[794] : 
                 (N9578)? mem[796] : 
                 (N9580)? mem[798] : 
                 (N9582)? mem[800] : 
                 (N9584)? mem[802] : 
                 (N9586)? mem[804] : 
                 (N9588)? mem[806] : 
                 (N9590)? mem[808] : 
                 (N9592)? mem[810] : 
                 (N9594)? mem[812] : 
                 (N9596)? mem[814] : 
                 (N9598)? mem[816] : 
                 (N9600)? mem[818] : 
                 (N9602)? mem[820] : 
                 (N9604)? mem[822] : 
                 (N9606)? mem[824] : 
                 (N9608)? mem[826] : 
                 (N9610)? mem[828] : 
                 (N9612)? mem[830] : 
                 (N9614)? mem[832] : 
                 (N9616)? mem[834] : 
                 (N9618)? mem[836] : 
                 (N9620)? mem[838] : 
                 (N9622)? mem[840] : 
                 (N9624)? mem[842] : 
                 (N9626)? mem[844] : 
                 (N9628)? mem[846] : 
                 (N9630)? mem[848] : 
                 (N9632)? mem[850] : 
                 (N9634)? mem[852] : 
                 (N9636)? mem[854] : 
                 (N9638)? mem[856] : 
                 (N9640)? mem[858] : 
                 (N9642)? mem[860] : 
                 (N9644)? mem[862] : 
                 (N9646)? mem[864] : 
                 (N9648)? mem[866] : 
                 (N9650)? mem[868] : 
                 (N9652)? mem[870] : 
                 (N9654)? mem[872] : 
                 (N9656)? mem[874] : 
                 (N9658)? mem[876] : 
                 (N9660)? mem[878] : 
                 (N9662)? mem[880] : 
                 (N9664)? mem[882] : 
                 (N9666)? mem[884] : 
                 (N9668)? mem[886] : 
                 (N9670)? mem[888] : 
                 (N9672)? mem[890] : 
                 (N9674)? mem[892] : 
                 (N9676)? mem[894] : 
                 (N8957)? mem[896] : 
                 (N8959)? mem[898] : 
                 (N8961)? mem[900] : 
                 (N8963)? mem[902] : 
                 (N8965)? mem[904] : 
                 (N8967)? mem[906] : 
                 (N8969)? mem[908] : 
                 (N8971)? mem[910] : 
                 (N3548)? mem[912] : 
                 (N3550)? mem[914] : 
                 (N3552)? mem[916] : 
                 (N3554)? mem[918] : 
                 (N3556)? mem[920] : 
                 (N3558)? mem[922] : 
                 (N3560)? mem[924] : 
                 (N3562)? mem[926] : 
                 (N8981)? mem[928] : 
                 (N8983)? mem[930] : 
                 (N8985)? mem[932] : 
                 (N8987)? mem[934] : 
                 (N8989)? mem[936] : 
                 (N8991)? mem[938] : 
                 (N8993)? mem[940] : 
                 (N8995)? mem[942] : 
                 (N3580)? mem[944] : 
                 (N3582)? mem[946] : 
                 (N3584)? mem[948] : 
                 (N3586)? mem[950] : 
                 (N3588)? mem[952] : 
                 (N3590)? mem[954] : 
                 (N3592)? mem[956] : 
                 (N3594)? mem[958] : 
                 (N6720)? mem[960] : 
                 (N6722)? mem[962] : 
                 (N6724)? mem[964] : 
                 (N6726)? mem[966] : 
                 (N6728)? mem[968] : 
                 (N6730)? mem[970] : 
                 (N6732)? mem[972] : 
                 (N6734)? mem[974] : 
                 (N3612)? mem[976] : 
                 (N3614)? mem[978] : 
                 (N3616)? mem[980] : 
                 (N3618)? mem[982] : 
                 (N3620)? mem[984] : 
                 (N3622)? mem[986] : 
                 (N3624)? mem[988] : 
                 (N3626)? mem[990] : 
                 (N12081)? mem[992] : 
                 (N12083)? mem[994] : 
                 (N12085)? mem[996] : 
                 (N12087)? mem[998] : 
                 (N12089)? mem[1000] : 
                 (N12091)? mem[1002] : 
                 (N12093)? mem[1004] : 
                 (N12095)? mem[1006] : 
                 (N12097)? mem[1008] : 
                 (N12099)? mem[1010] : 
                 (N12101)? mem[1012] : 
                 (N12103)? mem[1014] : 
                 (N12105)? mem[1016] : 
                 (N12107)? mem[1018] : 
                 (N12109)? mem[1020] : 
                 (N12111)? mem[1022] : 1'b0;
  assign N11087 = (N10607)? mem[1] : 
                  (N10609)? mem[3] : 
                  (N10611)? mem[5] : 
                  (N10613)? mem[7] : 
                  (N10615)? mem[9] : 
                  (N10617)? mem[11] : 
                  (N10619)? mem[13] : 
                  (N10621)? mem[15] : 
                  (N10623)? mem[17] : 
                  (N10625)? mem[19] : 
                  (N10627)? mem[21] : 
                  (N10629)? mem[23] : 
                  (N10631)? mem[25] : 
                  (N10633)? mem[27] : 
                  (N10635)? mem[29] : 
                  (N10637)? mem[31] : 
                  (N10639)? mem[33] : 
                  (N10641)? mem[35] : 
                  (N10643)? mem[37] : 
                  (N10645)? mem[39] : 
                  (N10647)? mem[41] : 
                  (N10649)? mem[43] : 
                  (N10651)? mem[45] : 
                  (N10653)? mem[47] : 
                  (N10655)? mem[49] : 
                  (N10657)? mem[51] : 
                  (N10659)? mem[53] : 
                  (N10661)? mem[55] : 
                  (N10663)? mem[57] : 
                  (N10665)? mem[59] : 
                  (N10667)? mem[61] : 
                  (N10669)? mem[63] : 
                  (N10671)? mem[65] : 
                  (N10673)? mem[67] : 
                  (N10675)? mem[69] : 
                  (N10677)? mem[71] : 
                  (N10679)? mem[73] : 
                  (N10681)? mem[75] : 
                  (N10683)? mem[77] : 
                  (N10685)? mem[79] : 
                  (N10687)? mem[81] : 
                  (N10689)? mem[83] : 
                  (N10691)? mem[85] : 
                  (N10693)? mem[87] : 
                  (N10695)? mem[89] : 
                  (N10697)? mem[91] : 
                  (N10699)? mem[93] : 
                  (N10701)? mem[95] : 
                  (N10703)? mem[97] : 
                  (N10705)? mem[99] : 
                  (N10707)? mem[101] : 
                  (N10709)? mem[103] : 
                  (N10711)? mem[105] : 
                  (N10713)? mem[107] : 
                  (N10715)? mem[109] : 
                  (N10717)? mem[111] : 
                  (N10719)? mem[113] : 
                  (N10721)? mem[115] : 
                  (N10723)? mem[117] : 
                  (N10725)? mem[119] : 
                  (N10727)? mem[121] : 
                  (N10729)? mem[123] : 
                  (N10731)? mem[125] : 
                  (N10733)? mem[127] : 
                  (N10735)? mem[129] : 
                  (N10737)? mem[131] : 
                  (N10739)? mem[133] : 
                  (N10741)? mem[135] : 
                  (N10743)? mem[137] : 
                  (N10745)? mem[139] : 
                  (N10747)? mem[141] : 
                  (N10749)? mem[143] : 
                  (N10751)? mem[145] : 
                  (N10753)? mem[147] : 
                  (N10755)? mem[149] : 
                  (N10757)? mem[151] : 
                  (N10759)? mem[153] : 
                  (N10761)? mem[155] : 
                  (N10763)? mem[157] : 
                  (N10765)? mem[159] : 
                  (N10767)? mem[161] : 
                  (N10769)? mem[163] : 
                  (N10771)? mem[165] : 
                  (N10773)? mem[167] : 
                  (N10775)? mem[169] : 
                  (N10777)? mem[171] : 
                  (N10779)? mem[173] : 
                  (N10781)? mem[175] : 
                  (N10783)? mem[177] : 
                  (N10785)? mem[179] : 
                  (N10787)? mem[181] : 
                  (N10789)? mem[183] : 
                  (N10791)? mem[185] : 
                  (N10793)? mem[187] : 
                  (N10795)? mem[189] : 
                  (N10797)? mem[191] : 
                  (N10799)? mem[193] : 
                  (N10801)? mem[195] : 
                  (N10803)? mem[197] : 
                  (N10805)? mem[199] : 
                  (N10807)? mem[201] : 
                  (N10809)? mem[203] : 
                  (N10811)? mem[205] : 
                  (N10813)? mem[207] : 
                  (N10815)? mem[209] : 
                  (N10817)? mem[211] : 
                  (N10819)? mem[213] : 
                  (N10821)? mem[215] : 
                  (N10823)? mem[217] : 
                  (N10825)? mem[219] : 
                  (N10827)? mem[221] : 
                  (N10829)? mem[223] : 
                  (N10831)? mem[225] : 
                  (N10833)? mem[227] : 
                  (N10835)? mem[229] : 
                  (N10837)? mem[231] : 
                  (N10839)? mem[233] : 
                  (N10841)? mem[235] : 
                  (N10843)? mem[237] : 
                  (N10845)? mem[239] : 
                  (N10847)? mem[241] : 
                  (N10849)? mem[243] : 
                  (N10851)? mem[245] : 
                  (N10853)? mem[247] : 
                  (N10855)? mem[249] : 
                  (N10857)? mem[251] : 
                  (N10859)? mem[253] : 
                  (N10861)? mem[255] : 
                  (N10863)? mem[257] : 
                  (N10865)? mem[259] : 
                  (N10867)? mem[261] : 
                  (N10869)? mem[263] : 
                  (N10871)? mem[265] : 
                  (N10873)? mem[267] : 
                  (N10875)? mem[269] : 
                  (N10877)? mem[271] : 
                  (N10879)? mem[273] : 
                  (N10881)? mem[275] : 
                  (N10883)? mem[277] : 
                  (N10885)? mem[279] : 
                  (N10887)? mem[281] : 
                  (N10889)? mem[283] : 
                  (N10891)? mem[285] : 
                  (N10893)? mem[287] : 
                  (N10895)? mem[289] : 
                  (N10897)? mem[291] : 
                  (N10899)? mem[293] : 
                  (N10901)? mem[295] : 
                  (N10903)? mem[297] : 
                  (N10905)? mem[299] : 
                  (N10907)? mem[301] : 
                  (N10909)? mem[303] : 
                  (N10911)? mem[305] : 
                  (N10913)? mem[307] : 
                  (N10915)? mem[309] : 
                  (N10917)? mem[311] : 
                  (N10919)? mem[313] : 
                  (N10921)? mem[315] : 
                  (N10923)? mem[317] : 
                  (N10925)? mem[319] : 
                  (N10927)? mem[321] : 
                  (N10929)? mem[323] : 
                  (N10931)? mem[325] : 
                  (N10933)? mem[327] : 
                  (N10935)? mem[329] : 
                  (N10937)? mem[331] : 
                  (N10939)? mem[333] : 
                  (N10941)? mem[335] : 
                  (N10943)? mem[337] : 
                  (N10945)? mem[339] : 
                  (N10947)? mem[341] : 
                  (N10949)? mem[343] : 
                  (N10951)? mem[345] : 
                  (N10953)? mem[347] : 
                  (N10955)? mem[349] : 
                  (N10957)? mem[351] : 
                  (N10959)? mem[353] : 
                  (N10961)? mem[355] : 
                  (N10963)? mem[357] : 
                  (N10965)? mem[359] : 
                  (N10967)? mem[361] : 
                  (N10969)? mem[363] : 
                  (N10971)? mem[365] : 
                  (N10973)? mem[367] : 
                  (N10975)? mem[369] : 
                  (N10977)? mem[371] : 
                  (N10979)? mem[373] : 
                  (N10981)? mem[375] : 
                  (N10983)? mem[377] : 
                  (N10985)? mem[379] : 
                  (N10987)? mem[381] : 
                  (N10989)? mem[383] : 
                  (N10991)? mem[385] : 
                  (N10993)? mem[387] : 
                  (N10995)? mem[389] : 
                  (N10997)? mem[391] : 
                  (N10999)? mem[393] : 
                  (N11001)? mem[395] : 
                  (N11003)? mem[397] : 
                  (N11005)? mem[399] : 
                  (N11007)? mem[401] : 
                  (N11009)? mem[403] : 
                  (N11011)? mem[405] : 
                  (N11013)? mem[407] : 
                  (N11015)? mem[409] : 
                  (N11017)? mem[411] : 
                  (N11019)? mem[413] : 
                  (N11021)? mem[415] : 
                  (N11023)? mem[417] : 
                  (N11025)? mem[419] : 
                  (N11027)? mem[421] : 
                  (N11029)? mem[423] : 
                  (N11031)? mem[425] : 
                  (N11033)? mem[427] : 
                  (N11035)? mem[429] : 
                  (N11037)? mem[431] : 
                  (N11039)? mem[433] : 
                  (N11041)? mem[435] : 
                  (N11043)? mem[437] : 
                  (N11045)? mem[439] : 
                  (N11047)? mem[441] : 
                  (N11049)? mem[443] : 
                  (N11051)? mem[445] : 
                  (N11053)? mem[447] : 
                  (N11055)? mem[449] : 
                  (N11056)? mem[451] : 
                  (N11057)? mem[453] : 
                  (N11058)? mem[455] : 
                  (N11059)? mem[457] : 
                  (N11060)? mem[459] : 
                  (N11061)? mem[461] : 
                  (N11062)? mem[463] : 
                  (N11063)? mem[465] : 
                  (N11064)? mem[467] : 
                  (N11065)? mem[469] : 
                  (N11066)? mem[471] : 
                  (N11067)? mem[473] : 
                  (N11068)? mem[475] : 
                  (N11069)? mem[477] : 
                  (N11070)? mem[479] : 
                  (N11071)? mem[481] : 
                  (N11072)? mem[483] : 
                  (N11073)? mem[485] : 
                  (N11074)? mem[487] : 
                  (N11075)? mem[489] : 
                  (N11076)? mem[491] : 
                  (N11077)? mem[493] : 
                  (N11078)? mem[495] : 
                  (N11079)? mem[497] : 
                  (N11080)? mem[499] : 
                  (N11081)? mem[501] : 
                  (N11082)? mem[503] : 
                  (N11083)? mem[505] : 
                  (N11084)? mem[507] : 
                  (N11085)? mem[509] : 
                  (N11086)? mem[511] : 
                  (N10608)? mem[513] : 
                  (N10610)? mem[515] : 
                  (N10612)? mem[517] : 
                  (N10614)? mem[519] : 
                  (N10616)? mem[521] : 
                  (N10618)? mem[523] : 
                  (N10620)? mem[525] : 
                  (N10622)? mem[527] : 
                  (N10624)? mem[529] : 
                  (N10626)? mem[531] : 
                  (N10628)? mem[533] : 
                  (N10630)? mem[535] : 
                  (N10632)? mem[537] : 
                  (N10634)? mem[539] : 
                  (N10636)? mem[541] : 
                  (N10638)? mem[543] : 
                  (N10640)? mem[545] : 
                  (N10642)? mem[547] : 
                  (N10644)? mem[549] : 
                  (N10646)? mem[551] : 
                  (N10648)? mem[553] : 
                  (N10650)? mem[555] : 
                  (N10652)? mem[557] : 
                  (N10654)? mem[559] : 
                  (N10656)? mem[561] : 
                  (N10658)? mem[563] : 
                  (N10660)? mem[565] : 
                  (N10662)? mem[567] : 
                  (N10664)? mem[569] : 
                  (N10666)? mem[571] : 
                  (N10668)? mem[573] : 
                  (N10670)? mem[575] : 
                  (N10672)? mem[577] : 
                  (N10674)? mem[579] : 
                  (N10676)? mem[581] : 
                  (N10678)? mem[583] : 
                  (N10680)? mem[585] : 
                  (N10682)? mem[587] : 
                  (N10684)? mem[589] : 
                  (N10686)? mem[591] : 
                  (N10688)? mem[593] : 
                  (N10690)? mem[595] : 
                  (N10692)? mem[597] : 
                  (N10694)? mem[599] : 
                  (N10696)? mem[601] : 
                  (N10698)? mem[603] : 
                  (N10700)? mem[605] : 
                  (N10702)? mem[607] : 
                  (N10704)? mem[609] : 
                  (N10706)? mem[611] : 
                  (N10708)? mem[613] : 
                  (N10710)? mem[615] : 
                  (N10712)? mem[617] : 
                  (N10714)? mem[619] : 
                  (N10716)? mem[621] : 
                  (N10718)? mem[623] : 
                  (N10720)? mem[625] : 
                  (N10722)? mem[627] : 
                  (N10724)? mem[629] : 
                  (N10726)? mem[631] : 
                  (N10728)? mem[633] : 
                  (N10730)? mem[635] : 
                  (N10732)? mem[637] : 
                  (N10734)? mem[639] : 
                  (N10736)? mem[641] : 
                  (N10738)? mem[643] : 
                  (N10740)? mem[645] : 
                  (N10742)? mem[647] : 
                  (N10744)? mem[649] : 
                  (N10746)? mem[651] : 
                  (N10748)? mem[653] : 
                  (N10750)? mem[655] : 
                  (N10752)? mem[657] : 
                  (N10754)? mem[659] : 
                  (N10756)? mem[661] : 
                  (N10758)? mem[663] : 
                  (N10760)? mem[665] : 
                  (N10762)? mem[667] : 
                  (N10764)? mem[669] : 
                  (N10766)? mem[671] : 
                  (N10768)? mem[673] : 
                  (N10770)? mem[675] : 
                  (N10772)? mem[677] : 
                  (N10774)? mem[679] : 
                  (N10776)? mem[681] : 
                  (N10778)? mem[683] : 
                  (N10780)? mem[685] : 
                  (N10782)? mem[687] : 
                  (N10784)? mem[689] : 
                  (N10786)? mem[691] : 
                  (N10788)? mem[693] : 
                  (N10790)? mem[695] : 
                  (N10792)? mem[697] : 
                  (N10794)? mem[699] : 
                  (N10796)? mem[701] : 
                  (N10798)? mem[703] : 
                  (N10800)? mem[705] : 
                  (N10802)? mem[707] : 
                  (N10804)? mem[709] : 
                  (N10806)? mem[711] : 
                  (N10808)? mem[713] : 
                  (N10810)? mem[715] : 
                  (N10812)? mem[717] : 
                  (N10814)? mem[719] : 
                  (N10816)? mem[721] : 
                  (N10818)? mem[723] : 
                  (N10820)? mem[725] : 
                  (N10822)? mem[727] : 
                  (N10824)? mem[729] : 
                  (N10826)? mem[731] : 
                  (N10828)? mem[733] : 
                  (N10830)? mem[735] : 
                  (N10832)? mem[737] : 
                  (N10834)? mem[739] : 
                  (N10836)? mem[741] : 
                  (N10838)? mem[743] : 
                  (N10840)? mem[745] : 
                  (N10842)? mem[747] : 
                  (N10844)? mem[749] : 
                  (N10846)? mem[751] : 
                  (N10848)? mem[753] : 
                  (N10850)? mem[755] : 
                  (N10852)? mem[757] : 
                  (N10854)? mem[759] : 
                  (N10856)? mem[761] : 
                  (N10858)? mem[763] : 
                  (N10860)? mem[765] : 
                  (N10862)? mem[767] : 
                  (N10864)? mem[769] : 
                  (N10866)? mem[771] : 
                  (N10868)? mem[773] : 
                  (N10870)? mem[775] : 
                  (N10872)? mem[777] : 
                  (N10874)? mem[779] : 
                  (N10876)? mem[781] : 
                  (N10878)? mem[783] : 
                  (N10880)? mem[785] : 
                  (N10882)? mem[787] : 
                  (N10884)? mem[789] : 
                  (N10886)? mem[791] : 
                  (N10888)? mem[793] : 
                  (N10890)? mem[795] : 
                  (N10892)? mem[797] : 
                  (N10894)? mem[799] : 
                  (N10896)? mem[801] : 
                  (N10898)? mem[803] : 
                  (N10900)? mem[805] : 
                  (N10902)? mem[807] : 
                  (N10904)? mem[809] : 
                  (N10906)? mem[811] : 
                  (N10908)? mem[813] : 
                  (N10910)? mem[815] : 
                  (N10912)? mem[817] : 
                  (N10914)? mem[819] : 
                  (N10916)? mem[821] : 
                  (N10918)? mem[823] : 
                  (N10920)? mem[825] : 
                  (N10922)? mem[827] : 
                  (N10924)? mem[829] : 
                  (N10926)? mem[831] : 
                  (N10928)? mem[833] : 
                  (N10930)? mem[835] : 
                  (N10932)? mem[837] : 
                  (N10934)? mem[839] : 
                  (N10936)? mem[841] : 
                  (N10938)? mem[843] : 
                  (N10940)? mem[845] : 
                  (N10942)? mem[847] : 
                  (N10944)? mem[849] : 
                  (N10946)? mem[851] : 
                  (N10948)? mem[853] : 
                  (N10950)? mem[855] : 
                  (N10952)? mem[857] : 
                  (N10954)? mem[859] : 
                  (N10956)? mem[861] : 
                  (N10958)? mem[863] : 
                  (N10960)? mem[865] : 
                  (N10962)? mem[867] : 
                  (N10964)? mem[869] : 
                  (N10966)? mem[871] : 
                  (N10968)? mem[873] : 
                  (N10970)? mem[875] : 
                  (N10972)? mem[877] : 
                  (N10974)? mem[879] : 
                  (N10976)? mem[881] : 
                  (N10978)? mem[883] : 
                  (N10980)? mem[885] : 
                  (N10982)? mem[887] : 
                  (N10984)? mem[889] : 
                  (N10986)? mem[891] : 
                  (N10988)? mem[893] : 
                  (N10990)? mem[895] : 
                  (N10992)? mem[897] : 
                  (N10994)? mem[899] : 
                  (N10996)? mem[901] : 
                  (N10998)? mem[903] : 
                  (N11000)? mem[905] : 
                  (N11002)? mem[907] : 
                  (N11004)? mem[909] : 
                  (N11006)? mem[911] : 
                  (N11008)? mem[913] : 
                  (N11010)? mem[915] : 
                  (N11012)? mem[917] : 
                  (N11014)? mem[919] : 
                  (N11016)? mem[921] : 
                  (N11018)? mem[923] : 
                  (N11020)? mem[925] : 
                  (N11022)? mem[927] : 
                  (N11024)? mem[929] : 
                  (N11026)? mem[931] : 
                  (N11028)? mem[933] : 
                  (N11030)? mem[935] : 
                  (N11032)? mem[937] : 
                  (N11034)? mem[939] : 
                  (N11036)? mem[941] : 
                  (N11038)? mem[943] : 
                  (N11040)? mem[945] : 
                  (N11042)? mem[947] : 
                  (N11044)? mem[949] : 
                  (N11046)? mem[951] : 
                  (N11048)? mem[953] : 
                  (N11050)? mem[955] : 
                  (N11052)? mem[957] : 
                  (N11054)? mem[959] : 
                  (N12049)? mem[961] : 
                  (N12051)? mem[963] : 
                  (N12053)? mem[965] : 
                  (N12055)? mem[967] : 
                  (N12057)? mem[969] : 
                  (N12059)? mem[971] : 
                  (N12061)? mem[973] : 
                  (N12063)? mem[975] : 
                  (N12065)? mem[977] : 
                  (N12067)? mem[979] : 
                  (N12069)? mem[981] : 
                  (N12071)? mem[983] : 
                  (N12073)? mem[985] : 
                  (N12075)? mem[987] : 
                  (N12077)? mem[989] : 
                  (N12079)? mem[991] : 
                  (N12081)? mem[993] : 
                  (N12083)? mem[995] : 
                  (N12085)? mem[997] : 
                  (N12087)? mem[999] : 
                  (N12089)? mem[1001] : 
                  (N12091)? mem[1003] : 
                  (N12093)? mem[1005] : 
                  (N12095)? mem[1007] : 
                  (N12097)? mem[1009] : 
                  (N12099)? mem[1011] : 
                  (N12101)? mem[1013] : 
                  (N12103)? mem[1015] : 
                  (N12105)? mem[1017] : 
                  (N12107)? mem[1019] : 
                  (N12109)? mem[1021] : 
                  (N12111)? mem[1023] : 1'b0;
  assign N11088 = (N10607)? mem[0] : 
                  (N10609)? mem[2] : 
                  (N10611)? mem[4] : 
                  (N10613)? mem[6] : 
                  (N10615)? mem[8] : 
                  (N10617)? mem[10] : 
                  (N10619)? mem[12] : 
                  (N10621)? mem[14] : 
                  (N10623)? mem[16] : 
                  (N10625)? mem[18] : 
                  (N10627)? mem[20] : 
                  (N10629)? mem[22] : 
                  (N10631)? mem[24] : 
                  (N10633)? mem[26] : 
                  (N10635)? mem[28] : 
                  (N10637)? mem[30] : 
                  (N10639)? mem[32] : 
                  (N10641)? mem[34] : 
                  (N10643)? mem[36] : 
                  (N10645)? mem[38] : 
                  (N10647)? mem[40] : 
                  (N10649)? mem[42] : 
                  (N10651)? mem[44] : 
                  (N10653)? mem[46] : 
                  (N10655)? mem[48] : 
                  (N10657)? mem[50] : 
                  (N10659)? mem[52] : 
                  (N10661)? mem[54] : 
                  (N10663)? mem[56] : 
                  (N10665)? mem[58] : 
                  (N10667)? mem[60] : 
                  (N10669)? mem[62] : 
                  (N10671)? mem[64] : 
                  (N10673)? mem[66] : 
                  (N10675)? mem[68] : 
                  (N10677)? mem[70] : 
                  (N10679)? mem[72] : 
                  (N10681)? mem[74] : 
                  (N10683)? mem[76] : 
                  (N10685)? mem[78] : 
                  (N10687)? mem[80] : 
                  (N10689)? mem[82] : 
                  (N10691)? mem[84] : 
                  (N10693)? mem[86] : 
                  (N10695)? mem[88] : 
                  (N10697)? mem[90] : 
                  (N10699)? mem[92] : 
                  (N10701)? mem[94] : 
                  (N10703)? mem[96] : 
                  (N10705)? mem[98] : 
                  (N10707)? mem[100] : 
                  (N10709)? mem[102] : 
                  (N10711)? mem[104] : 
                  (N10713)? mem[106] : 
                  (N10715)? mem[108] : 
                  (N10717)? mem[110] : 
                  (N10719)? mem[112] : 
                  (N10721)? mem[114] : 
                  (N10723)? mem[116] : 
                  (N10725)? mem[118] : 
                  (N10727)? mem[120] : 
                  (N10729)? mem[122] : 
                  (N10731)? mem[124] : 
                  (N10733)? mem[126] : 
                  (N10735)? mem[128] : 
                  (N10737)? mem[130] : 
                  (N10739)? mem[132] : 
                  (N10741)? mem[134] : 
                  (N10743)? mem[136] : 
                  (N10745)? mem[138] : 
                  (N10747)? mem[140] : 
                  (N10749)? mem[142] : 
                  (N10751)? mem[144] : 
                  (N10753)? mem[146] : 
                  (N10755)? mem[148] : 
                  (N10757)? mem[150] : 
                  (N10759)? mem[152] : 
                  (N10761)? mem[154] : 
                  (N10763)? mem[156] : 
                  (N10765)? mem[158] : 
                  (N10767)? mem[160] : 
                  (N10769)? mem[162] : 
                  (N10771)? mem[164] : 
                  (N10773)? mem[166] : 
                  (N10775)? mem[168] : 
                  (N10777)? mem[170] : 
                  (N10779)? mem[172] : 
                  (N10781)? mem[174] : 
                  (N10783)? mem[176] : 
                  (N10785)? mem[178] : 
                  (N10787)? mem[180] : 
                  (N10789)? mem[182] : 
                  (N10791)? mem[184] : 
                  (N10793)? mem[186] : 
                  (N10795)? mem[188] : 
                  (N10797)? mem[190] : 
                  (N10799)? mem[192] : 
                  (N10801)? mem[194] : 
                  (N10803)? mem[196] : 
                  (N10805)? mem[198] : 
                  (N10807)? mem[200] : 
                  (N10809)? mem[202] : 
                  (N10811)? mem[204] : 
                  (N10813)? mem[206] : 
                  (N10815)? mem[208] : 
                  (N10817)? mem[210] : 
                  (N10819)? mem[212] : 
                  (N10821)? mem[214] : 
                  (N10823)? mem[216] : 
                  (N10825)? mem[218] : 
                  (N10827)? mem[220] : 
                  (N10829)? mem[222] : 
                  (N10831)? mem[224] : 
                  (N10833)? mem[226] : 
                  (N10835)? mem[228] : 
                  (N10837)? mem[230] : 
                  (N10839)? mem[232] : 
                  (N10841)? mem[234] : 
                  (N10843)? mem[236] : 
                  (N10845)? mem[238] : 
                  (N10847)? mem[240] : 
                  (N10849)? mem[242] : 
                  (N10851)? mem[244] : 
                  (N10853)? mem[246] : 
                  (N10855)? mem[248] : 
                  (N10857)? mem[250] : 
                  (N10859)? mem[252] : 
                  (N10861)? mem[254] : 
                  (N10863)? mem[256] : 
                  (N10865)? mem[258] : 
                  (N10867)? mem[260] : 
                  (N10869)? mem[262] : 
                  (N10871)? mem[264] : 
                  (N10873)? mem[266] : 
                  (N10875)? mem[268] : 
                  (N10877)? mem[270] : 
                  (N10879)? mem[272] : 
                  (N10881)? mem[274] : 
                  (N10883)? mem[276] : 
                  (N10885)? mem[278] : 
                  (N10887)? mem[280] : 
                  (N10889)? mem[282] : 
                  (N10891)? mem[284] : 
                  (N10893)? mem[286] : 
                  (N10895)? mem[288] : 
                  (N10897)? mem[290] : 
                  (N10899)? mem[292] : 
                  (N10901)? mem[294] : 
                  (N10903)? mem[296] : 
                  (N10905)? mem[298] : 
                  (N10907)? mem[300] : 
                  (N10909)? mem[302] : 
                  (N10911)? mem[304] : 
                  (N10913)? mem[306] : 
                  (N10915)? mem[308] : 
                  (N10917)? mem[310] : 
                  (N10919)? mem[312] : 
                  (N10921)? mem[314] : 
                  (N10923)? mem[316] : 
                  (N10925)? mem[318] : 
                  (N10927)? mem[320] : 
                  (N10929)? mem[322] : 
                  (N10931)? mem[324] : 
                  (N10933)? mem[326] : 
                  (N10935)? mem[328] : 
                  (N10937)? mem[330] : 
                  (N10939)? mem[332] : 
                  (N10941)? mem[334] : 
                  (N10943)? mem[336] : 
                  (N10945)? mem[338] : 
                  (N10947)? mem[340] : 
                  (N10949)? mem[342] : 
                  (N10951)? mem[344] : 
                  (N10953)? mem[346] : 
                  (N10955)? mem[348] : 
                  (N10957)? mem[350] : 
                  (N10959)? mem[352] : 
                  (N10961)? mem[354] : 
                  (N10963)? mem[356] : 
                  (N10965)? mem[358] : 
                  (N10967)? mem[360] : 
                  (N10969)? mem[362] : 
                  (N10971)? mem[364] : 
                  (N10973)? mem[366] : 
                  (N10975)? mem[368] : 
                  (N10977)? mem[370] : 
                  (N10979)? mem[372] : 
                  (N10981)? mem[374] : 
                  (N10983)? mem[376] : 
                  (N10985)? mem[378] : 
                  (N10987)? mem[380] : 
                  (N10989)? mem[382] : 
                  (N10991)? mem[384] : 
                  (N10993)? mem[386] : 
                  (N10995)? mem[388] : 
                  (N10997)? mem[390] : 
                  (N10999)? mem[392] : 
                  (N11001)? mem[394] : 
                  (N11003)? mem[396] : 
                  (N11005)? mem[398] : 
                  (N11007)? mem[400] : 
                  (N11009)? mem[402] : 
                  (N11011)? mem[404] : 
                  (N11013)? mem[406] : 
                  (N11015)? mem[408] : 
                  (N11017)? mem[410] : 
                  (N11019)? mem[412] : 
                  (N11021)? mem[414] : 
                  (N11023)? mem[416] : 
                  (N11025)? mem[418] : 
                  (N11027)? mem[420] : 
                  (N11029)? mem[422] : 
                  (N11031)? mem[424] : 
                  (N11033)? mem[426] : 
                  (N11035)? mem[428] : 
                  (N11037)? mem[430] : 
                  (N11039)? mem[432] : 
                  (N11041)? mem[434] : 
                  (N11043)? mem[436] : 
                  (N11045)? mem[438] : 
                  (N11047)? mem[440] : 
                  (N11049)? mem[442] : 
                  (N11051)? mem[444] : 
                  (N11053)? mem[446] : 
                  (N11055)? mem[448] : 
                  (N11056)? mem[450] : 
                  (N11057)? mem[452] : 
                  (N11058)? mem[454] : 
                  (N11059)? mem[456] : 
                  (N11060)? mem[458] : 
                  (N11061)? mem[460] : 
                  (N11062)? mem[462] : 
                  (N11063)? mem[464] : 
                  (N11064)? mem[466] : 
                  (N11065)? mem[468] : 
                  (N11066)? mem[470] : 
                  (N11067)? mem[472] : 
                  (N11068)? mem[474] : 
                  (N11069)? mem[476] : 
                  (N11070)? mem[478] : 
                  (N11071)? mem[480] : 
                  (N11072)? mem[482] : 
                  (N11073)? mem[484] : 
                  (N11074)? mem[486] : 
                  (N11075)? mem[488] : 
                  (N11076)? mem[490] : 
                  (N11077)? mem[492] : 
                  (N11078)? mem[494] : 
                  (N11079)? mem[496] : 
                  (N11080)? mem[498] : 
                  (N11081)? mem[500] : 
                  (N11082)? mem[502] : 
                  (N11083)? mem[504] : 
                  (N11084)? mem[506] : 
                  (N11085)? mem[508] : 
                  (N11086)? mem[510] : 
                  (N10608)? mem[512] : 
                  (N10610)? mem[514] : 
                  (N10612)? mem[516] : 
                  (N10614)? mem[518] : 
                  (N10616)? mem[520] : 
                  (N10618)? mem[522] : 
                  (N10620)? mem[524] : 
                  (N10622)? mem[526] : 
                  (N10624)? mem[528] : 
                  (N10626)? mem[530] : 
                  (N10628)? mem[532] : 
                  (N10630)? mem[534] : 
                  (N10632)? mem[536] : 
                  (N10634)? mem[538] : 
                  (N10636)? mem[540] : 
                  (N10638)? mem[542] : 
                  (N10640)? mem[544] : 
                  (N10642)? mem[546] : 
                  (N10644)? mem[548] : 
                  (N10646)? mem[550] : 
                  (N10648)? mem[552] : 
                  (N10650)? mem[554] : 
                  (N10652)? mem[556] : 
                  (N10654)? mem[558] : 
                  (N10656)? mem[560] : 
                  (N10658)? mem[562] : 
                  (N10660)? mem[564] : 
                  (N10662)? mem[566] : 
                  (N10664)? mem[568] : 
                  (N10666)? mem[570] : 
                  (N10668)? mem[572] : 
                  (N10670)? mem[574] : 
                  (N10672)? mem[576] : 
                  (N10674)? mem[578] : 
                  (N10676)? mem[580] : 
                  (N10678)? mem[582] : 
                  (N10680)? mem[584] : 
                  (N10682)? mem[586] : 
                  (N10684)? mem[588] : 
                  (N10686)? mem[590] : 
                  (N10688)? mem[592] : 
                  (N10690)? mem[594] : 
                  (N10692)? mem[596] : 
                  (N10694)? mem[598] : 
                  (N10696)? mem[600] : 
                  (N10698)? mem[602] : 
                  (N10700)? mem[604] : 
                  (N10702)? mem[606] : 
                  (N10704)? mem[608] : 
                  (N10706)? mem[610] : 
                  (N10708)? mem[612] : 
                  (N10710)? mem[614] : 
                  (N10712)? mem[616] : 
                  (N10714)? mem[618] : 
                  (N10716)? mem[620] : 
                  (N10718)? mem[622] : 
                  (N10720)? mem[624] : 
                  (N10722)? mem[626] : 
                  (N10724)? mem[628] : 
                  (N10726)? mem[630] : 
                  (N10728)? mem[632] : 
                  (N10730)? mem[634] : 
                  (N10732)? mem[636] : 
                  (N10734)? mem[638] : 
                  (N10736)? mem[640] : 
                  (N10738)? mem[642] : 
                  (N10740)? mem[644] : 
                  (N10742)? mem[646] : 
                  (N10744)? mem[648] : 
                  (N10746)? mem[650] : 
                  (N10748)? mem[652] : 
                  (N10750)? mem[654] : 
                  (N10752)? mem[656] : 
                  (N10754)? mem[658] : 
                  (N10756)? mem[660] : 
                  (N10758)? mem[662] : 
                  (N10760)? mem[664] : 
                  (N10762)? mem[666] : 
                  (N10764)? mem[668] : 
                  (N10766)? mem[670] : 
                  (N10768)? mem[672] : 
                  (N10770)? mem[674] : 
                  (N10772)? mem[676] : 
                  (N10774)? mem[678] : 
                  (N10776)? mem[680] : 
                  (N10778)? mem[682] : 
                  (N10780)? mem[684] : 
                  (N10782)? mem[686] : 
                  (N10784)? mem[688] : 
                  (N10786)? mem[690] : 
                  (N10788)? mem[692] : 
                  (N10790)? mem[694] : 
                  (N10792)? mem[696] : 
                  (N10794)? mem[698] : 
                  (N10796)? mem[700] : 
                  (N10798)? mem[702] : 
                  (N10800)? mem[704] : 
                  (N10802)? mem[706] : 
                  (N10804)? mem[708] : 
                  (N10806)? mem[710] : 
                  (N10808)? mem[712] : 
                  (N10810)? mem[714] : 
                  (N10812)? mem[716] : 
                  (N10814)? mem[718] : 
                  (N10816)? mem[720] : 
                  (N10818)? mem[722] : 
                  (N10820)? mem[724] : 
                  (N10822)? mem[726] : 
                  (N10824)? mem[728] : 
                  (N10826)? mem[730] : 
                  (N10828)? mem[732] : 
                  (N10830)? mem[734] : 
                  (N10832)? mem[736] : 
                  (N10834)? mem[738] : 
                  (N10836)? mem[740] : 
                  (N10838)? mem[742] : 
                  (N10840)? mem[744] : 
                  (N10842)? mem[746] : 
                  (N10844)? mem[748] : 
                  (N10846)? mem[750] : 
                  (N10848)? mem[752] : 
                  (N10850)? mem[754] : 
                  (N10852)? mem[756] : 
                  (N10854)? mem[758] : 
                  (N10856)? mem[760] : 
                  (N10858)? mem[762] : 
                  (N10860)? mem[764] : 
                  (N10862)? mem[766] : 
                  (N10864)? mem[768] : 
                  (N10866)? mem[770] : 
                  (N10868)? mem[772] : 
                  (N10870)? mem[774] : 
                  (N10872)? mem[776] : 
                  (N10874)? mem[778] : 
                  (N10876)? mem[780] : 
                  (N10878)? mem[782] : 
                  (N10880)? mem[784] : 
                  (N10882)? mem[786] : 
                  (N10884)? mem[788] : 
                  (N10886)? mem[790] : 
                  (N10888)? mem[792] : 
                  (N10890)? mem[794] : 
                  (N10892)? mem[796] : 
                  (N10894)? mem[798] : 
                  (N10896)? mem[800] : 
                  (N10898)? mem[802] : 
                  (N10900)? mem[804] : 
                  (N10902)? mem[806] : 
                  (N10904)? mem[808] : 
                  (N10906)? mem[810] : 
                  (N10908)? mem[812] : 
                  (N10910)? mem[814] : 
                  (N10912)? mem[816] : 
                  (N10914)? mem[818] : 
                  (N10916)? mem[820] : 
                  (N10918)? mem[822] : 
                  (N10920)? mem[824] : 
                  (N10922)? mem[826] : 
                  (N10924)? mem[828] : 
                  (N10926)? mem[830] : 
                  (N10928)? mem[832] : 
                  (N10930)? mem[834] : 
                  (N10932)? mem[836] : 
                  (N10934)? mem[838] : 
                  (N10936)? mem[840] : 
                  (N10938)? mem[842] : 
                  (N10940)? mem[844] : 
                  (N10942)? mem[846] : 
                  (N10944)? mem[848] : 
                  (N10946)? mem[850] : 
                  (N10948)? mem[852] : 
                  (N10950)? mem[854] : 
                  (N10952)? mem[856] : 
                  (N10954)? mem[858] : 
                  (N10956)? mem[860] : 
                  (N10958)? mem[862] : 
                  (N10960)? mem[864] : 
                  (N10962)? mem[866] : 
                  (N10964)? mem[868] : 
                  (N10966)? mem[870] : 
                  (N10968)? mem[872] : 
                  (N10970)? mem[874] : 
                  (N10972)? mem[876] : 
                  (N10974)? mem[878] : 
                  (N10976)? mem[880] : 
                  (N10978)? mem[882] : 
                  (N10980)? mem[884] : 
                  (N10982)? mem[886] : 
                  (N10984)? mem[888] : 
                  (N10986)? mem[890] : 
                  (N10988)? mem[892] : 
                  (N10990)? mem[894] : 
                  (N10992)? mem[896] : 
                  (N10994)? mem[898] : 
                  (N10996)? mem[900] : 
                  (N10998)? mem[902] : 
                  (N11000)? mem[904] : 
                  (N11002)? mem[906] : 
                  (N11004)? mem[908] : 
                  (N11006)? mem[910] : 
                  (N11008)? mem[912] : 
                  (N11010)? mem[914] : 
                  (N11012)? mem[916] : 
                  (N11014)? mem[918] : 
                  (N11016)? mem[920] : 
                  (N11018)? mem[922] : 
                  (N11020)? mem[924] : 
                  (N11022)? mem[926] : 
                  (N11024)? mem[928] : 
                  (N11026)? mem[930] : 
                  (N11028)? mem[932] : 
                  (N11030)? mem[934] : 
                  (N11032)? mem[936] : 
                  (N11034)? mem[938] : 
                  (N11036)? mem[940] : 
                  (N11038)? mem[942] : 
                  (N11040)? mem[944] : 
                  (N11042)? mem[946] : 
                  (N11044)? mem[948] : 
                  (N11046)? mem[950] : 
                  (N11048)? mem[952] : 
                  (N11050)? mem[954] : 
                  (N11052)? mem[956] : 
                  (N11054)? mem[958] : 
                  (N12049)? mem[960] : 
                  (N12051)? mem[962] : 
                  (N12053)? mem[964] : 
                  (N12055)? mem[966] : 
                  (N12057)? mem[968] : 
                  (N12059)? mem[970] : 
                  (N12061)? mem[972] : 
                  (N12063)? mem[974] : 
                  (N12065)? mem[976] : 
                  (N12067)? mem[978] : 
                  (N12069)? mem[980] : 
                  (N12071)? mem[982] : 
                  (N12073)? mem[984] : 
                  (N12075)? mem[986] : 
                  (N12077)? mem[988] : 
                  (N12079)? mem[990] : 
                  (N12081)? mem[992] : 
                  (N12083)? mem[994] : 
                  (N12085)? mem[996] : 
                  (N12087)? mem[998] : 
                  (N12089)? mem[1000] : 
                  (N12091)? mem[1002] : 
                  (N12093)? mem[1004] : 
                  (N12095)? mem[1006] : 
                  (N12097)? mem[1008] : 
                  (N12099)? mem[1010] : 
                  (N12101)? mem[1012] : 
                  (N12103)? mem[1014] : 
                  (N12105)? mem[1016] : 
                  (N12107)? mem[1018] : 
                  (N12109)? mem[1020] : 
                  (N12111)? mem[1022] : 1'b0;
  assign N12112 = (N11600)? mem[1] : 
                  (N11602)? mem[3] : 
                  (N11604)? mem[5] : 
                  (N11606)? mem[7] : 
                  (N11608)? mem[9] : 
                  (N11610)? mem[11] : 
                  (N11612)? mem[13] : 
                  (N11614)? mem[15] : 
                  (N11616)? mem[17] : 
                  (N11618)? mem[19] : 
                  (N11620)? mem[21] : 
                  (N11622)? mem[23] : 
                  (N11624)? mem[25] : 
                  (N11626)? mem[27] : 
                  (N11628)? mem[29] : 
                  (N11630)? mem[31] : 
                  (N11632)? mem[33] : 
                  (N11634)? mem[35] : 
                  (N11636)? mem[37] : 
                  (N11638)? mem[39] : 
                  (N11640)? mem[41] : 
                  (N11642)? mem[43] : 
                  (N11644)? mem[45] : 
                  (N11646)? mem[47] : 
                  (N11648)? mem[49] : 
                  (N11650)? mem[51] : 
                  (N11652)? mem[53] : 
                  (N11654)? mem[55] : 
                  (N11656)? mem[57] : 
                  (N11658)? mem[59] : 
                  (N11660)? mem[61] : 
                  (N11662)? mem[63] : 
                  (N11664)? mem[65] : 
                  (N11666)? mem[67] : 
                  (N11668)? mem[69] : 
                  (N11670)? mem[71] : 
                  (N11672)? mem[73] : 
                  (N11674)? mem[75] : 
                  (N11676)? mem[77] : 
                  (N11678)? mem[79] : 
                  (N11680)? mem[81] : 
                  (N11682)? mem[83] : 
                  (N11684)? mem[85] : 
                  (N11686)? mem[87] : 
                  (N11688)? mem[89] : 
                  (N11690)? mem[91] : 
                  (N11692)? mem[93] : 
                  (N11694)? mem[95] : 
                  (N11696)? mem[97] : 
                  (N11698)? mem[99] : 
                  (N11700)? mem[101] : 
                  (N11702)? mem[103] : 
                  (N11704)? mem[105] : 
                  (N11706)? mem[107] : 
                  (N11708)? mem[109] : 
                  (N11710)? mem[111] : 
                  (N11712)? mem[113] : 
                  (N11714)? mem[115] : 
                  (N11716)? mem[117] : 
                  (N11718)? mem[119] : 
                  (N11720)? mem[121] : 
                  (N11722)? mem[123] : 
                  (N11724)? mem[125] : 
                  (N11726)? mem[127] : 
                  (N11728)? mem[129] : 
                  (N11730)? mem[131] : 
                  (N11732)? mem[133] : 
                  (N11734)? mem[135] : 
                  (N11736)? mem[137] : 
                  (N11738)? mem[139] : 
                  (N11740)? mem[141] : 
                  (N11742)? mem[143] : 
                  (N11744)? mem[145] : 
                  (N11746)? mem[147] : 
                  (N11748)? mem[149] : 
                  (N11750)? mem[151] : 
                  (N11752)? mem[153] : 
                  (N11754)? mem[155] : 
                  (N11756)? mem[157] : 
                  (N11758)? mem[159] : 
                  (N11760)? mem[161] : 
                  (N11762)? mem[163] : 
                  (N11764)? mem[165] : 
                  (N11766)? mem[167] : 
                  (N11768)? mem[169] : 
                  (N11770)? mem[171] : 
                  (N11772)? mem[173] : 
                  (N11774)? mem[175] : 
                  (N11776)? mem[177] : 
                  (N11778)? mem[179] : 
                  (N11780)? mem[181] : 
                  (N11782)? mem[183] : 
                  (N11784)? mem[185] : 
                  (N11786)? mem[187] : 
                  (N11788)? mem[189] : 
                  (N11790)? mem[191] : 
                  (N11792)? mem[193] : 
                  (N11794)? mem[195] : 
                  (N11796)? mem[197] : 
                  (N11798)? mem[199] : 
                  (N11800)? mem[201] : 
                  (N11802)? mem[203] : 
                  (N11804)? mem[205] : 
                  (N11806)? mem[207] : 
                  (N11808)? mem[209] : 
                  (N11810)? mem[211] : 
                  (N11812)? mem[213] : 
                  (N11814)? mem[215] : 
                  (N11816)? mem[217] : 
                  (N11818)? mem[219] : 
                  (N11820)? mem[221] : 
                  (N11822)? mem[223] : 
                  (N11824)? mem[225] : 
                  (N11826)? mem[227] : 
                  (N11828)? mem[229] : 
                  (N11830)? mem[231] : 
                  (N11832)? mem[233] : 
                  (N11834)? mem[235] : 
                  (N11836)? mem[237] : 
                  (N11838)? mem[239] : 
                  (N11840)? mem[241] : 
                  (N11842)? mem[243] : 
                  (N11844)? mem[245] : 
                  (N11846)? mem[247] : 
                  (N11848)? mem[249] : 
                  (N11850)? mem[251] : 
                  (N11852)? mem[253] : 
                  (N11854)? mem[255] : 
                  (N11856)? mem[257] : 
                  (N11858)? mem[259] : 
                  (N11860)? mem[261] : 
                  (N11862)? mem[263] : 
                  (N11864)? mem[265] : 
                  (N11866)? mem[267] : 
                  (N11868)? mem[269] : 
                  (N11870)? mem[271] : 
                  (N11872)? mem[273] : 
                  (N11874)? mem[275] : 
                  (N11876)? mem[277] : 
                  (N11878)? mem[279] : 
                  (N11880)? mem[281] : 
                  (N11882)? mem[283] : 
                  (N11884)? mem[285] : 
                  (N11886)? mem[287] : 
                  (N11888)? mem[289] : 
                  (N11890)? mem[291] : 
                  (N11892)? mem[293] : 
                  (N11894)? mem[295] : 
                  (N11896)? mem[297] : 
                  (N11898)? mem[299] : 
                  (N11900)? mem[301] : 
                  (N11902)? mem[303] : 
                  (N11904)? mem[305] : 
                  (N11906)? mem[307] : 
                  (N11908)? mem[309] : 
                  (N11910)? mem[311] : 
                  (N11912)? mem[313] : 
                  (N11914)? mem[315] : 
                  (N11916)? mem[317] : 
                  (N11918)? mem[319] : 
                  (N11920)? mem[321] : 
                  (N11922)? mem[323] : 
                  (N11924)? mem[325] : 
                  (N11926)? mem[327] : 
                  (N11928)? mem[329] : 
                  (N11930)? mem[331] : 
                  (N11932)? mem[333] : 
                  (N11934)? mem[335] : 
                  (N11936)? mem[337] : 
                  (N11938)? mem[339] : 
                  (N11940)? mem[341] : 
                  (N11942)? mem[343] : 
                  (N11944)? mem[345] : 
                  (N11946)? mem[347] : 
                  (N11948)? mem[349] : 
                  (N11950)? mem[351] : 
                  (N11952)? mem[353] : 
                  (N11954)? mem[355] : 
                  (N11956)? mem[357] : 
                  (N11958)? mem[359] : 
                  (N11960)? mem[361] : 
                  (N11962)? mem[363] : 
                  (N11964)? mem[365] : 
                  (N11966)? mem[367] : 
                  (N11968)? mem[369] : 
                  (N11970)? mem[371] : 
                  (N11972)? mem[373] : 
                  (N11974)? mem[375] : 
                  (N11976)? mem[377] : 
                  (N11978)? mem[379] : 
                  (N11980)? mem[381] : 
                  (N11982)? mem[383] : 
                  (N11984)? mem[385] : 
                  (N11986)? mem[387] : 
                  (N11988)? mem[389] : 
                  (N11990)? mem[391] : 
                  (N11992)? mem[393] : 
                  (N11994)? mem[395] : 
                  (N11996)? mem[397] : 
                  (N11998)? mem[399] : 
                  (N12000)? mem[401] : 
                  (N12002)? mem[403] : 
                  (N12004)? mem[405] : 
                  (N12006)? mem[407] : 
                  (N12008)? mem[409] : 
                  (N12010)? mem[411] : 
                  (N12012)? mem[413] : 
                  (N12014)? mem[415] : 
                  (N12016)? mem[417] : 
                  (N12018)? mem[419] : 
                  (N12020)? mem[421] : 
                  (N12022)? mem[423] : 
                  (N12024)? mem[425] : 
                  (N12026)? mem[427] : 
                  (N12028)? mem[429] : 
                  (N12030)? mem[431] : 
                  (N12032)? mem[433] : 
                  (N12034)? mem[435] : 
                  (N12036)? mem[437] : 
                  (N12038)? mem[439] : 
                  (N12040)? mem[441] : 
                  (N12042)? mem[443] : 
                  (N12044)? mem[445] : 
                  (N12046)? mem[447] : 
                  (N12048)? mem[449] : 
                  (N12050)? mem[451] : 
                  (N12052)? mem[453] : 
                  (N12054)? mem[455] : 
                  (N12056)? mem[457] : 
                  (N12058)? mem[459] : 
                  (N12060)? mem[461] : 
                  (N12062)? mem[463] : 
                  (N12064)? mem[465] : 
                  (N12066)? mem[467] : 
                  (N12068)? mem[469] : 
                  (N12070)? mem[471] : 
                  (N12072)? mem[473] : 
                  (N12074)? mem[475] : 
                  (N12076)? mem[477] : 
                  (N12078)? mem[479] : 
                  (N12080)? mem[481] : 
                  (N12082)? mem[483] : 
                  (N12084)? mem[485] : 
                  (N12086)? mem[487] : 
                  (N12088)? mem[489] : 
                  (N12090)? mem[491] : 
                  (N12092)? mem[493] : 
                  (N12094)? mem[495] : 
                  (N12096)? mem[497] : 
                  (N12098)? mem[499] : 
                  (N12100)? mem[501] : 
                  (N12102)? mem[503] : 
                  (N12104)? mem[505] : 
                  (N12106)? mem[507] : 
                  (N12108)? mem[509] : 
                  (N12110)? mem[511] : 
                  (N11601)? mem[513] : 
                  (N11603)? mem[515] : 
                  (N11605)? mem[517] : 
                  (N11607)? mem[519] : 
                  (N11609)? mem[521] : 
                  (N11611)? mem[523] : 
                  (N11613)? mem[525] : 
                  (N11615)? mem[527] : 
                  (N11617)? mem[529] : 
                  (N11619)? mem[531] : 
                  (N11621)? mem[533] : 
                  (N11623)? mem[535] : 
                  (N11625)? mem[537] : 
                  (N11627)? mem[539] : 
                  (N11629)? mem[541] : 
                  (N11631)? mem[543] : 
                  (N11633)? mem[545] : 
                  (N11635)? mem[547] : 
                  (N11637)? mem[549] : 
                  (N11639)? mem[551] : 
                  (N11641)? mem[553] : 
                  (N11643)? mem[555] : 
                  (N11645)? mem[557] : 
                  (N11647)? mem[559] : 
                  (N11649)? mem[561] : 
                  (N11651)? mem[563] : 
                  (N11653)? mem[565] : 
                  (N11655)? mem[567] : 
                  (N11657)? mem[569] : 
                  (N11659)? mem[571] : 
                  (N11661)? mem[573] : 
                  (N11663)? mem[575] : 
                  (N11665)? mem[577] : 
                  (N11667)? mem[579] : 
                  (N11669)? mem[581] : 
                  (N11671)? mem[583] : 
                  (N11673)? mem[585] : 
                  (N11675)? mem[587] : 
                  (N11677)? mem[589] : 
                  (N11679)? mem[591] : 
                  (N11681)? mem[593] : 
                  (N11683)? mem[595] : 
                  (N11685)? mem[597] : 
                  (N11687)? mem[599] : 
                  (N11689)? mem[601] : 
                  (N11691)? mem[603] : 
                  (N11693)? mem[605] : 
                  (N11695)? mem[607] : 
                  (N11697)? mem[609] : 
                  (N11699)? mem[611] : 
                  (N11701)? mem[613] : 
                  (N11703)? mem[615] : 
                  (N11705)? mem[617] : 
                  (N11707)? mem[619] : 
                  (N11709)? mem[621] : 
                  (N11711)? mem[623] : 
                  (N11713)? mem[625] : 
                  (N11715)? mem[627] : 
                  (N11717)? mem[629] : 
                  (N11719)? mem[631] : 
                  (N11721)? mem[633] : 
                  (N11723)? mem[635] : 
                  (N11725)? mem[637] : 
                  (N11727)? mem[639] : 
                  (N11729)? mem[641] : 
                  (N11731)? mem[643] : 
                  (N11733)? mem[645] : 
                  (N11735)? mem[647] : 
                  (N11737)? mem[649] : 
                  (N11739)? mem[651] : 
                  (N11741)? mem[653] : 
                  (N11743)? mem[655] : 
                  (N11745)? mem[657] : 
                  (N11747)? mem[659] : 
                  (N11749)? mem[661] : 
                  (N11751)? mem[663] : 
                  (N11753)? mem[665] : 
                  (N11755)? mem[667] : 
                  (N11757)? mem[669] : 
                  (N11759)? mem[671] : 
                  (N11761)? mem[673] : 
                  (N11763)? mem[675] : 
                  (N11765)? mem[677] : 
                  (N11767)? mem[679] : 
                  (N11769)? mem[681] : 
                  (N11771)? mem[683] : 
                  (N11773)? mem[685] : 
                  (N11775)? mem[687] : 
                  (N11777)? mem[689] : 
                  (N11779)? mem[691] : 
                  (N11781)? mem[693] : 
                  (N11783)? mem[695] : 
                  (N11785)? mem[697] : 
                  (N11787)? mem[699] : 
                  (N11789)? mem[701] : 
                  (N11791)? mem[703] : 
                  (N11793)? mem[705] : 
                  (N11795)? mem[707] : 
                  (N11797)? mem[709] : 
                  (N11799)? mem[711] : 
                  (N11801)? mem[713] : 
                  (N11803)? mem[715] : 
                  (N11805)? mem[717] : 
                  (N11807)? mem[719] : 
                  (N11809)? mem[721] : 
                  (N11811)? mem[723] : 
                  (N11813)? mem[725] : 
                  (N11815)? mem[727] : 
                  (N11817)? mem[729] : 
                  (N11819)? mem[731] : 
                  (N11821)? mem[733] : 
                  (N11823)? mem[735] : 
                  (N11825)? mem[737] : 
                  (N11827)? mem[739] : 
                  (N11829)? mem[741] : 
                  (N11831)? mem[743] : 
                  (N11833)? mem[745] : 
                  (N11835)? mem[747] : 
                  (N11837)? mem[749] : 
                  (N11839)? mem[751] : 
                  (N11841)? mem[753] : 
                  (N11843)? mem[755] : 
                  (N11845)? mem[757] : 
                  (N11847)? mem[759] : 
                  (N11849)? mem[761] : 
                  (N11851)? mem[763] : 
                  (N11853)? mem[765] : 
                  (N11855)? mem[767] : 
                  (N11857)? mem[769] : 
                  (N11859)? mem[771] : 
                  (N11861)? mem[773] : 
                  (N11863)? mem[775] : 
                  (N11865)? mem[777] : 
                  (N11867)? mem[779] : 
                  (N11869)? mem[781] : 
                  (N11871)? mem[783] : 
                  (N11873)? mem[785] : 
                  (N11875)? mem[787] : 
                  (N11877)? mem[789] : 
                  (N11879)? mem[791] : 
                  (N11881)? mem[793] : 
                  (N11883)? mem[795] : 
                  (N11885)? mem[797] : 
                  (N11887)? mem[799] : 
                  (N11889)? mem[801] : 
                  (N11891)? mem[803] : 
                  (N11893)? mem[805] : 
                  (N11895)? mem[807] : 
                  (N11897)? mem[809] : 
                  (N11899)? mem[811] : 
                  (N11901)? mem[813] : 
                  (N11903)? mem[815] : 
                  (N11905)? mem[817] : 
                  (N11907)? mem[819] : 
                  (N11909)? mem[821] : 
                  (N11911)? mem[823] : 
                  (N11913)? mem[825] : 
                  (N11915)? mem[827] : 
                  (N11917)? mem[829] : 
                  (N11919)? mem[831] : 
                  (N11921)? mem[833] : 
                  (N11923)? mem[835] : 
                  (N11925)? mem[837] : 
                  (N11927)? mem[839] : 
                  (N11929)? mem[841] : 
                  (N11931)? mem[843] : 
                  (N11933)? mem[845] : 
                  (N11935)? mem[847] : 
                  (N11937)? mem[849] : 
                  (N11939)? mem[851] : 
                  (N11941)? mem[853] : 
                  (N11943)? mem[855] : 
                  (N11945)? mem[857] : 
                  (N11947)? mem[859] : 
                  (N11949)? mem[861] : 
                  (N11951)? mem[863] : 
                  (N11953)? mem[865] : 
                  (N11955)? mem[867] : 
                  (N11957)? mem[869] : 
                  (N11959)? mem[871] : 
                  (N11961)? mem[873] : 
                  (N11963)? mem[875] : 
                  (N11965)? mem[877] : 
                  (N11967)? mem[879] : 
                  (N11969)? mem[881] : 
                  (N11971)? mem[883] : 
                  (N11973)? mem[885] : 
                  (N11975)? mem[887] : 
                  (N11977)? mem[889] : 
                  (N11979)? mem[891] : 
                  (N11981)? mem[893] : 
                  (N11983)? mem[895] : 
                  (N11985)? mem[897] : 
                  (N11987)? mem[899] : 
                  (N11989)? mem[901] : 
                  (N11991)? mem[903] : 
                  (N11993)? mem[905] : 
                  (N11995)? mem[907] : 
                  (N11997)? mem[909] : 
                  (N11999)? mem[911] : 
                  (N12001)? mem[913] : 
                  (N12003)? mem[915] : 
                  (N12005)? mem[917] : 
                  (N12007)? mem[919] : 
                  (N12009)? mem[921] : 
                  (N12011)? mem[923] : 
                  (N12013)? mem[925] : 
                  (N12015)? mem[927] : 
                  (N12017)? mem[929] : 
                  (N12019)? mem[931] : 
                  (N12021)? mem[933] : 
                  (N12023)? mem[935] : 
                  (N12025)? mem[937] : 
                  (N12027)? mem[939] : 
                  (N12029)? mem[941] : 
                  (N12031)? mem[943] : 
                  (N12033)? mem[945] : 
                  (N12035)? mem[947] : 
                  (N12037)? mem[949] : 
                  (N12039)? mem[951] : 
                  (N12041)? mem[953] : 
                  (N12043)? mem[955] : 
                  (N12045)? mem[957] : 
                  (N12047)? mem[959] : 
                  (N12049)? mem[961] : 
                  (N12051)? mem[963] : 
                  (N12053)? mem[965] : 
                  (N12055)? mem[967] : 
                  (N12057)? mem[969] : 
                  (N12059)? mem[971] : 
                  (N12061)? mem[973] : 
                  (N12063)? mem[975] : 
                  (N12065)? mem[977] : 
                  (N12067)? mem[979] : 
                  (N12069)? mem[981] : 
                  (N12071)? mem[983] : 
                  (N12073)? mem[985] : 
                  (N12075)? mem[987] : 
                  (N12077)? mem[989] : 
                  (N12079)? mem[991] : 
                  (N12081)? mem[993] : 
                  (N12083)? mem[995] : 
                  (N12085)? mem[997] : 
                  (N12087)? mem[999] : 
                  (N12089)? mem[1001] : 
                  (N12091)? mem[1003] : 
                  (N12093)? mem[1005] : 
                  (N12095)? mem[1007] : 
                  (N12097)? mem[1009] : 
                  (N12099)? mem[1011] : 
                  (N12101)? mem[1013] : 
                  (N12103)? mem[1015] : 
                  (N12105)? mem[1017] : 
                  (N12107)? mem[1019] : 
                  (N12109)? mem[1021] : 
                  (N12111)? mem[1023] : 1'b0;
  assign N12817 = (N12369)? mem[0] : 
                  (N12371)? mem[2] : 
                  (N12373)? mem[4] : 
                  (N12375)? mem[6] : 
                  (N12377)? mem[8] : 
                  (N12379)? mem[10] : 
                  (N12381)? mem[12] : 
                  (N12383)? mem[14] : 
                  (N12385)? mem[16] : 
                  (N12387)? mem[18] : 
                  (N12389)? mem[20] : 
                  (N12391)? mem[22] : 
                  (N12393)? mem[24] : 
                  (N12395)? mem[26] : 
                  (N12397)? mem[28] : 
                  (N12399)? mem[30] : 
                  (N12401)? mem[32] : 
                  (N12403)? mem[34] : 
                  (N12405)? mem[36] : 
                  (N12407)? mem[38] : 
                  (N12409)? mem[40] : 
                  (N12411)? mem[42] : 
                  (N12413)? mem[44] : 
                  (N12415)? mem[46] : 
                  (N12417)? mem[48] : 
                  (N12419)? mem[50] : 
                  (N12421)? mem[52] : 
                  (N12423)? mem[54] : 
                  (N12425)? mem[56] : 
                  (N12427)? mem[58] : 
                  (N12429)? mem[60] : 
                  (N12431)? mem[62] : 
                  (N12433)? mem[64] : 
                  (N12435)? mem[66] : 
                  (N12437)? mem[68] : 
                  (N12439)? mem[70] : 
                  (N12441)? mem[72] : 
                  (N12443)? mem[74] : 
                  (N12445)? mem[76] : 
                  (N12447)? mem[78] : 
                  (N12449)? mem[80] : 
                  (N12451)? mem[82] : 
                  (N12453)? mem[84] : 
                  (N12455)? mem[86] : 
                  (N12457)? mem[88] : 
                  (N12459)? mem[90] : 
                  (N12461)? mem[92] : 
                  (N12463)? mem[94] : 
                  (N12465)? mem[96] : 
                  (N12467)? mem[98] : 
                  (N12469)? mem[100] : 
                  (N12471)? mem[102] : 
                  (N12473)? mem[104] : 
                  (N12475)? mem[106] : 
                  (N12477)? mem[108] : 
                  (N12479)? mem[110] : 
                  (N12481)? mem[112] : 
                  (N12483)? mem[114] : 
                  (N12485)? mem[116] : 
                  (N12487)? mem[118] : 
                  (N12489)? mem[120] : 
                  (N12491)? mem[122] : 
                  (N12493)? mem[124] : 
                  (N12495)? mem[126] : 
                  (N12497)? mem[128] : 
                  (N12499)? mem[130] : 
                  (N12501)? mem[132] : 
                  (N12503)? mem[134] : 
                  (N12505)? mem[136] : 
                  (N12507)? mem[138] : 
                  (N12509)? mem[140] : 
                  (N12511)? mem[142] : 
                  (N12513)? mem[144] : 
                  (N12515)? mem[146] : 
                  (N12517)? mem[148] : 
                  (N12519)? mem[150] : 
                  (N12521)? mem[152] : 
                  (N12523)? mem[154] : 
                  (N12525)? mem[156] : 
                  (N12527)? mem[158] : 
                  (N12529)? mem[160] : 
                  (N12531)? mem[162] : 
                  (N12533)? mem[164] : 
                  (N12535)? mem[166] : 
                  (N12537)? mem[168] : 
                  (N12539)? mem[170] : 
                  (N12541)? mem[172] : 
                  (N12543)? mem[174] : 
                  (N12545)? mem[176] : 
                  (N12547)? mem[178] : 
                  (N12549)? mem[180] : 
                  (N12551)? mem[182] : 
                  (N12553)? mem[184] : 
                  (N12555)? mem[186] : 
                  (N12557)? mem[188] : 
                  (N12559)? mem[190] : 
                  (N12561)? mem[192] : 
                  (N12563)? mem[194] : 
                  (N12565)? mem[196] : 
                  (N12567)? mem[198] : 
                  (N12569)? mem[200] : 
                  (N12571)? mem[202] : 
                  (N12573)? mem[204] : 
                  (N12575)? mem[206] : 
                  (N12577)? mem[208] : 
                  (N12579)? mem[210] : 
                  (N12581)? mem[212] : 
                  (N12583)? mem[214] : 
                  (N12585)? mem[216] : 
                  (N12587)? mem[218] : 
                  (N12589)? mem[220] : 
                  (N12591)? mem[222] : 
                  (N12593)? mem[224] : 
                  (N12595)? mem[226] : 
                  (N12597)? mem[228] : 
                  (N12599)? mem[230] : 
                  (N12601)? mem[232] : 
                  (N12603)? mem[234] : 
                  (N12605)? mem[236] : 
                  (N12607)? mem[238] : 
                  (N12609)? mem[240] : 
                  (N12611)? mem[242] : 
                  (N12613)? mem[244] : 
                  (N12615)? mem[246] : 
                  (N12617)? mem[248] : 
                  (N12619)? mem[250] : 
                  (N12621)? mem[252] : 
                  (N12623)? mem[254] : 
                  (N12625)? mem[256] : 
                  (N12627)? mem[258] : 
                  (N12629)? mem[260] : 
                  (N12631)? mem[262] : 
                  (N12633)? mem[264] : 
                  (N12635)? mem[266] : 
                  (N12637)? mem[268] : 
                  (N12639)? mem[270] : 
                  (N12641)? mem[272] : 
                  (N12643)? mem[274] : 
                  (N12645)? mem[276] : 
                  (N12647)? mem[278] : 
                  (N12649)? mem[280] : 
                  (N12651)? mem[282] : 
                  (N12653)? mem[284] : 
                  (N12655)? mem[286] : 
                  (N12657)? mem[288] : 
                  (N12659)? mem[290] : 
                  (N12661)? mem[292] : 
                  (N12663)? mem[294] : 
                  (N12665)? mem[296] : 
                  (N12667)? mem[298] : 
                  (N12669)? mem[300] : 
                  (N12671)? mem[302] : 
                  (N12673)? mem[304] : 
                  (N12675)? mem[306] : 
                  (N12677)? mem[308] : 
                  (N12679)? mem[310] : 
                  (N12681)? mem[312] : 
                  (N12683)? mem[314] : 
                  (N12685)? mem[316] : 
                  (N12687)? mem[318] : 
                  (N12689)? mem[320] : 
                  (N12691)? mem[322] : 
                  (N12693)? mem[324] : 
                  (N12695)? mem[326] : 
                  (N12697)? mem[328] : 
                  (N12699)? mem[330] : 
                  (N12701)? mem[332] : 
                  (N12703)? mem[334] : 
                  (N12705)? mem[336] : 
                  (N12707)? mem[338] : 
                  (N12709)? mem[340] : 
                  (N12711)? mem[342] : 
                  (N12713)? mem[344] : 
                  (N12715)? mem[346] : 
                  (N12717)? mem[348] : 
                  (N12719)? mem[350] : 
                  (N12721)? mem[352] : 
                  (N12723)? mem[354] : 
                  (N12725)? mem[356] : 
                  (N12727)? mem[358] : 
                  (N12729)? mem[360] : 
                  (N12731)? mem[362] : 
                  (N12733)? mem[364] : 
                  (N12735)? mem[366] : 
                  (N12737)? mem[368] : 
                  (N12739)? mem[370] : 
                  (N12741)? mem[372] : 
                  (N12743)? mem[374] : 
                  (N12745)? mem[376] : 
                  (N12747)? mem[378] : 
                  (N12749)? mem[380] : 
                  (N12751)? mem[382] : 
                  (N12753)? mem[384] : 
                  (N12754)? mem[386] : 
                  (N12755)? mem[388] : 
                  (N12756)? mem[390] : 
                  (N12757)? mem[392] : 
                  (N12758)? mem[394] : 
                  (N12759)? mem[396] : 
                  (N12760)? mem[398] : 
                  (N12761)? mem[400] : 
                  (N12762)? mem[402] : 
                  (N12763)? mem[404] : 
                  (N12764)? mem[406] : 
                  (N12765)? mem[408] : 
                  (N12766)? mem[410] : 
                  (N12767)? mem[412] : 
                  (N12768)? mem[414] : 
                  (N12769)? mem[416] : 
                  (N12770)? mem[418] : 
                  (N12771)? mem[420] : 
                  (N12772)? mem[422] : 
                  (N12773)? mem[424] : 
                  (N12774)? mem[426] : 
                  (N12775)? mem[428] : 
                  (N12776)? mem[430] : 
                  (N12777)? mem[432] : 
                  (N12778)? mem[434] : 
                  (N12779)? mem[436] : 
                  (N12780)? mem[438] : 
                  (N12781)? mem[440] : 
                  (N12782)? mem[442] : 
                  (N12783)? mem[444] : 
                  (N12784)? mem[446] : 
                  (N12785)? mem[448] : 
                  (N12786)? mem[450] : 
                  (N12787)? mem[452] : 
                  (N12788)? mem[454] : 
                  (N12789)? mem[456] : 
                  (N12790)? mem[458] : 
                  (N12791)? mem[460] : 
                  (N12792)? mem[462] : 
                  (N12793)? mem[464] : 
                  (N12794)? mem[466] : 
                  (N12795)? mem[468] : 
                  (N12796)? mem[470] : 
                  (N12797)? mem[472] : 
                  (N12798)? mem[474] : 
                  (N12799)? mem[476] : 
                  (N12800)? mem[478] : 
                  (N12801)? mem[480] : 
                  (N12802)? mem[482] : 
                  (N12803)? mem[484] : 
                  (N12804)? mem[486] : 
                  (N12805)? mem[488] : 
                  (N12806)? mem[490] : 
                  (N12807)? mem[492] : 
                  (N12808)? mem[494] : 
                  (N12809)? mem[496] : 
                  (N12810)? mem[498] : 
                  (N12811)? mem[500] : 
                  (N12812)? mem[502] : 
                  (N12813)? mem[504] : 
                  (N12814)? mem[506] : 
                  (N12815)? mem[508] : 
                  (N12816)? mem[510] : 
                  (N12370)? mem[512] : 
                  (N12372)? mem[514] : 
                  (N12374)? mem[516] : 
                  (N12376)? mem[518] : 
                  (N12378)? mem[520] : 
                  (N12380)? mem[522] : 
                  (N12382)? mem[524] : 
                  (N12384)? mem[526] : 
                  (N12386)? mem[528] : 
                  (N12388)? mem[530] : 
                  (N12390)? mem[532] : 
                  (N12392)? mem[534] : 
                  (N12394)? mem[536] : 
                  (N12396)? mem[538] : 
                  (N12398)? mem[540] : 
                  (N12400)? mem[542] : 
                  (N12402)? mem[544] : 
                  (N12404)? mem[546] : 
                  (N12406)? mem[548] : 
                  (N12408)? mem[550] : 
                  (N12410)? mem[552] : 
                  (N12412)? mem[554] : 
                  (N12414)? mem[556] : 
                  (N12416)? mem[558] : 
                  (N12418)? mem[560] : 
                  (N12420)? mem[562] : 
                  (N12422)? mem[564] : 
                  (N12424)? mem[566] : 
                  (N12426)? mem[568] : 
                  (N12428)? mem[570] : 
                  (N12430)? mem[572] : 
                  (N12432)? mem[574] : 
                  (N12434)? mem[576] : 
                  (N12436)? mem[578] : 
                  (N12438)? mem[580] : 
                  (N12440)? mem[582] : 
                  (N12442)? mem[584] : 
                  (N12444)? mem[586] : 
                  (N12446)? mem[588] : 
                  (N12448)? mem[590] : 
                  (N12450)? mem[592] : 
                  (N12452)? mem[594] : 
                  (N12454)? mem[596] : 
                  (N12456)? mem[598] : 
                  (N12458)? mem[600] : 
                  (N12460)? mem[602] : 
                  (N12462)? mem[604] : 
                  (N12464)? mem[606] : 
                  (N12466)? mem[608] : 
                  (N12468)? mem[610] : 
                  (N12470)? mem[612] : 
                  (N12472)? mem[614] : 
                  (N12474)? mem[616] : 
                  (N12476)? mem[618] : 
                  (N12478)? mem[620] : 
                  (N12480)? mem[622] : 
                  (N12482)? mem[624] : 
                  (N12484)? mem[626] : 
                  (N12486)? mem[628] : 
                  (N12488)? mem[630] : 
                  (N12490)? mem[632] : 
                  (N12492)? mem[634] : 
                  (N12494)? mem[636] : 
                  (N12496)? mem[638] : 
                  (N12498)? mem[640] : 
                  (N12500)? mem[642] : 
                  (N12502)? mem[644] : 
                  (N12504)? mem[646] : 
                  (N12506)? mem[648] : 
                  (N12508)? mem[650] : 
                  (N12510)? mem[652] : 
                  (N12512)? mem[654] : 
                  (N12514)? mem[656] : 
                  (N12516)? mem[658] : 
                  (N12518)? mem[660] : 
                  (N12520)? mem[662] : 
                  (N12522)? mem[664] : 
                  (N12524)? mem[666] : 
                  (N12526)? mem[668] : 
                  (N12528)? mem[670] : 
                  (N12530)? mem[672] : 
                  (N12532)? mem[674] : 
                  (N12534)? mem[676] : 
                  (N12536)? mem[678] : 
                  (N12538)? mem[680] : 
                  (N12540)? mem[682] : 
                  (N12542)? mem[684] : 
                  (N12544)? mem[686] : 
                  (N12546)? mem[688] : 
                  (N12548)? mem[690] : 
                  (N12550)? mem[692] : 
                  (N12552)? mem[694] : 
                  (N12554)? mem[696] : 
                  (N12556)? mem[698] : 
                  (N12558)? mem[700] : 
                  (N12560)? mem[702] : 
                  (N12562)? mem[704] : 
                  (N12564)? mem[706] : 
                  (N12566)? mem[708] : 
                  (N12568)? mem[710] : 
                  (N12570)? mem[712] : 
                  (N12572)? mem[714] : 
                  (N12574)? mem[716] : 
                  (N12576)? mem[718] : 
                  (N12578)? mem[720] : 
                  (N12580)? mem[722] : 
                  (N12582)? mem[724] : 
                  (N12584)? mem[726] : 
                  (N12586)? mem[728] : 
                  (N12588)? mem[730] : 
                  (N12590)? mem[732] : 
                  (N12592)? mem[734] : 
                  (N12594)? mem[736] : 
                  (N12596)? mem[738] : 
                  (N12598)? mem[740] : 
                  (N12600)? mem[742] : 
                  (N12602)? mem[744] : 
                  (N12604)? mem[746] : 
                  (N12606)? mem[748] : 
                  (N12608)? mem[750] : 
                  (N12610)? mem[752] : 
                  (N12612)? mem[754] : 
                  (N12614)? mem[756] : 
                  (N12616)? mem[758] : 
                  (N12618)? mem[760] : 
                  (N12620)? mem[762] : 
                  (N12622)? mem[764] : 
                  (N12624)? mem[766] : 
                  (N12626)? mem[768] : 
                  (N12628)? mem[770] : 
                  (N12630)? mem[772] : 
                  (N12632)? mem[774] : 
                  (N12634)? mem[776] : 
                  (N12636)? mem[778] : 
                  (N12638)? mem[780] : 
                  (N12640)? mem[782] : 
                  (N12642)? mem[784] : 
                  (N12644)? mem[786] : 
                  (N12646)? mem[788] : 
                  (N12648)? mem[790] : 
                  (N12650)? mem[792] : 
                  (N12652)? mem[794] : 
                  (N12654)? mem[796] : 
                  (N12656)? mem[798] : 
                  (N12658)? mem[800] : 
                  (N12660)? mem[802] : 
                  (N12662)? mem[804] : 
                  (N12664)? mem[806] : 
                  (N12666)? mem[808] : 
                  (N12668)? mem[810] : 
                  (N12670)? mem[812] : 
                  (N12672)? mem[814] : 
                  (N12674)? mem[816] : 
                  (N12676)? mem[818] : 
                  (N12678)? mem[820] : 
                  (N12680)? mem[822] : 
                  (N12682)? mem[824] : 
                  (N12684)? mem[826] : 
                  (N12686)? mem[828] : 
                  (N12688)? mem[830] : 
                  (N12690)? mem[832] : 
                  (N12692)? mem[834] : 
                  (N12694)? mem[836] : 
                  (N12696)? mem[838] : 
                  (N12698)? mem[840] : 
                  (N12700)? mem[842] : 
                  (N12702)? mem[844] : 
                  (N12704)? mem[846] : 
                  (N12706)? mem[848] : 
                  (N12708)? mem[850] : 
                  (N12710)? mem[852] : 
                  (N12712)? mem[854] : 
                  (N12714)? mem[856] : 
                  (N12716)? mem[858] : 
                  (N12718)? mem[860] : 
                  (N12720)? mem[862] : 
                  (N12722)? mem[864] : 
                  (N12724)? mem[866] : 
                  (N12726)? mem[868] : 
                  (N12728)? mem[870] : 
                  (N12730)? mem[872] : 
                  (N12732)? mem[874] : 
                  (N12734)? mem[876] : 
                  (N12736)? mem[878] : 
                  (N12738)? mem[880] : 
                  (N12740)? mem[882] : 
                  (N12742)? mem[884] : 
                  (N12744)? mem[886] : 
                  (N12746)? mem[888] : 
                  (N12748)? mem[890] : 
                  (N12750)? mem[892] : 
                  (N12752)? mem[894] : 
                  (N10992)? mem[896] : 
                  (N10994)? mem[898] : 
                  (N10996)? mem[900] : 
                  (N10998)? mem[902] : 
                  (N11000)? mem[904] : 
                  (N11002)? mem[906] : 
                  (N11004)? mem[908] : 
                  (N11006)? mem[910] : 
                  (N11008)? mem[912] : 
                  (N11010)? mem[914] : 
                  (N11012)? mem[916] : 
                  (N11014)? mem[918] : 
                  (N11016)? mem[920] : 
                  (N11018)? mem[922] : 
                  (N11020)? mem[924] : 
                  (N11022)? mem[926] : 
                  (N11024)? mem[928] : 
                  (N11026)? mem[930] : 
                  (N11028)? mem[932] : 
                  (N11030)? mem[934] : 
                  (N11032)? mem[936] : 
                  (N11034)? mem[938] : 
                  (N11036)? mem[940] : 
                  (N11038)? mem[942] : 
                  (N11040)? mem[944] : 
                  (N11042)? mem[946] : 
                  (N11044)? mem[948] : 
                  (N11046)? mem[950] : 
                  (N11048)? mem[952] : 
                  (N11050)? mem[954] : 
                  (N11052)? mem[956] : 
                  (N11054)? mem[958] : 
                  (N12049)? mem[960] : 
                  (N12051)? mem[962] : 
                  (N12053)? mem[964] : 
                  (N12055)? mem[966] : 
                  (N12057)? mem[968] : 
                  (N12059)? mem[970] : 
                  (N12061)? mem[972] : 
                  (N12063)? mem[974] : 
                  (N12065)? mem[976] : 
                  (N12067)? mem[978] : 
                  (N12069)? mem[980] : 
                  (N12071)? mem[982] : 
                  (N12073)? mem[984] : 
                  (N12075)? mem[986] : 
                  (N12077)? mem[988] : 
                  (N12079)? mem[990] : 
                  (N12081)? mem[992] : 
                  (N12083)? mem[994] : 
                  (N12085)? mem[996] : 
                  (N12087)? mem[998] : 
                  (N12089)? mem[1000] : 
                  (N12091)? mem[1002] : 
                  (N12093)? mem[1004] : 
                  (N12095)? mem[1006] : 
                  (N12097)? mem[1008] : 
                  (N12099)? mem[1010] : 
                  (N12101)? mem[1012] : 
                  (N12103)? mem[1014] : 
                  (N12105)? mem[1016] : 
                  (N12107)? mem[1018] : 
                  (N12109)? mem[1020] : 
                  (N12111)? mem[1022] : 1'b0;
  assign N13523 = (N13075)? mem[1] : 
                  (N13077)? mem[3] : 
                  (N13079)? mem[5] : 
                  (N13081)? mem[7] : 
                  (N13083)? mem[9] : 
                  (N13085)? mem[11] : 
                  (N13087)? mem[13] : 
                  (N13089)? mem[15] : 
                  (N13091)? mem[17] : 
                  (N13093)? mem[19] : 
                  (N13095)? mem[21] : 
                  (N13097)? mem[23] : 
                  (N13099)? mem[25] : 
                  (N13101)? mem[27] : 
                  (N13103)? mem[29] : 
                  (N13105)? mem[31] : 
                  (N13107)? mem[33] : 
                  (N13109)? mem[35] : 
                  (N13111)? mem[37] : 
                  (N13113)? mem[39] : 
                  (N13115)? mem[41] : 
                  (N13117)? mem[43] : 
                  (N13119)? mem[45] : 
                  (N13121)? mem[47] : 
                  (N13123)? mem[49] : 
                  (N13125)? mem[51] : 
                  (N13127)? mem[53] : 
                  (N13129)? mem[55] : 
                  (N13131)? mem[57] : 
                  (N13133)? mem[59] : 
                  (N13135)? mem[61] : 
                  (N13137)? mem[63] : 
                  (N13139)? mem[65] : 
                  (N13141)? mem[67] : 
                  (N13143)? mem[69] : 
                  (N13145)? mem[71] : 
                  (N13147)? mem[73] : 
                  (N13149)? mem[75] : 
                  (N13151)? mem[77] : 
                  (N13153)? mem[79] : 
                  (N13155)? mem[81] : 
                  (N13157)? mem[83] : 
                  (N13159)? mem[85] : 
                  (N13161)? mem[87] : 
                  (N13163)? mem[89] : 
                  (N13165)? mem[91] : 
                  (N13167)? mem[93] : 
                  (N13169)? mem[95] : 
                  (N13171)? mem[97] : 
                  (N13173)? mem[99] : 
                  (N13175)? mem[101] : 
                  (N13177)? mem[103] : 
                  (N13179)? mem[105] : 
                  (N13181)? mem[107] : 
                  (N13183)? mem[109] : 
                  (N13185)? mem[111] : 
                  (N13187)? mem[113] : 
                  (N13189)? mem[115] : 
                  (N13191)? mem[117] : 
                  (N13193)? mem[119] : 
                  (N13195)? mem[121] : 
                  (N13197)? mem[123] : 
                  (N13199)? mem[125] : 
                  (N13201)? mem[127] : 
                  (N13203)? mem[129] : 
                  (N13205)? mem[131] : 
                  (N13207)? mem[133] : 
                  (N13209)? mem[135] : 
                  (N13211)? mem[137] : 
                  (N13213)? mem[139] : 
                  (N13215)? mem[141] : 
                  (N13217)? mem[143] : 
                  (N13219)? mem[145] : 
                  (N13221)? mem[147] : 
                  (N13223)? mem[149] : 
                  (N13225)? mem[151] : 
                  (N13227)? mem[153] : 
                  (N13229)? mem[155] : 
                  (N13231)? mem[157] : 
                  (N13233)? mem[159] : 
                  (N13235)? mem[161] : 
                  (N13237)? mem[163] : 
                  (N13239)? mem[165] : 
                  (N13241)? mem[167] : 
                  (N13243)? mem[169] : 
                  (N13245)? mem[171] : 
                  (N13247)? mem[173] : 
                  (N13249)? mem[175] : 
                  (N13251)? mem[177] : 
                  (N13253)? mem[179] : 
                  (N13255)? mem[181] : 
                  (N13257)? mem[183] : 
                  (N13259)? mem[185] : 
                  (N13261)? mem[187] : 
                  (N13263)? mem[189] : 
                  (N13265)? mem[191] : 
                  (N13267)? mem[193] : 
                  (N13269)? mem[195] : 
                  (N13271)? mem[197] : 
                  (N13273)? mem[199] : 
                  (N13275)? mem[201] : 
                  (N13277)? mem[203] : 
                  (N13279)? mem[205] : 
                  (N13281)? mem[207] : 
                  (N13283)? mem[209] : 
                  (N13285)? mem[211] : 
                  (N13287)? mem[213] : 
                  (N13289)? mem[215] : 
                  (N13291)? mem[217] : 
                  (N13293)? mem[219] : 
                  (N13295)? mem[221] : 
                  (N13297)? mem[223] : 
                  (N13299)? mem[225] : 
                  (N13301)? mem[227] : 
                  (N13303)? mem[229] : 
                  (N13305)? mem[231] : 
                  (N13307)? mem[233] : 
                  (N13309)? mem[235] : 
                  (N13311)? mem[237] : 
                  (N13313)? mem[239] : 
                  (N13315)? mem[241] : 
                  (N13317)? mem[243] : 
                  (N13319)? mem[245] : 
                  (N13321)? mem[247] : 
                  (N13323)? mem[249] : 
                  (N13325)? mem[251] : 
                  (N13327)? mem[253] : 
                  (N13329)? mem[255] : 
                  (N13331)? mem[257] : 
                  (N13333)? mem[259] : 
                  (N13335)? mem[261] : 
                  (N13337)? mem[263] : 
                  (N13339)? mem[265] : 
                  (N13341)? mem[267] : 
                  (N13343)? mem[269] : 
                  (N13345)? mem[271] : 
                  (N13347)? mem[273] : 
                  (N13349)? mem[275] : 
                  (N13351)? mem[277] : 
                  (N13353)? mem[279] : 
                  (N13355)? mem[281] : 
                  (N13357)? mem[283] : 
                  (N13359)? mem[285] : 
                  (N13361)? mem[287] : 
                  (N13363)? mem[289] : 
                  (N13365)? mem[291] : 
                  (N13367)? mem[293] : 
                  (N13369)? mem[295] : 
                  (N13371)? mem[297] : 
                  (N13373)? mem[299] : 
                  (N13375)? mem[301] : 
                  (N13377)? mem[303] : 
                  (N13379)? mem[305] : 
                  (N13381)? mem[307] : 
                  (N13383)? mem[309] : 
                  (N13385)? mem[311] : 
                  (N13387)? mem[313] : 
                  (N13389)? mem[315] : 
                  (N13391)? mem[317] : 
                  (N13393)? mem[319] : 
                  (N13395)? mem[321] : 
                  (N13397)? mem[323] : 
                  (N13399)? mem[325] : 
                  (N13401)? mem[327] : 
                  (N13403)? mem[329] : 
                  (N13405)? mem[331] : 
                  (N13407)? mem[333] : 
                  (N13409)? mem[335] : 
                  (N13411)? mem[337] : 
                  (N13413)? mem[339] : 
                  (N13415)? mem[341] : 
                  (N13417)? mem[343] : 
                  (N13419)? mem[345] : 
                  (N13421)? mem[347] : 
                  (N13423)? mem[349] : 
                  (N13425)? mem[351] : 
                  (N13427)? mem[353] : 
                  (N13429)? mem[355] : 
                  (N13431)? mem[357] : 
                  (N13433)? mem[359] : 
                  (N13435)? mem[361] : 
                  (N13437)? mem[363] : 
                  (N13439)? mem[365] : 
                  (N13441)? mem[367] : 
                  (N13443)? mem[369] : 
                  (N13445)? mem[371] : 
                  (N13447)? mem[373] : 
                  (N13449)? mem[375] : 
                  (N13451)? mem[377] : 
                  (N13453)? mem[379] : 
                  (N13455)? mem[381] : 
                  (N13457)? mem[383] : 
                  (N13459)? mem[385] : 
                  (N13460)? mem[387] : 
                  (N13461)? mem[389] : 
                  (N13462)? mem[391] : 
                  (N13463)? mem[393] : 
                  (N13464)? mem[395] : 
                  (N13465)? mem[397] : 
                  (N13466)? mem[399] : 
                  (N13467)? mem[401] : 
                  (N13468)? mem[403] : 
                  (N13469)? mem[405] : 
                  (N13470)? mem[407] : 
                  (N13471)? mem[409] : 
                  (N13472)? mem[411] : 
                  (N13473)? mem[413] : 
                  (N13474)? mem[415] : 
                  (N13475)? mem[417] : 
                  (N13476)? mem[419] : 
                  (N13477)? mem[421] : 
                  (N13478)? mem[423] : 
                  (N13479)? mem[425] : 
                  (N13480)? mem[427] : 
                  (N13481)? mem[429] : 
                  (N13482)? mem[431] : 
                  (N13483)? mem[433] : 
                  (N13484)? mem[435] : 
                  (N13485)? mem[437] : 
                  (N13486)? mem[439] : 
                  (N13487)? mem[441] : 
                  (N13488)? mem[443] : 
                  (N13489)? mem[445] : 
                  (N13490)? mem[447] : 
                  (N13491)? mem[449] : 
                  (N13492)? mem[451] : 
                  (N13493)? mem[453] : 
                  (N13494)? mem[455] : 
                  (N13495)? mem[457] : 
                  (N13496)? mem[459] : 
                  (N13497)? mem[461] : 
                  (N13498)? mem[463] : 
                  (N13499)? mem[465] : 
                  (N13500)? mem[467] : 
                  (N13501)? mem[469] : 
                  (N13502)? mem[471] : 
                  (N13503)? mem[473] : 
                  (N13504)? mem[475] : 
                  (N13505)? mem[477] : 
                  (N13506)? mem[479] : 
                  (N13507)? mem[481] : 
                  (N13508)? mem[483] : 
                  (N13509)? mem[485] : 
                  (N13510)? mem[487] : 
                  (N13511)? mem[489] : 
                  (N13512)? mem[491] : 
                  (N13513)? mem[493] : 
                  (N13514)? mem[495] : 
                  (N13515)? mem[497] : 
                  (N13516)? mem[499] : 
                  (N13517)? mem[501] : 
                  (N13518)? mem[503] : 
                  (N13519)? mem[505] : 
                  (N13520)? mem[507] : 
                  (N13521)? mem[509] : 
                  (N13522)? mem[511] : 
                  (N13076)? mem[513] : 
                  (N13078)? mem[515] : 
                  (N13080)? mem[517] : 
                  (N13082)? mem[519] : 
                  (N13084)? mem[521] : 
                  (N13086)? mem[523] : 
                  (N13088)? mem[525] : 
                  (N13090)? mem[527] : 
                  (N13092)? mem[529] : 
                  (N13094)? mem[531] : 
                  (N13096)? mem[533] : 
                  (N13098)? mem[535] : 
                  (N13100)? mem[537] : 
                  (N13102)? mem[539] : 
                  (N13104)? mem[541] : 
                  (N13106)? mem[543] : 
                  (N13108)? mem[545] : 
                  (N13110)? mem[547] : 
                  (N13112)? mem[549] : 
                  (N13114)? mem[551] : 
                  (N13116)? mem[553] : 
                  (N13118)? mem[555] : 
                  (N13120)? mem[557] : 
                  (N13122)? mem[559] : 
                  (N13124)? mem[561] : 
                  (N13126)? mem[563] : 
                  (N13128)? mem[565] : 
                  (N13130)? mem[567] : 
                  (N13132)? mem[569] : 
                  (N13134)? mem[571] : 
                  (N13136)? mem[573] : 
                  (N13138)? mem[575] : 
                  (N13140)? mem[577] : 
                  (N13142)? mem[579] : 
                  (N13144)? mem[581] : 
                  (N13146)? mem[583] : 
                  (N13148)? mem[585] : 
                  (N13150)? mem[587] : 
                  (N13152)? mem[589] : 
                  (N13154)? mem[591] : 
                  (N13156)? mem[593] : 
                  (N13158)? mem[595] : 
                  (N13160)? mem[597] : 
                  (N13162)? mem[599] : 
                  (N13164)? mem[601] : 
                  (N13166)? mem[603] : 
                  (N13168)? mem[605] : 
                  (N13170)? mem[607] : 
                  (N13172)? mem[609] : 
                  (N13174)? mem[611] : 
                  (N13176)? mem[613] : 
                  (N13178)? mem[615] : 
                  (N13180)? mem[617] : 
                  (N13182)? mem[619] : 
                  (N13184)? mem[621] : 
                  (N13186)? mem[623] : 
                  (N13188)? mem[625] : 
                  (N13190)? mem[627] : 
                  (N13192)? mem[629] : 
                  (N13194)? mem[631] : 
                  (N13196)? mem[633] : 
                  (N13198)? mem[635] : 
                  (N13200)? mem[637] : 
                  (N13202)? mem[639] : 
                  (N13204)? mem[641] : 
                  (N13206)? mem[643] : 
                  (N13208)? mem[645] : 
                  (N13210)? mem[647] : 
                  (N13212)? mem[649] : 
                  (N13214)? mem[651] : 
                  (N13216)? mem[653] : 
                  (N13218)? mem[655] : 
                  (N13220)? mem[657] : 
                  (N13222)? mem[659] : 
                  (N13224)? mem[661] : 
                  (N13226)? mem[663] : 
                  (N13228)? mem[665] : 
                  (N13230)? mem[667] : 
                  (N13232)? mem[669] : 
                  (N13234)? mem[671] : 
                  (N13236)? mem[673] : 
                  (N13238)? mem[675] : 
                  (N13240)? mem[677] : 
                  (N13242)? mem[679] : 
                  (N13244)? mem[681] : 
                  (N13246)? mem[683] : 
                  (N13248)? mem[685] : 
                  (N13250)? mem[687] : 
                  (N13252)? mem[689] : 
                  (N13254)? mem[691] : 
                  (N13256)? mem[693] : 
                  (N13258)? mem[695] : 
                  (N13260)? mem[697] : 
                  (N13262)? mem[699] : 
                  (N13264)? mem[701] : 
                  (N13266)? mem[703] : 
                  (N13268)? mem[705] : 
                  (N13270)? mem[707] : 
                  (N13272)? mem[709] : 
                  (N13274)? mem[711] : 
                  (N13276)? mem[713] : 
                  (N13278)? mem[715] : 
                  (N13280)? mem[717] : 
                  (N13282)? mem[719] : 
                  (N13284)? mem[721] : 
                  (N13286)? mem[723] : 
                  (N13288)? mem[725] : 
                  (N13290)? mem[727] : 
                  (N13292)? mem[729] : 
                  (N13294)? mem[731] : 
                  (N13296)? mem[733] : 
                  (N13298)? mem[735] : 
                  (N13300)? mem[737] : 
                  (N13302)? mem[739] : 
                  (N13304)? mem[741] : 
                  (N13306)? mem[743] : 
                  (N13308)? mem[745] : 
                  (N13310)? mem[747] : 
                  (N13312)? mem[749] : 
                  (N13314)? mem[751] : 
                  (N13316)? mem[753] : 
                  (N13318)? mem[755] : 
                  (N13320)? mem[757] : 
                  (N13322)? mem[759] : 
                  (N13324)? mem[761] : 
                  (N13326)? mem[763] : 
                  (N13328)? mem[765] : 
                  (N13330)? mem[767] : 
                  (N13332)? mem[769] : 
                  (N13334)? mem[771] : 
                  (N13336)? mem[773] : 
                  (N13338)? mem[775] : 
                  (N13340)? mem[777] : 
                  (N13342)? mem[779] : 
                  (N13344)? mem[781] : 
                  (N13346)? mem[783] : 
                  (N13348)? mem[785] : 
                  (N13350)? mem[787] : 
                  (N13352)? mem[789] : 
                  (N13354)? mem[791] : 
                  (N13356)? mem[793] : 
                  (N13358)? mem[795] : 
                  (N13360)? mem[797] : 
                  (N13362)? mem[799] : 
                  (N13364)? mem[801] : 
                  (N13366)? mem[803] : 
                  (N13368)? mem[805] : 
                  (N13370)? mem[807] : 
                  (N13372)? mem[809] : 
                  (N13374)? mem[811] : 
                  (N13376)? mem[813] : 
                  (N13378)? mem[815] : 
                  (N13380)? mem[817] : 
                  (N13382)? mem[819] : 
                  (N13384)? mem[821] : 
                  (N13386)? mem[823] : 
                  (N13388)? mem[825] : 
                  (N13390)? mem[827] : 
                  (N13392)? mem[829] : 
                  (N13394)? mem[831] : 
                  (N13396)? mem[833] : 
                  (N13398)? mem[835] : 
                  (N13400)? mem[837] : 
                  (N13402)? mem[839] : 
                  (N13404)? mem[841] : 
                  (N13406)? mem[843] : 
                  (N13408)? mem[845] : 
                  (N13410)? mem[847] : 
                  (N13412)? mem[849] : 
                  (N13414)? mem[851] : 
                  (N13416)? mem[853] : 
                  (N13418)? mem[855] : 
                  (N13420)? mem[857] : 
                  (N13422)? mem[859] : 
                  (N13424)? mem[861] : 
                  (N13426)? mem[863] : 
                  (N13428)? mem[865] : 
                  (N13430)? mem[867] : 
                  (N13432)? mem[869] : 
                  (N13434)? mem[871] : 
                  (N13436)? mem[873] : 
                  (N13438)? mem[875] : 
                  (N13440)? mem[877] : 
                  (N13442)? mem[879] : 
                  (N13444)? mem[881] : 
                  (N13446)? mem[883] : 
                  (N13448)? mem[885] : 
                  (N13450)? mem[887] : 
                  (N13452)? mem[889] : 
                  (N13454)? mem[891] : 
                  (N13456)? mem[893] : 
                  (N13458)? mem[895] : 
                  (N10992)? mem[897] : 
                  (N10994)? mem[899] : 
                  (N10996)? mem[901] : 
                  (N10998)? mem[903] : 
                  (N11000)? mem[905] : 
                  (N11002)? mem[907] : 
                  (N11004)? mem[909] : 
                  (N11006)? mem[911] : 
                  (N11008)? mem[913] : 
                  (N11010)? mem[915] : 
                  (N11012)? mem[917] : 
                  (N11014)? mem[919] : 
                  (N11016)? mem[921] : 
                  (N11018)? mem[923] : 
                  (N11020)? mem[925] : 
                  (N11022)? mem[927] : 
                  (N11024)? mem[929] : 
                  (N11026)? mem[931] : 
                  (N11028)? mem[933] : 
                  (N11030)? mem[935] : 
                  (N11032)? mem[937] : 
                  (N11034)? mem[939] : 
                  (N11036)? mem[941] : 
                  (N11038)? mem[943] : 
                  (N11040)? mem[945] : 
                  (N11042)? mem[947] : 
                  (N11044)? mem[949] : 
                  (N11046)? mem[951] : 
                  (N11048)? mem[953] : 
                  (N11050)? mem[955] : 
                  (N11052)? mem[957] : 
                  (N11054)? mem[959] : 
                  (N12049)? mem[961] : 
                  (N12051)? mem[963] : 
                  (N12053)? mem[965] : 
                  (N12055)? mem[967] : 
                  (N12057)? mem[969] : 
                  (N12059)? mem[971] : 
                  (N12061)? mem[973] : 
                  (N12063)? mem[975] : 
                  (N12065)? mem[977] : 
                  (N12067)? mem[979] : 
                  (N12069)? mem[981] : 
                  (N12071)? mem[983] : 
                  (N12073)? mem[985] : 
                  (N12075)? mem[987] : 
                  (N12077)? mem[989] : 
                  (N12079)? mem[991] : 
                  (N12081)? mem[993] : 
                  (N12083)? mem[995] : 
                  (N12085)? mem[997] : 
                  (N12087)? mem[999] : 
                  (N12089)? mem[1001] : 
                  (N12091)? mem[1003] : 
                  (N12093)? mem[1005] : 
                  (N12095)? mem[1007] : 
                  (N12097)? mem[1009] : 
                  (N12099)? mem[1011] : 
                  (N12101)? mem[1013] : 
                  (N12103)? mem[1015] : 
                  (N12105)? mem[1017] : 
                  (N12107)? mem[1019] : 
                  (N12109)? mem[1021] : 
                  (N12111)? mem[1023] : 1'b0;
  assign N13524 = (N13075)? mem[0] : 
                  (N13077)? mem[2] : 
                  (N13079)? mem[4] : 
                  (N13081)? mem[6] : 
                  (N13083)? mem[8] : 
                  (N13085)? mem[10] : 
                  (N13087)? mem[12] : 
                  (N13089)? mem[14] : 
                  (N13091)? mem[16] : 
                  (N13093)? mem[18] : 
                  (N13095)? mem[20] : 
                  (N13097)? mem[22] : 
                  (N13099)? mem[24] : 
                  (N13101)? mem[26] : 
                  (N13103)? mem[28] : 
                  (N13105)? mem[30] : 
                  (N13107)? mem[32] : 
                  (N13109)? mem[34] : 
                  (N13111)? mem[36] : 
                  (N13113)? mem[38] : 
                  (N13115)? mem[40] : 
                  (N13117)? mem[42] : 
                  (N13119)? mem[44] : 
                  (N13121)? mem[46] : 
                  (N13123)? mem[48] : 
                  (N13125)? mem[50] : 
                  (N13127)? mem[52] : 
                  (N13129)? mem[54] : 
                  (N13131)? mem[56] : 
                  (N13133)? mem[58] : 
                  (N13135)? mem[60] : 
                  (N13137)? mem[62] : 
                  (N13139)? mem[64] : 
                  (N13141)? mem[66] : 
                  (N13143)? mem[68] : 
                  (N13145)? mem[70] : 
                  (N13147)? mem[72] : 
                  (N13149)? mem[74] : 
                  (N13151)? mem[76] : 
                  (N13153)? mem[78] : 
                  (N13155)? mem[80] : 
                  (N13157)? mem[82] : 
                  (N13159)? mem[84] : 
                  (N13161)? mem[86] : 
                  (N13163)? mem[88] : 
                  (N13165)? mem[90] : 
                  (N13167)? mem[92] : 
                  (N13169)? mem[94] : 
                  (N13171)? mem[96] : 
                  (N13173)? mem[98] : 
                  (N13175)? mem[100] : 
                  (N13177)? mem[102] : 
                  (N13179)? mem[104] : 
                  (N13181)? mem[106] : 
                  (N13183)? mem[108] : 
                  (N13185)? mem[110] : 
                  (N13187)? mem[112] : 
                  (N13189)? mem[114] : 
                  (N13191)? mem[116] : 
                  (N13193)? mem[118] : 
                  (N13195)? mem[120] : 
                  (N13197)? mem[122] : 
                  (N13199)? mem[124] : 
                  (N13201)? mem[126] : 
                  (N13203)? mem[128] : 
                  (N13205)? mem[130] : 
                  (N13207)? mem[132] : 
                  (N13209)? mem[134] : 
                  (N13211)? mem[136] : 
                  (N13213)? mem[138] : 
                  (N13215)? mem[140] : 
                  (N13217)? mem[142] : 
                  (N13219)? mem[144] : 
                  (N13221)? mem[146] : 
                  (N13223)? mem[148] : 
                  (N13225)? mem[150] : 
                  (N13227)? mem[152] : 
                  (N13229)? mem[154] : 
                  (N13231)? mem[156] : 
                  (N13233)? mem[158] : 
                  (N13235)? mem[160] : 
                  (N13237)? mem[162] : 
                  (N13239)? mem[164] : 
                  (N13241)? mem[166] : 
                  (N13243)? mem[168] : 
                  (N13245)? mem[170] : 
                  (N13247)? mem[172] : 
                  (N13249)? mem[174] : 
                  (N13251)? mem[176] : 
                  (N13253)? mem[178] : 
                  (N13255)? mem[180] : 
                  (N13257)? mem[182] : 
                  (N13259)? mem[184] : 
                  (N13261)? mem[186] : 
                  (N13263)? mem[188] : 
                  (N13265)? mem[190] : 
                  (N13267)? mem[192] : 
                  (N13269)? mem[194] : 
                  (N13271)? mem[196] : 
                  (N13273)? mem[198] : 
                  (N13275)? mem[200] : 
                  (N13277)? mem[202] : 
                  (N13279)? mem[204] : 
                  (N13281)? mem[206] : 
                  (N13283)? mem[208] : 
                  (N13285)? mem[210] : 
                  (N13287)? mem[212] : 
                  (N13289)? mem[214] : 
                  (N13291)? mem[216] : 
                  (N13293)? mem[218] : 
                  (N13295)? mem[220] : 
                  (N13297)? mem[222] : 
                  (N13299)? mem[224] : 
                  (N13301)? mem[226] : 
                  (N13303)? mem[228] : 
                  (N13305)? mem[230] : 
                  (N13307)? mem[232] : 
                  (N13309)? mem[234] : 
                  (N13311)? mem[236] : 
                  (N13313)? mem[238] : 
                  (N13315)? mem[240] : 
                  (N13317)? mem[242] : 
                  (N13319)? mem[244] : 
                  (N13321)? mem[246] : 
                  (N13323)? mem[248] : 
                  (N13325)? mem[250] : 
                  (N13327)? mem[252] : 
                  (N13329)? mem[254] : 
                  (N13331)? mem[256] : 
                  (N13333)? mem[258] : 
                  (N13335)? mem[260] : 
                  (N13337)? mem[262] : 
                  (N13339)? mem[264] : 
                  (N13341)? mem[266] : 
                  (N13343)? mem[268] : 
                  (N13345)? mem[270] : 
                  (N13347)? mem[272] : 
                  (N13349)? mem[274] : 
                  (N13351)? mem[276] : 
                  (N13353)? mem[278] : 
                  (N13355)? mem[280] : 
                  (N13357)? mem[282] : 
                  (N13359)? mem[284] : 
                  (N13361)? mem[286] : 
                  (N13363)? mem[288] : 
                  (N13365)? mem[290] : 
                  (N13367)? mem[292] : 
                  (N13369)? mem[294] : 
                  (N13371)? mem[296] : 
                  (N13373)? mem[298] : 
                  (N13375)? mem[300] : 
                  (N13377)? mem[302] : 
                  (N13379)? mem[304] : 
                  (N13381)? mem[306] : 
                  (N13383)? mem[308] : 
                  (N13385)? mem[310] : 
                  (N13387)? mem[312] : 
                  (N13389)? mem[314] : 
                  (N13391)? mem[316] : 
                  (N13393)? mem[318] : 
                  (N13395)? mem[320] : 
                  (N13397)? mem[322] : 
                  (N13399)? mem[324] : 
                  (N13401)? mem[326] : 
                  (N13403)? mem[328] : 
                  (N13405)? mem[330] : 
                  (N13407)? mem[332] : 
                  (N13409)? mem[334] : 
                  (N13411)? mem[336] : 
                  (N13413)? mem[338] : 
                  (N13415)? mem[340] : 
                  (N13417)? mem[342] : 
                  (N13419)? mem[344] : 
                  (N13421)? mem[346] : 
                  (N13423)? mem[348] : 
                  (N13425)? mem[350] : 
                  (N13427)? mem[352] : 
                  (N13429)? mem[354] : 
                  (N13431)? mem[356] : 
                  (N13433)? mem[358] : 
                  (N13435)? mem[360] : 
                  (N13437)? mem[362] : 
                  (N13439)? mem[364] : 
                  (N13441)? mem[366] : 
                  (N13443)? mem[368] : 
                  (N13445)? mem[370] : 
                  (N13447)? mem[372] : 
                  (N13449)? mem[374] : 
                  (N13451)? mem[376] : 
                  (N13453)? mem[378] : 
                  (N13455)? mem[380] : 
                  (N13457)? mem[382] : 
                  (N13459)? mem[384] : 
                  (N13460)? mem[386] : 
                  (N13461)? mem[388] : 
                  (N13462)? mem[390] : 
                  (N13463)? mem[392] : 
                  (N13464)? mem[394] : 
                  (N13465)? mem[396] : 
                  (N13466)? mem[398] : 
                  (N13467)? mem[400] : 
                  (N13468)? mem[402] : 
                  (N13469)? mem[404] : 
                  (N13470)? mem[406] : 
                  (N13471)? mem[408] : 
                  (N13472)? mem[410] : 
                  (N13473)? mem[412] : 
                  (N13474)? mem[414] : 
                  (N13475)? mem[416] : 
                  (N13476)? mem[418] : 
                  (N13477)? mem[420] : 
                  (N13478)? mem[422] : 
                  (N13479)? mem[424] : 
                  (N13480)? mem[426] : 
                  (N13481)? mem[428] : 
                  (N13482)? mem[430] : 
                  (N13483)? mem[432] : 
                  (N13484)? mem[434] : 
                  (N13485)? mem[436] : 
                  (N13486)? mem[438] : 
                  (N13487)? mem[440] : 
                  (N13488)? mem[442] : 
                  (N13489)? mem[444] : 
                  (N13490)? mem[446] : 
                  (N13491)? mem[448] : 
                  (N13492)? mem[450] : 
                  (N13493)? mem[452] : 
                  (N13494)? mem[454] : 
                  (N13495)? mem[456] : 
                  (N13496)? mem[458] : 
                  (N13497)? mem[460] : 
                  (N13498)? mem[462] : 
                  (N13499)? mem[464] : 
                  (N13500)? mem[466] : 
                  (N13501)? mem[468] : 
                  (N13502)? mem[470] : 
                  (N13503)? mem[472] : 
                  (N13504)? mem[474] : 
                  (N13505)? mem[476] : 
                  (N13506)? mem[478] : 
                  (N13507)? mem[480] : 
                  (N13508)? mem[482] : 
                  (N13509)? mem[484] : 
                  (N13510)? mem[486] : 
                  (N13511)? mem[488] : 
                  (N13512)? mem[490] : 
                  (N13513)? mem[492] : 
                  (N13514)? mem[494] : 
                  (N13515)? mem[496] : 
                  (N13516)? mem[498] : 
                  (N13517)? mem[500] : 
                  (N13518)? mem[502] : 
                  (N13519)? mem[504] : 
                  (N13520)? mem[506] : 
                  (N13521)? mem[508] : 
                  (N13522)? mem[510] : 
                  (N13076)? mem[512] : 
                  (N13078)? mem[514] : 
                  (N13080)? mem[516] : 
                  (N13082)? mem[518] : 
                  (N13084)? mem[520] : 
                  (N13086)? mem[522] : 
                  (N13088)? mem[524] : 
                  (N13090)? mem[526] : 
                  (N13092)? mem[528] : 
                  (N13094)? mem[530] : 
                  (N13096)? mem[532] : 
                  (N13098)? mem[534] : 
                  (N13100)? mem[536] : 
                  (N13102)? mem[538] : 
                  (N13104)? mem[540] : 
                  (N13106)? mem[542] : 
                  (N13108)? mem[544] : 
                  (N13110)? mem[546] : 
                  (N13112)? mem[548] : 
                  (N13114)? mem[550] : 
                  (N13116)? mem[552] : 
                  (N13118)? mem[554] : 
                  (N13120)? mem[556] : 
                  (N13122)? mem[558] : 
                  (N13124)? mem[560] : 
                  (N13126)? mem[562] : 
                  (N13128)? mem[564] : 
                  (N13130)? mem[566] : 
                  (N13132)? mem[568] : 
                  (N13134)? mem[570] : 
                  (N13136)? mem[572] : 
                  (N13138)? mem[574] : 
                  (N13140)? mem[576] : 
                  (N13142)? mem[578] : 
                  (N13144)? mem[580] : 
                  (N13146)? mem[582] : 
                  (N13148)? mem[584] : 
                  (N13150)? mem[586] : 
                  (N13152)? mem[588] : 
                  (N13154)? mem[590] : 
                  (N13156)? mem[592] : 
                  (N13158)? mem[594] : 
                  (N13160)? mem[596] : 
                  (N13162)? mem[598] : 
                  (N13164)? mem[600] : 
                  (N13166)? mem[602] : 
                  (N13168)? mem[604] : 
                  (N13170)? mem[606] : 
                  (N13172)? mem[608] : 
                  (N13174)? mem[610] : 
                  (N13176)? mem[612] : 
                  (N13178)? mem[614] : 
                  (N13180)? mem[616] : 
                  (N13182)? mem[618] : 
                  (N13184)? mem[620] : 
                  (N13186)? mem[622] : 
                  (N13188)? mem[624] : 
                  (N13190)? mem[626] : 
                  (N13192)? mem[628] : 
                  (N13194)? mem[630] : 
                  (N13196)? mem[632] : 
                  (N13198)? mem[634] : 
                  (N13200)? mem[636] : 
                  (N13202)? mem[638] : 
                  (N13204)? mem[640] : 
                  (N13206)? mem[642] : 
                  (N13208)? mem[644] : 
                  (N13210)? mem[646] : 
                  (N13212)? mem[648] : 
                  (N13214)? mem[650] : 
                  (N13216)? mem[652] : 
                  (N13218)? mem[654] : 
                  (N13220)? mem[656] : 
                  (N13222)? mem[658] : 
                  (N13224)? mem[660] : 
                  (N13226)? mem[662] : 
                  (N13228)? mem[664] : 
                  (N13230)? mem[666] : 
                  (N13232)? mem[668] : 
                  (N13234)? mem[670] : 
                  (N13236)? mem[672] : 
                  (N13238)? mem[674] : 
                  (N13240)? mem[676] : 
                  (N13242)? mem[678] : 
                  (N13244)? mem[680] : 
                  (N13246)? mem[682] : 
                  (N13248)? mem[684] : 
                  (N13250)? mem[686] : 
                  (N13252)? mem[688] : 
                  (N13254)? mem[690] : 
                  (N13256)? mem[692] : 
                  (N13258)? mem[694] : 
                  (N13260)? mem[696] : 
                  (N13262)? mem[698] : 
                  (N13264)? mem[700] : 
                  (N13266)? mem[702] : 
                  (N13268)? mem[704] : 
                  (N13270)? mem[706] : 
                  (N13272)? mem[708] : 
                  (N13274)? mem[710] : 
                  (N13276)? mem[712] : 
                  (N13278)? mem[714] : 
                  (N13280)? mem[716] : 
                  (N13282)? mem[718] : 
                  (N13284)? mem[720] : 
                  (N13286)? mem[722] : 
                  (N13288)? mem[724] : 
                  (N13290)? mem[726] : 
                  (N13292)? mem[728] : 
                  (N13294)? mem[730] : 
                  (N13296)? mem[732] : 
                  (N13298)? mem[734] : 
                  (N13300)? mem[736] : 
                  (N13302)? mem[738] : 
                  (N13304)? mem[740] : 
                  (N13306)? mem[742] : 
                  (N13308)? mem[744] : 
                  (N13310)? mem[746] : 
                  (N13312)? mem[748] : 
                  (N13314)? mem[750] : 
                  (N13316)? mem[752] : 
                  (N13318)? mem[754] : 
                  (N13320)? mem[756] : 
                  (N13322)? mem[758] : 
                  (N13324)? mem[760] : 
                  (N13326)? mem[762] : 
                  (N13328)? mem[764] : 
                  (N13330)? mem[766] : 
                  (N13332)? mem[768] : 
                  (N13334)? mem[770] : 
                  (N13336)? mem[772] : 
                  (N13338)? mem[774] : 
                  (N13340)? mem[776] : 
                  (N13342)? mem[778] : 
                  (N13344)? mem[780] : 
                  (N13346)? mem[782] : 
                  (N13348)? mem[784] : 
                  (N13350)? mem[786] : 
                  (N13352)? mem[788] : 
                  (N13354)? mem[790] : 
                  (N13356)? mem[792] : 
                  (N13358)? mem[794] : 
                  (N13360)? mem[796] : 
                  (N13362)? mem[798] : 
                  (N13364)? mem[800] : 
                  (N13366)? mem[802] : 
                  (N13368)? mem[804] : 
                  (N13370)? mem[806] : 
                  (N13372)? mem[808] : 
                  (N13374)? mem[810] : 
                  (N13376)? mem[812] : 
                  (N13378)? mem[814] : 
                  (N13380)? mem[816] : 
                  (N13382)? mem[818] : 
                  (N13384)? mem[820] : 
                  (N13386)? mem[822] : 
                  (N13388)? mem[824] : 
                  (N13390)? mem[826] : 
                  (N13392)? mem[828] : 
                  (N13394)? mem[830] : 
                  (N13396)? mem[832] : 
                  (N13398)? mem[834] : 
                  (N13400)? mem[836] : 
                  (N13402)? mem[838] : 
                  (N13404)? mem[840] : 
                  (N13406)? mem[842] : 
                  (N13408)? mem[844] : 
                  (N13410)? mem[846] : 
                  (N13412)? mem[848] : 
                  (N13414)? mem[850] : 
                  (N13416)? mem[852] : 
                  (N13418)? mem[854] : 
                  (N13420)? mem[856] : 
                  (N13422)? mem[858] : 
                  (N13424)? mem[860] : 
                  (N13426)? mem[862] : 
                  (N13428)? mem[864] : 
                  (N13430)? mem[866] : 
                  (N13432)? mem[868] : 
                  (N13434)? mem[870] : 
                  (N13436)? mem[872] : 
                  (N13438)? mem[874] : 
                  (N13440)? mem[876] : 
                  (N13442)? mem[878] : 
                  (N13444)? mem[880] : 
                  (N13446)? mem[882] : 
                  (N13448)? mem[884] : 
                  (N13450)? mem[886] : 
                  (N13452)? mem[888] : 
                  (N13454)? mem[890] : 
                  (N13456)? mem[892] : 
                  (N13458)? mem[894] : 
                  (N10992)? mem[896] : 
                  (N10994)? mem[898] : 
                  (N10996)? mem[900] : 
                  (N10998)? mem[902] : 
                  (N11000)? mem[904] : 
                  (N11002)? mem[906] : 
                  (N11004)? mem[908] : 
                  (N11006)? mem[910] : 
                  (N11008)? mem[912] : 
                  (N11010)? mem[914] : 
                  (N11012)? mem[916] : 
                  (N11014)? mem[918] : 
                  (N11016)? mem[920] : 
                  (N11018)? mem[922] : 
                  (N11020)? mem[924] : 
                  (N11022)? mem[926] : 
                  (N11024)? mem[928] : 
                  (N11026)? mem[930] : 
                  (N11028)? mem[932] : 
                  (N11030)? mem[934] : 
                  (N11032)? mem[936] : 
                  (N11034)? mem[938] : 
                  (N11036)? mem[940] : 
                  (N11038)? mem[942] : 
                  (N11040)? mem[944] : 
                  (N11042)? mem[946] : 
                  (N11044)? mem[948] : 
                  (N11046)? mem[950] : 
                  (N11048)? mem[952] : 
                  (N11050)? mem[954] : 
                  (N11052)? mem[956] : 
                  (N11054)? mem[958] : 
                  (N12049)? mem[960] : 
                  (N12051)? mem[962] : 
                  (N12053)? mem[964] : 
                  (N12055)? mem[966] : 
                  (N12057)? mem[968] : 
                  (N12059)? mem[970] : 
                  (N12061)? mem[972] : 
                  (N12063)? mem[974] : 
                  (N12065)? mem[976] : 
                  (N12067)? mem[978] : 
                  (N12069)? mem[980] : 
                  (N12071)? mem[982] : 
                  (N12073)? mem[984] : 
                  (N12075)? mem[986] : 
                  (N12077)? mem[988] : 
                  (N12079)? mem[990] : 
                  (N12081)? mem[992] : 
                  (N12083)? mem[994] : 
                  (N12085)? mem[996] : 
                  (N12087)? mem[998] : 
                  (N12089)? mem[1000] : 
                  (N12091)? mem[1002] : 
                  (N12093)? mem[1004] : 
                  (N12095)? mem[1006] : 
                  (N12097)? mem[1008] : 
                  (N12099)? mem[1010] : 
                  (N12101)? mem[1012] : 
                  (N12103)? mem[1014] : 
                  (N12105)? mem[1016] : 
                  (N12107)? mem[1018] : 
                  (N12109)? mem[1020] : 
                  (N12111)? mem[1022] : 1'b0;
  assign N14741 = (N14293)? mem[1] : 
                  (N14295)? mem[3] : 
                  (N14297)? mem[5] : 
                  (N14299)? mem[7] : 
                  (N14301)? mem[9] : 
                  (N14303)? mem[11] : 
                  (N14305)? mem[13] : 
                  (N14307)? mem[15] : 
                  (N14309)? mem[17] : 
                  (N14311)? mem[19] : 
                  (N14313)? mem[21] : 
                  (N14315)? mem[23] : 
                  (N14317)? mem[25] : 
                  (N14319)? mem[27] : 
                  (N14321)? mem[29] : 
                  (N14323)? mem[31] : 
                  (N14325)? mem[33] : 
                  (N14327)? mem[35] : 
                  (N14329)? mem[37] : 
                  (N14331)? mem[39] : 
                  (N14333)? mem[41] : 
                  (N14335)? mem[43] : 
                  (N14337)? mem[45] : 
                  (N14339)? mem[47] : 
                  (N14341)? mem[49] : 
                  (N14343)? mem[51] : 
                  (N14345)? mem[53] : 
                  (N14347)? mem[55] : 
                  (N14349)? mem[57] : 
                  (N14351)? mem[59] : 
                  (N14353)? mem[61] : 
                  (N14355)? mem[63] : 
                  (N14357)? mem[65] : 
                  (N14359)? mem[67] : 
                  (N14361)? mem[69] : 
                  (N14363)? mem[71] : 
                  (N14365)? mem[73] : 
                  (N14367)? mem[75] : 
                  (N14369)? mem[77] : 
                  (N14371)? mem[79] : 
                  (N14373)? mem[81] : 
                  (N14375)? mem[83] : 
                  (N14377)? mem[85] : 
                  (N14379)? mem[87] : 
                  (N14381)? mem[89] : 
                  (N14383)? mem[91] : 
                  (N14385)? mem[93] : 
                  (N14387)? mem[95] : 
                  (N14389)? mem[97] : 
                  (N14391)? mem[99] : 
                  (N14393)? mem[101] : 
                  (N14395)? mem[103] : 
                  (N14397)? mem[105] : 
                  (N14399)? mem[107] : 
                  (N14401)? mem[109] : 
                  (N14403)? mem[111] : 
                  (N14405)? mem[113] : 
                  (N14407)? mem[115] : 
                  (N14409)? mem[117] : 
                  (N14411)? mem[119] : 
                  (N14413)? mem[121] : 
                  (N14415)? mem[123] : 
                  (N14417)? mem[125] : 
                  (N14419)? mem[127] : 
                  (N14421)? mem[129] : 
                  (N14423)? mem[131] : 
                  (N14425)? mem[133] : 
                  (N14427)? mem[135] : 
                  (N14429)? mem[137] : 
                  (N14431)? mem[139] : 
                  (N14433)? mem[141] : 
                  (N14435)? mem[143] : 
                  (N14437)? mem[145] : 
                  (N14439)? mem[147] : 
                  (N14441)? mem[149] : 
                  (N14443)? mem[151] : 
                  (N14445)? mem[153] : 
                  (N14447)? mem[155] : 
                  (N14449)? mem[157] : 
                  (N14451)? mem[159] : 
                  (N14453)? mem[161] : 
                  (N14455)? mem[163] : 
                  (N14457)? mem[165] : 
                  (N14459)? mem[167] : 
                  (N14461)? mem[169] : 
                  (N14463)? mem[171] : 
                  (N14465)? mem[173] : 
                  (N14467)? mem[175] : 
                  (N14469)? mem[177] : 
                  (N14471)? mem[179] : 
                  (N14473)? mem[181] : 
                  (N14475)? mem[183] : 
                  (N14477)? mem[185] : 
                  (N14479)? mem[187] : 
                  (N14481)? mem[189] : 
                  (N14483)? mem[191] : 
                  (N14485)? mem[193] : 
                  (N14487)? mem[195] : 
                  (N14489)? mem[197] : 
                  (N14491)? mem[199] : 
                  (N14493)? mem[201] : 
                  (N14495)? mem[203] : 
                  (N14497)? mem[205] : 
                  (N14499)? mem[207] : 
                  (N14501)? mem[209] : 
                  (N14503)? mem[211] : 
                  (N14505)? mem[213] : 
                  (N14507)? mem[215] : 
                  (N14509)? mem[217] : 
                  (N14511)? mem[219] : 
                  (N14513)? mem[221] : 
                  (N14515)? mem[223] : 
                  (N14517)? mem[225] : 
                  (N14519)? mem[227] : 
                  (N14521)? mem[229] : 
                  (N14523)? mem[231] : 
                  (N14525)? mem[233] : 
                  (N14527)? mem[235] : 
                  (N14529)? mem[237] : 
                  (N14531)? mem[239] : 
                  (N14533)? mem[241] : 
                  (N14535)? mem[243] : 
                  (N14537)? mem[245] : 
                  (N14539)? mem[247] : 
                  (N14541)? mem[249] : 
                  (N14543)? mem[251] : 
                  (N14545)? mem[253] : 
                  (N14547)? mem[255] : 
                  (N14549)? mem[257] : 
                  (N14551)? mem[259] : 
                  (N14553)? mem[261] : 
                  (N14555)? mem[263] : 
                  (N14557)? mem[265] : 
                  (N14559)? mem[267] : 
                  (N14561)? mem[269] : 
                  (N14563)? mem[271] : 
                  (N14565)? mem[273] : 
                  (N14567)? mem[275] : 
                  (N14569)? mem[277] : 
                  (N14571)? mem[279] : 
                  (N14573)? mem[281] : 
                  (N14575)? mem[283] : 
                  (N14577)? mem[285] : 
                  (N14579)? mem[287] : 
                  (N14581)? mem[289] : 
                  (N14583)? mem[291] : 
                  (N14585)? mem[293] : 
                  (N14587)? mem[295] : 
                  (N14589)? mem[297] : 
                  (N14591)? mem[299] : 
                  (N14593)? mem[301] : 
                  (N14595)? mem[303] : 
                  (N14597)? mem[305] : 
                  (N14599)? mem[307] : 
                  (N14601)? mem[309] : 
                  (N14603)? mem[311] : 
                  (N14605)? mem[313] : 
                  (N14607)? mem[315] : 
                  (N14609)? mem[317] : 
                  (N14611)? mem[319] : 
                  (N14613)? mem[321] : 
                  (N14615)? mem[323] : 
                  (N14617)? mem[325] : 
                  (N14619)? mem[327] : 
                  (N14621)? mem[329] : 
                  (N14623)? mem[331] : 
                  (N14625)? mem[333] : 
                  (N14627)? mem[335] : 
                  (N14629)? mem[337] : 
                  (N14631)? mem[339] : 
                  (N14633)? mem[341] : 
                  (N14635)? mem[343] : 
                  (N14637)? mem[345] : 
                  (N14639)? mem[347] : 
                  (N14641)? mem[349] : 
                  (N14643)? mem[351] : 
                  (N14645)? mem[353] : 
                  (N14647)? mem[355] : 
                  (N14649)? mem[357] : 
                  (N14651)? mem[359] : 
                  (N14653)? mem[361] : 
                  (N14655)? mem[363] : 
                  (N14657)? mem[365] : 
                  (N14659)? mem[367] : 
                  (N14661)? mem[369] : 
                  (N14663)? mem[371] : 
                  (N14665)? mem[373] : 
                  (N14667)? mem[375] : 
                  (N14669)? mem[377] : 
                  (N14671)? mem[379] : 
                  (N14673)? mem[381] : 
                  (N14675)? mem[383] : 
                  (N14677)? mem[385] : 
                  (N14678)? mem[387] : 
                  (N14679)? mem[389] : 
                  (N14680)? mem[391] : 
                  (N14681)? mem[393] : 
                  (N14682)? mem[395] : 
                  (N14683)? mem[397] : 
                  (N14684)? mem[399] : 
                  (N14685)? mem[401] : 
                  (N14686)? mem[403] : 
                  (N14687)? mem[405] : 
                  (N14688)? mem[407] : 
                  (N14689)? mem[409] : 
                  (N14690)? mem[411] : 
                  (N14691)? mem[413] : 
                  (N14692)? mem[415] : 
                  (N14693)? mem[417] : 
                  (N14694)? mem[419] : 
                  (N14695)? mem[421] : 
                  (N14696)? mem[423] : 
                  (N14697)? mem[425] : 
                  (N14698)? mem[427] : 
                  (N14699)? mem[429] : 
                  (N14700)? mem[431] : 
                  (N14701)? mem[433] : 
                  (N14702)? mem[435] : 
                  (N14703)? mem[437] : 
                  (N14704)? mem[439] : 
                  (N14705)? mem[441] : 
                  (N14706)? mem[443] : 
                  (N14707)? mem[445] : 
                  (N14708)? mem[447] : 
                  (N14709)? mem[449] : 
                  (N14710)? mem[451] : 
                  (N14711)? mem[453] : 
                  (N14712)? mem[455] : 
                  (N14713)? mem[457] : 
                  (N14714)? mem[459] : 
                  (N14715)? mem[461] : 
                  (N14716)? mem[463] : 
                  (N14717)? mem[465] : 
                  (N14718)? mem[467] : 
                  (N14719)? mem[469] : 
                  (N14720)? mem[471] : 
                  (N14721)? mem[473] : 
                  (N14722)? mem[475] : 
                  (N14723)? mem[477] : 
                  (N14724)? mem[479] : 
                  (N14725)? mem[481] : 
                  (N14726)? mem[483] : 
                  (N14727)? mem[485] : 
                  (N14728)? mem[487] : 
                  (N14729)? mem[489] : 
                  (N14730)? mem[491] : 
                  (N14731)? mem[493] : 
                  (N14732)? mem[495] : 
                  (N14733)? mem[497] : 
                  (N14734)? mem[499] : 
                  (N14735)? mem[501] : 
                  (N14736)? mem[503] : 
                  (N14737)? mem[505] : 
                  (N14738)? mem[507] : 
                  (N14739)? mem[509] : 
                  (N14740)? mem[511] : 
                  (N14294)? mem[513] : 
                  (N14296)? mem[515] : 
                  (N14298)? mem[517] : 
                  (N14300)? mem[519] : 
                  (N14302)? mem[521] : 
                  (N14304)? mem[523] : 
                  (N14306)? mem[525] : 
                  (N14308)? mem[527] : 
                  (N14310)? mem[529] : 
                  (N14312)? mem[531] : 
                  (N14314)? mem[533] : 
                  (N14316)? mem[535] : 
                  (N14318)? mem[537] : 
                  (N14320)? mem[539] : 
                  (N14322)? mem[541] : 
                  (N14324)? mem[543] : 
                  (N14326)? mem[545] : 
                  (N14328)? mem[547] : 
                  (N14330)? mem[549] : 
                  (N14332)? mem[551] : 
                  (N14334)? mem[553] : 
                  (N14336)? mem[555] : 
                  (N14338)? mem[557] : 
                  (N14340)? mem[559] : 
                  (N14342)? mem[561] : 
                  (N14344)? mem[563] : 
                  (N14346)? mem[565] : 
                  (N14348)? mem[567] : 
                  (N14350)? mem[569] : 
                  (N14352)? mem[571] : 
                  (N14354)? mem[573] : 
                  (N14356)? mem[575] : 
                  (N14358)? mem[577] : 
                  (N14360)? mem[579] : 
                  (N14362)? mem[581] : 
                  (N14364)? mem[583] : 
                  (N14366)? mem[585] : 
                  (N14368)? mem[587] : 
                  (N14370)? mem[589] : 
                  (N14372)? mem[591] : 
                  (N14374)? mem[593] : 
                  (N14376)? mem[595] : 
                  (N14378)? mem[597] : 
                  (N14380)? mem[599] : 
                  (N14382)? mem[601] : 
                  (N14384)? mem[603] : 
                  (N14386)? mem[605] : 
                  (N14388)? mem[607] : 
                  (N14390)? mem[609] : 
                  (N14392)? mem[611] : 
                  (N14394)? mem[613] : 
                  (N14396)? mem[615] : 
                  (N14398)? mem[617] : 
                  (N14400)? mem[619] : 
                  (N14402)? mem[621] : 
                  (N14404)? mem[623] : 
                  (N14406)? mem[625] : 
                  (N14408)? mem[627] : 
                  (N14410)? mem[629] : 
                  (N14412)? mem[631] : 
                  (N14414)? mem[633] : 
                  (N14416)? mem[635] : 
                  (N14418)? mem[637] : 
                  (N14420)? mem[639] : 
                  (N14422)? mem[641] : 
                  (N14424)? mem[643] : 
                  (N14426)? mem[645] : 
                  (N14428)? mem[647] : 
                  (N14430)? mem[649] : 
                  (N14432)? mem[651] : 
                  (N14434)? mem[653] : 
                  (N14436)? mem[655] : 
                  (N14438)? mem[657] : 
                  (N14440)? mem[659] : 
                  (N14442)? mem[661] : 
                  (N14444)? mem[663] : 
                  (N14446)? mem[665] : 
                  (N14448)? mem[667] : 
                  (N14450)? mem[669] : 
                  (N14452)? mem[671] : 
                  (N14454)? mem[673] : 
                  (N14456)? mem[675] : 
                  (N14458)? mem[677] : 
                  (N14460)? mem[679] : 
                  (N14462)? mem[681] : 
                  (N14464)? mem[683] : 
                  (N14466)? mem[685] : 
                  (N14468)? mem[687] : 
                  (N14470)? mem[689] : 
                  (N14472)? mem[691] : 
                  (N14474)? mem[693] : 
                  (N14476)? mem[695] : 
                  (N14478)? mem[697] : 
                  (N14480)? mem[699] : 
                  (N14482)? mem[701] : 
                  (N14484)? mem[703] : 
                  (N14486)? mem[705] : 
                  (N14488)? mem[707] : 
                  (N14490)? mem[709] : 
                  (N14492)? mem[711] : 
                  (N14494)? mem[713] : 
                  (N14496)? mem[715] : 
                  (N14498)? mem[717] : 
                  (N14500)? mem[719] : 
                  (N14502)? mem[721] : 
                  (N14504)? mem[723] : 
                  (N14506)? mem[725] : 
                  (N14508)? mem[727] : 
                  (N14510)? mem[729] : 
                  (N14512)? mem[731] : 
                  (N14514)? mem[733] : 
                  (N14516)? mem[735] : 
                  (N14518)? mem[737] : 
                  (N14520)? mem[739] : 
                  (N14522)? mem[741] : 
                  (N14524)? mem[743] : 
                  (N14526)? mem[745] : 
                  (N14528)? mem[747] : 
                  (N14530)? mem[749] : 
                  (N14532)? mem[751] : 
                  (N14534)? mem[753] : 
                  (N14536)? mem[755] : 
                  (N14538)? mem[757] : 
                  (N14540)? mem[759] : 
                  (N14542)? mem[761] : 
                  (N14544)? mem[763] : 
                  (N14546)? mem[765] : 
                  (N14548)? mem[767] : 
                  (N14550)? mem[769] : 
                  (N14552)? mem[771] : 
                  (N14554)? mem[773] : 
                  (N14556)? mem[775] : 
                  (N14558)? mem[777] : 
                  (N14560)? mem[779] : 
                  (N14562)? mem[781] : 
                  (N14564)? mem[783] : 
                  (N14566)? mem[785] : 
                  (N14568)? mem[787] : 
                  (N14570)? mem[789] : 
                  (N14572)? mem[791] : 
                  (N14574)? mem[793] : 
                  (N14576)? mem[795] : 
                  (N14578)? mem[797] : 
                  (N14580)? mem[799] : 
                  (N14582)? mem[801] : 
                  (N14584)? mem[803] : 
                  (N14586)? mem[805] : 
                  (N14588)? mem[807] : 
                  (N14590)? mem[809] : 
                  (N14592)? mem[811] : 
                  (N14594)? mem[813] : 
                  (N14596)? mem[815] : 
                  (N14598)? mem[817] : 
                  (N14600)? mem[819] : 
                  (N14602)? mem[821] : 
                  (N14604)? mem[823] : 
                  (N14606)? mem[825] : 
                  (N14608)? mem[827] : 
                  (N14610)? mem[829] : 
                  (N14612)? mem[831] : 
                  (N14614)? mem[833] : 
                  (N14616)? mem[835] : 
                  (N14618)? mem[837] : 
                  (N14620)? mem[839] : 
                  (N14622)? mem[841] : 
                  (N14624)? mem[843] : 
                  (N14626)? mem[845] : 
                  (N14628)? mem[847] : 
                  (N14630)? mem[849] : 
                  (N14632)? mem[851] : 
                  (N14634)? mem[853] : 
                  (N14636)? mem[855] : 
                  (N14638)? mem[857] : 
                  (N14640)? mem[859] : 
                  (N14642)? mem[861] : 
                  (N14644)? mem[863] : 
                  (N14646)? mem[865] : 
                  (N14648)? mem[867] : 
                  (N14650)? mem[869] : 
                  (N14652)? mem[871] : 
                  (N14654)? mem[873] : 
                  (N14656)? mem[875] : 
                  (N14658)? mem[877] : 
                  (N14660)? mem[879] : 
                  (N14662)? mem[881] : 
                  (N14664)? mem[883] : 
                  (N14666)? mem[885] : 
                  (N14668)? mem[887] : 
                  (N14670)? mem[889] : 
                  (N14672)? mem[891] : 
                  (N14674)? mem[893] : 
                  (N14676)? mem[895] : 
                  (N11985)? mem[897] : 
                  (N11987)? mem[899] : 
                  (N11989)? mem[901] : 
                  (N11991)? mem[903] : 
                  (N11993)? mem[905] : 
                  (N11995)? mem[907] : 
                  (N11997)? mem[909] : 
                  (N11999)? mem[911] : 
                  (N12001)? mem[913] : 
                  (N12003)? mem[915] : 
                  (N12005)? mem[917] : 
                  (N12007)? mem[919] : 
                  (N12009)? mem[921] : 
                  (N12011)? mem[923] : 
                  (N12013)? mem[925] : 
                  (N12015)? mem[927] : 
                  (N12017)? mem[929] : 
                  (N12019)? mem[931] : 
                  (N12021)? mem[933] : 
                  (N12023)? mem[935] : 
                  (N12025)? mem[937] : 
                  (N12027)? mem[939] : 
                  (N12029)? mem[941] : 
                  (N12031)? mem[943] : 
                  (N12033)? mem[945] : 
                  (N12035)? mem[947] : 
                  (N12037)? mem[949] : 
                  (N12039)? mem[951] : 
                  (N12041)? mem[953] : 
                  (N12043)? mem[955] : 
                  (N12045)? mem[957] : 
                  (N12047)? mem[959] : 
                  (N12049)? mem[961] : 
                  (N12051)? mem[963] : 
                  (N12053)? mem[965] : 
                  (N12055)? mem[967] : 
                  (N12057)? mem[969] : 
                  (N12059)? mem[971] : 
                  (N12061)? mem[973] : 
                  (N12063)? mem[975] : 
                  (N12065)? mem[977] : 
                  (N12067)? mem[979] : 
                  (N12069)? mem[981] : 
                  (N12071)? mem[983] : 
                  (N12073)? mem[985] : 
                  (N12075)? mem[987] : 
                  (N12077)? mem[989] : 
                  (N12079)? mem[991] : 
                  (N12081)? mem[993] : 
                  (N12083)? mem[995] : 
                  (N12085)? mem[997] : 
                  (N12087)? mem[999] : 
                  (N12089)? mem[1001] : 
                  (N12091)? mem[1003] : 
                  (N12093)? mem[1005] : 
                  (N12095)? mem[1007] : 
                  (N12097)? mem[1009] : 
                  (N12099)? mem[1011] : 
                  (N12101)? mem[1013] : 
                  (N12103)? mem[1015] : 
                  (N12105)? mem[1017] : 
                  (N12107)? mem[1019] : 
                  (N12109)? mem[1021] : 
                  (N12111)? mem[1023] : 1'b0;
  assign N15446 = (N14998)? mem[0] : 
                  (N15000)? mem[2] : 
                  (N15002)? mem[4] : 
                  (N15004)? mem[6] : 
                  (N15006)? mem[8] : 
                  (N15008)? mem[10] : 
                  (N15010)? mem[12] : 
                  (N15012)? mem[14] : 
                  (N15014)? mem[16] : 
                  (N15016)? mem[18] : 
                  (N15018)? mem[20] : 
                  (N15020)? mem[22] : 
                  (N15022)? mem[24] : 
                  (N15024)? mem[26] : 
                  (N15026)? mem[28] : 
                  (N15028)? mem[30] : 
                  (N15030)? mem[32] : 
                  (N15032)? mem[34] : 
                  (N15034)? mem[36] : 
                  (N15036)? mem[38] : 
                  (N15038)? mem[40] : 
                  (N15040)? mem[42] : 
                  (N15042)? mem[44] : 
                  (N15044)? mem[46] : 
                  (N15046)? mem[48] : 
                  (N15048)? mem[50] : 
                  (N15050)? mem[52] : 
                  (N15052)? mem[54] : 
                  (N15054)? mem[56] : 
                  (N15056)? mem[58] : 
                  (N15058)? mem[60] : 
                  (N15060)? mem[62] : 
                  (N15062)? mem[64] : 
                  (N15064)? mem[66] : 
                  (N15066)? mem[68] : 
                  (N15068)? mem[70] : 
                  (N15070)? mem[72] : 
                  (N15072)? mem[74] : 
                  (N15074)? mem[76] : 
                  (N15076)? mem[78] : 
                  (N15078)? mem[80] : 
                  (N15080)? mem[82] : 
                  (N15082)? mem[84] : 
                  (N15084)? mem[86] : 
                  (N15086)? mem[88] : 
                  (N15088)? mem[90] : 
                  (N15090)? mem[92] : 
                  (N15092)? mem[94] : 
                  (N15094)? mem[96] : 
                  (N15096)? mem[98] : 
                  (N15098)? mem[100] : 
                  (N15100)? mem[102] : 
                  (N15102)? mem[104] : 
                  (N15104)? mem[106] : 
                  (N15106)? mem[108] : 
                  (N15108)? mem[110] : 
                  (N15110)? mem[112] : 
                  (N15112)? mem[114] : 
                  (N15114)? mem[116] : 
                  (N15116)? mem[118] : 
                  (N15118)? mem[120] : 
                  (N15120)? mem[122] : 
                  (N15122)? mem[124] : 
                  (N15124)? mem[126] : 
                  (N15126)? mem[128] : 
                  (N15128)? mem[130] : 
                  (N15130)? mem[132] : 
                  (N15132)? mem[134] : 
                  (N15134)? mem[136] : 
                  (N15136)? mem[138] : 
                  (N15138)? mem[140] : 
                  (N15140)? mem[142] : 
                  (N15142)? mem[144] : 
                  (N15144)? mem[146] : 
                  (N15146)? mem[148] : 
                  (N15148)? mem[150] : 
                  (N15150)? mem[152] : 
                  (N15152)? mem[154] : 
                  (N15154)? mem[156] : 
                  (N15156)? mem[158] : 
                  (N15158)? mem[160] : 
                  (N15160)? mem[162] : 
                  (N15162)? mem[164] : 
                  (N15164)? mem[166] : 
                  (N15166)? mem[168] : 
                  (N15168)? mem[170] : 
                  (N15170)? mem[172] : 
                  (N15172)? mem[174] : 
                  (N15174)? mem[176] : 
                  (N15176)? mem[178] : 
                  (N15178)? mem[180] : 
                  (N15180)? mem[182] : 
                  (N15182)? mem[184] : 
                  (N15184)? mem[186] : 
                  (N15186)? mem[188] : 
                  (N15188)? mem[190] : 
                  (N15190)? mem[192] : 
                  (N15192)? mem[194] : 
                  (N15194)? mem[196] : 
                  (N15196)? mem[198] : 
                  (N15198)? mem[200] : 
                  (N15200)? mem[202] : 
                  (N15202)? mem[204] : 
                  (N15204)? mem[206] : 
                  (N15206)? mem[208] : 
                  (N15208)? mem[210] : 
                  (N15210)? mem[212] : 
                  (N15212)? mem[214] : 
                  (N15214)? mem[216] : 
                  (N15216)? mem[218] : 
                  (N15218)? mem[220] : 
                  (N15220)? mem[222] : 
                  (N15222)? mem[224] : 
                  (N15224)? mem[226] : 
                  (N15226)? mem[228] : 
                  (N15228)? mem[230] : 
                  (N15230)? mem[232] : 
                  (N15232)? mem[234] : 
                  (N15234)? mem[236] : 
                  (N15236)? mem[238] : 
                  (N15238)? mem[240] : 
                  (N15240)? mem[242] : 
                  (N15242)? mem[244] : 
                  (N15244)? mem[246] : 
                  (N15246)? mem[248] : 
                  (N15248)? mem[250] : 
                  (N15250)? mem[252] : 
                  (N15252)? mem[254] : 
                  (N15254)? mem[256] : 
                  (N15256)? mem[258] : 
                  (N15258)? mem[260] : 
                  (N15260)? mem[262] : 
                  (N15262)? mem[264] : 
                  (N15264)? mem[266] : 
                  (N15266)? mem[268] : 
                  (N15268)? mem[270] : 
                  (N15270)? mem[272] : 
                  (N15272)? mem[274] : 
                  (N15274)? mem[276] : 
                  (N15276)? mem[278] : 
                  (N15278)? mem[280] : 
                  (N15280)? mem[282] : 
                  (N15282)? mem[284] : 
                  (N15284)? mem[286] : 
                  (N15286)? mem[288] : 
                  (N15288)? mem[290] : 
                  (N15290)? mem[292] : 
                  (N15292)? mem[294] : 
                  (N15294)? mem[296] : 
                  (N15296)? mem[298] : 
                  (N15298)? mem[300] : 
                  (N15300)? mem[302] : 
                  (N15302)? mem[304] : 
                  (N15304)? mem[306] : 
                  (N15306)? mem[308] : 
                  (N15308)? mem[310] : 
                  (N15310)? mem[312] : 
                  (N15312)? mem[314] : 
                  (N15314)? mem[316] : 
                  (N15316)? mem[318] : 
                  (N15318)? mem[320] : 
                  (N15320)? mem[322] : 
                  (N15322)? mem[324] : 
                  (N15324)? mem[326] : 
                  (N15326)? mem[328] : 
                  (N15328)? mem[330] : 
                  (N15330)? mem[332] : 
                  (N15332)? mem[334] : 
                  (N15334)? mem[336] : 
                  (N15336)? mem[338] : 
                  (N15338)? mem[340] : 
                  (N15340)? mem[342] : 
                  (N15342)? mem[344] : 
                  (N15344)? mem[346] : 
                  (N15346)? mem[348] : 
                  (N15348)? mem[350] : 
                  (N15350)? mem[352] : 
                  (N15352)? mem[354] : 
                  (N15354)? mem[356] : 
                  (N15356)? mem[358] : 
                  (N15358)? mem[360] : 
                  (N15360)? mem[362] : 
                  (N15362)? mem[364] : 
                  (N15364)? mem[366] : 
                  (N15366)? mem[368] : 
                  (N15368)? mem[370] : 
                  (N15370)? mem[372] : 
                  (N15372)? mem[374] : 
                  (N15374)? mem[376] : 
                  (N15376)? mem[378] : 
                  (N15378)? mem[380] : 
                  (N15380)? mem[382] : 
                  (N15382)? mem[384] : 
                  (N15383)? mem[386] : 
                  (N15384)? mem[388] : 
                  (N15385)? mem[390] : 
                  (N15386)? mem[392] : 
                  (N15387)? mem[394] : 
                  (N15388)? mem[396] : 
                  (N15389)? mem[398] : 
                  (N15390)? mem[400] : 
                  (N15391)? mem[402] : 
                  (N15392)? mem[404] : 
                  (N15393)? mem[406] : 
                  (N15394)? mem[408] : 
                  (N15395)? mem[410] : 
                  (N15396)? mem[412] : 
                  (N15397)? mem[414] : 
                  (N15398)? mem[416] : 
                  (N15399)? mem[418] : 
                  (N15400)? mem[420] : 
                  (N15401)? mem[422] : 
                  (N15402)? mem[424] : 
                  (N15403)? mem[426] : 
                  (N15404)? mem[428] : 
                  (N15405)? mem[430] : 
                  (N15406)? mem[432] : 
                  (N15407)? mem[434] : 
                  (N15408)? mem[436] : 
                  (N15409)? mem[438] : 
                  (N15410)? mem[440] : 
                  (N15411)? mem[442] : 
                  (N15412)? mem[444] : 
                  (N15413)? mem[446] : 
                  (N15414)? mem[448] : 
                  (N15415)? mem[450] : 
                  (N15416)? mem[452] : 
                  (N15417)? mem[454] : 
                  (N15418)? mem[456] : 
                  (N15419)? mem[458] : 
                  (N15420)? mem[460] : 
                  (N15421)? mem[462] : 
                  (N15422)? mem[464] : 
                  (N15423)? mem[466] : 
                  (N15424)? mem[468] : 
                  (N15425)? mem[470] : 
                  (N15426)? mem[472] : 
                  (N15427)? mem[474] : 
                  (N15428)? mem[476] : 
                  (N15429)? mem[478] : 
                  (N15430)? mem[480] : 
                  (N15431)? mem[482] : 
                  (N15432)? mem[484] : 
                  (N15433)? mem[486] : 
                  (N15434)? mem[488] : 
                  (N15435)? mem[490] : 
                  (N15436)? mem[492] : 
                  (N15437)? mem[494] : 
                  (N15438)? mem[496] : 
                  (N15439)? mem[498] : 
                  (N15440)? mem[500] : 
                  (N15441)? mem[502] : 
                  (N15442)? mem[504] : 
                  (N15443)? mem[506] : 
                  (N15444)? mem[508] : 
                  (N15445)? mem[510] : 
                  (N14999)? mem[512] : 
                  (N15001)? mem[514] : 
                  (N15003)? mem[516] : 
                  (N15005)? mem[518] : 
                  (N15007)? mem[520] : 
                  (N15009)? mem[522] : 
                  (N15011)? mem[524] : 
                  (N15013)? mem[526] : 
                  (N15015)? mem[528] : 
                  (N15017)? mem[530] : 
                  (N15019)? mem[532] : 
                  (N15021)? mem[534] : 
                  (N15023)? mem[536] : 
                  (N15025)? mem[538] : 
                  (N15027)? mem[540] : 
                  (N15029)? mem[542] : 
                  (N15031)? mem[544] : 
                  (N15033)? mem[546] : 
                  (N15035)? mem[548] : 
                  (N15037)? mem[550] : 
                  (N15039)? mem[552] : 
                  (N15041)? mem[554] : 
                  (N15043)? mem[556] : 
                  (N15045)? mem[558] : 
                  (N15047)? mem[560] : 
                  (N15049)? mem[562] : 
                  (N15051)? mem[564] : 
                  (N15053)? mem[566] : 
                  (N15055)? mem[568] : 
                  (N15057)? mem[570] : 
                  (N15059)? mem[572] : 
                  (N15061)? mem[574] : 
                  (N15063)? mem[576] : 
                  (N15065)? mem[578] : 
                  (N15067)? mem[580] : 
                  (N15069)? mem[582] : 
                  (N15071)? mem[584] : 
                  (N15073)? mem[586] : 
                  (N15075)? mem[588] : 
                  (N15077)? mem[590] : 
                  (N15079)? mem[592] : 
                  (N15081)? mem[594] : 
                  (N15083)? mem[596] : 
                  (N15085)? mem[598] : 
                  (N15087)? mem[600] : 
                  (N15089)? mem[602] : 
                  (N15091)? mem[604] : 
                  (N15093)? mem[606] : 
                  (N15095)? mem[608] : 
                  (N15097)? mem[610] : 
                  (N15099)? mem[612] : 
                  (N15101)? mem[614] : 
                  (N15103)? mem[616] : 
                  (N15105)? mem[618] : 
                  (N15107)? mem[620] : 
                  (N15109)? mem[622] : 
                  (N15111)? mem[624] : 
                  (N15113)? mem[626] : 
                  (N15115)? mem[628] : 
                  (N15117)? mem[630] : 
                  (N15119)? mem[632] : 
                  (N15121)? mem[634] : 
                  (N15123)? mem[636] : 
                  (N15125)? mem[638] : 
                  (N15127)? mem[640] : 
                  (N15129)? mem[642] : 
                  (N15131)? mem[644] : 
                  (N15133)? mem[646] : 
                  (N15135)? mem[648] : 
                  (N15137)? mem[650] : 
                  (N15139)? mem[652] : 
                  (N15141)? mem[654] : 
                  (N15143)? mem[656] : 
                  (N15145)? mem[658] : 
                  (N15147)? mem[660] : 
                  (N15149)? mem[662] : 
                  (N15151)? mem[664] : 
                  (N15153)? mem[666] : 
                  (N15155)? mem[668] : 
                  (N15157)? mem[670] : 
                  (N15159)? mem[672] : 
                  (N15161)? mem[674] : 
                  (N15163)? mem[676] : 
                  (N15165)? mem[678] : 
                  (N15167)? mem[680] : 
                  (N15169)? mem[682] : 
                  (N15171)? mem[684] : 
                  (N15173)? mem[686] : 
                  (N15175)? mem[688] : 
                  (N15177)? mem[690] : 
                  (N15179)? mem[692] : 
                  (N15181)? mem[694] : 
                  (N15183)? mem[696] : 
                  (N15185)? mem[698] : 
                  (N15187)? mem[700] : 
                  (N15189)? mem[702] : 
                  (N15191)? mem[704] : 
                  (N15193)? mem[706] : 
                  (N15195)? mem[708] : 
                  (N15197)? mem[710] : 
                  (N15199)? mem[712] : 
                  (N15201)? mem[714] : 
                  (N15203)? mem[716] : 
                  (N15205)? mem[718] : 
                  (N15207)? mem[720] : 
                  (N15209)? mem[722] : 
                  (N15211)? mem[724] : 
                  (N15213)? mem[726] : 
                  (N15215)? mem[728] : 
                  (N15217)? mem[730] : 
                  (N15219)? mem[732] : 
                  (N15221)? mem[734] : 
                  (N15223)? mem[736] : 
                  (N15225)? mem[738] : 
                  (N15227)? mem[740] : 
                  (N15229)? mem[742] : 
                  (N15231)? mem[744] : 
                  (N15233)? mem[746] : 
                  (N15235)? mem[748] : 
                  (N15237)? mem[750] : 
                  (N15239)? mem[752] : 
                  (N15241)? mem[754] : 
                  (N15243)? mem[756] : 
                  (N15245)? mem[758] : 
                  (N15247)? mem[760] : 
                  (N15249)? mem[762] : 
                  (N15251)? mem[764] : 
                  (N15253)? mem[766] : 
                  (N15255)? mem[768] : 
                  (N15257)? mem[770] : 
                  (N15259)? mem[772] : 
                  (N15261)? mem[774] : 
                  (N15263)? mem[776] : 
                  (N15265)? mem[778] : 
                  (N15267)? mem[780] : 
                  (N15269)? mem[782] : 
                  (N15271)? mem[784] : 
                  (N15273)? mem[786] : 
                  (N15275)? mem[788] : 
                  (N15277)? mem[790] : 
                  (N15279)? mem[792] : 
                  (N15281)? mem[794] : 
                  (N15283)? mem[796] : 
                  (N15285)? mem[798] : 
                  (N15287)? mem[800] : 
                  (N15289)? mem[802] : 
                  (N15291)? mem[804] : 
                  (N15293)? mem[806] : 
                  (N15295)? mem[808] : 
                  (N15297)? mem[810] : 
                  (N15299)? mem[812] : 
                  (N15301)? mem[814] : 
                  (N15303)? mem[816] : 
                  (N15305)? mem[818] : 
                  (N15307)? mem[820] : 
                  (N15309)? mem[822] : 
                  (N15311)? mem[824] : 
                  (N15313)? mem[826] : 
                  (N15315)? mem[828] : 
                  (N15317)? mem[830] : 
                  (N15319)? mem[832] : 
                  (N15321)? mem[834] : 
                  (N15323)? mem[836] : 
                  (N15325)? mem[838] : 
                  (N15327)? mem[840] : 
                  (N15329)? mem[842] : 
                  (N15331)? mem[844] : 
                  (N15333)? mem[846] : 
                  (N15335)? mem[848] : 
                  (N15337)? mem[850] : 
                  (N15339)? mem[852] : 
                  (N15341)? mem[854] : 
                  (N15343)? mem[856] : 
                  (N15345)? mem[858] : 
                  (N15347)? mem[860] : 
                  (N15349)? mem[862] : 
                  (N15351)? mem[864] : 
                  (N15353)? mem[866] : 
                  (N15355)? mem[868] : 
                  (N15357)? mem[870] : 
                  (N15359)? mem[872] : 
                  (N15361)? mem[874] : 
                  (N15363)? mem[876] : 
                  (N15365)? mem[878] : 
                  (N15367)? mem[880] : 
                  (N15369)? mem[882] : 
                  (N15371)? mem[884] : 
                  (N15373)? mem[886] : 
                  (N15375)? mem[888] : 
                  (N15377)? mem[890] : 
                  (N15379)? mem[892] : 
                  (N15381)? mem[894] : 
                  (N11985)? mem[896] : 
                  (N11987)? mem[898] : 
                  (N11989)? mem[900] : 
                  (N11991)? mem[902] : 
                  (N11993)? mem[904] : 
                  (N11995)? mem[906] : 
                  (N11997)? mem[908] : 
                  (N11999)? mem[910] : 
                  (N12001)? mem[912] : 
                  (N12003)? mem[914] : 
                  (N12005)? mem[916] : 
                  (N12007)? mem[918] : 
                  (N12009)? mem[920] : 
                  (N12011)? mem[922] : 
                  (N12013)? mem[924] : 
                  (N12015)? mem[926] : 
                  (N12017)? mem[928] : 
                  (N12019)? mem[930] : 
                  (N12021)? mem[932] : 
                  (N12023)? mem[934] : 
                  (N12025)? mem[936] : 
                  (N12027)? mem[938] : 
                  (N12029)? mem[940] : 
                  (N12031)? mem[942] : 
                  (N12033)? mem[944] : 
                  (N12035)? mem[946] : 
                  (N12037)? mem[948] : 
                  (N12039)? mem[950] : 
                  (N12041)? mem[952] : 
                  (N12043)? mem[954] : 
                  (N12045)? mem[956] : 
                  (N12047)? mem[958] : 
                  (N12049)? mem[960] : 
                  (N12051)? mem[962] : 
                  (N12053)? mem[964] : 
                  (N12055)? mem[966] : 
                  (N12057)? mem[968] : 
                  (N12059)? mem[970] : 
                  (N12061)? mem[972] : 
                  (N12063)? mem[974] : 
                  (N12065)? mem[976] : 
                  (N12067)? mem[978] : 
                  (N12069)? mem[980] : 
                  (N12071)? mem[982] : 
                  (N12073)? mem[984] : 
                  (N12075)? mem[986] : 
                  (N12077)? mem[988] : 
                  (N12079)? mem[990] : 
                  (N12081)? mem[992] : 
                  (N12083)? mem[994] : 
                  (N12085)? mem[996] : 
                  (N12087)? mem[998] : 
                  (N12089)? mem[1000] : 
                  (N12091)? mem[1002] : 
                  (N12093)? mem[1004] : 
                  (N12095)? mem[1006] : 
                  (N12097)? mem[1008] : 
                  (N12099)? mem[1010] : 
                  (N12101)? mem[1012] : 
                  (N12103)? mem[1014] : 
                  (N12105)? mem[1016] : 
                  (N12107)? mem[1018] : 
                  (N12109)? mem[1020] : 
                  (N12111)? mem[1022] : 1'b0;

  always @(posedge clk_i) begin
    if(N16495) begin
      mem_1023_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16495) begin
      mem_1022_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16494) begin
      mem_1021_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16494) begin
      mem_1020_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16493) begin
      mem_1019_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16493) begin
      mem_1018_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16492) begin
      mem_1017_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16492) begin
      mem_1016_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16491) begin
      mem_1015_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16491) begin
      mem_1014_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16490) begin
      mem_1013_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16490) begin
      mem_1012_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16489) begin
      mem_1011_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16489) begin
      mem_1010_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16488) begin
      mem_1009_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16488) begin
      mem_1008_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16487) begin
      mem_1007_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16487) begin
      mem_1006_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16486) begin
      mem_1005_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16486) begin
      mem_1004_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16485) begin
      mem_1003_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16485) begin
      mem_1002_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16484) begin
      mem_1001_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16484) begin
      mem_1000_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16483) begin
      mem_999_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16483) begin
      mem_998_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16482) begin
      mem_997_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16482) begin
      mem_996_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16481) begin
      mem_995_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16481) begin
      mem_994_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16480) begin
      mem_993_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16480) begin
      mem_992_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16479) begin
      mem_991_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16479) begin
      mem_990_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16478) begin
      mem_989_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16478) begin
      mem_988_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16477) begin
      mem_987_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16477) begin
      mem_986_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16476) begin
      mem_985_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16476) begin
      mem_984_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16475) begin
      mem_983_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16475) begin
      mem_982_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16474) begin
      mem_981_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16474) begin
      mem_980_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16473) begin
      mem_979_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16473) begin
      mem_978_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16472) begin
      mem_977_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16472) begin
      mem_976_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16471) begin
      mem_975_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16471) begin
      mem_974_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16470) begin
      mem_973_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16470) begin
      mem_972_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16469) begin
      mem_971_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16469) begin
      mem_970_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16468) begin
      mem_969_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16468) begin
      mem_968_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16467) begin
      mem_967_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16467) begin
      mem_966_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16466) begin
      mem_965_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16466) begin
      mem_964_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16465) begin
      mem_963_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16465) begin
      mem_962_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16464) begin
      mem_961_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16464) begin
      mem_960_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16463) begin
      mem_959_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16463) begin
      mem_958_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16462) begin
      mem_957_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16462) begin
      mem_956_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16461) begin
      mem_955_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16461) begin
      mem_954_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16460) begin
      mem_953_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16460) begin
      mem_952_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16459) begin
      mem_951_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16459) begin
      mem_950_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16458) begin
      mem_949_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16458) begin
      mem_948_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16457) begin
      mem_947_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16457) begin
      mem_946_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16456) begin
      mem_945_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16456) begin
      mem_944_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16455) begin
      mem_943_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16455) begin
      mem_942_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16454) begin
      mem_941_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16454) begin
      mem_940_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16453) begin
      mem_939_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16453) begin
      mem_938_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16452) begin
      mem_937_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16452) begin
      mem_936_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16451) begin
      mem_935_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16451) begin
      mem_934_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16450) begin
      mem_933_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16450) begin
      mem_932_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16449) begin
      mem_931_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16449) begin
      mem_930_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16448) begin
      mem_929_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16448) begin
      mem_928_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16447) begin
      mem_927_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16447) begin
      mem_926_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16446) begin
      mem_925_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16446) begin
      mem_924_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16445) begin
      mem_923_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16445) begin
      mem_922_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16444) begin
      mem_921_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16444) begin
      mem_920_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16443) begin
      mem_919_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16443) begin
      mem_918_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16442) begin
      mem_917_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16442) begin
      mem_916_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16441) begin
      mem_915_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16441) begin
      mem_914_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16440) begin
      mem_913_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16440) begin
      mem_912_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16439) begin
      mem_911_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16439) begin
      mem_910_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16438) begin
      mem_909_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16438) begin
      mem_908_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16437) begin
      mem_907_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16437) begin
      mem_906_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16436) begin
      mem_905_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16436) begin
      mem_904_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16435) begin
      mem_903_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16435) begin
      mem_902_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16434) begin
      mem_901_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16434) begin
      mem_900_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16433) begin
      mem_899_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16433) begin
      mem_898_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16432) begin
      mem_897_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16432) begin
      mem_896_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16431) begin
      mem_895_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16431) begin
      mem_894_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16430) begin
      mem_893_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16430) begin
      mem_892_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16429) begin
      mem_891_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16429) begin
      mem_890_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16428) begin
      mem_889_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16428) begin
      mem_888_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16427) begin
      mem_887_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16427) begin
      mem_886_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16426) begin
      mem_885_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16426) begin
      mem_884_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16425) begin
      mem_883_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16425) begin
      mem_882_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16424) begin
      mem_881_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16424) begin
      mem_880_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16423) begin
      mem_879_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16423) begin
      mem_878_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16422) begin
      mem_877_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16422) begin
      mem_876_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16421) begin
      mem_875_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16421) begin
      mem_874_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16420) begin
      mem_873_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16420) begin
      mem_872_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16419) begin
      mem_871_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16419) begin
      mem_870_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16418) begin
      mem_869_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16418) begin
      mem_868_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16417) begin
      mem_867_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16417) begin
      mem_866_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16416) begin
      mem_865_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16416) begin
      mem_864_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16415) begin
      mem_863_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16415) begin
      mem_862_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16414) begin
      mem_861_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16414) begin
      mem_860_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16413) begin
      mem_859_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16413) begin
      mem_858_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16412) begin
      mem_857_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16412) begin
      mem_856_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16411) begin
      mem_855_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16411) begin
      mem_854_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16410) begin
      mem_853_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16410) begin
      mem_852_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16409) begin
      mem_851_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16409) begin
      mem_850_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16408) begin
      mem_849_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16408) begin
      mem_848_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16407) begin
      mem_847_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16407) begin
      mem_846_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16406) begin
      mem_845_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16406) begin
      mem_844_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16405) begin
      mem_843_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16405) begin
      mem_842_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16404) begin
      mem_841_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16404) begin
      mem_840_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16403) begin
      mem_839_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16403) begin
      mem_838_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16402) begin
      mem_837_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16402) begin
      mem_836_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16401) begin
      mem_835_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16401) begin
      mem_834_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16400) begin
      mem_833_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16400) begin
      mem_832_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16399) begin
      mem_831_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16399) begin
      mem_830_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16398) begin
      mem_829_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16398) begin
      mem_828_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16397) begin
      mem_827_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N16397) begin
      mem_826_sv2v_reg <= N15973;
    end 
  end


  always @(posedge clk_i) begin
    if(N16396) begin
      mem_825_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16396) begin
      mem_824_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16395) begin
      mem_823_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16395) begin
      mem_822_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16394) begin
      mem_821_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16394) begin
      mem_820_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16393) begin
      mem_819_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16393) begin
      mem_818_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16392) begin
      mem_817_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16392) begin
      mem_816_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16391) begin
      mem_815_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16391) begin
      mem_814_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16390) begin
      mem_813_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16390) begin
      mem_812_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16389) begin
      mem_811_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16389) begin
      mem_810_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16388) begin
      mem_809_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16388) begin
      mem_808_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16387) begin
      mem_807_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16387) begin
      mem_806_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16386) begin
      mem_805_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16386) begin
      mem_804_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16385) begin
      mem_803_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16385) begin
      mem_802_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16384) begin
      mem_801_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16384) begin
      mem_800_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16383) begin
      mem_799_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16383) begin
      mem_798_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16382) begin
      mem_797_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16382) begin
      mem_796_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16381) begin
      mem_795_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16381) begin
      mem_794_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16380) begin
      mem_793_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16380) begin
      mem_792_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16379) begin
      mem_791_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16379) begin
      mem_790_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16378) begin
      mem_789_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16378) begin
      mem_788_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16377) begin
      mem_787_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16377) begin
      mem_786_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16376) begin
      mem_785_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16376) begin
      mem_784_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16375) begin
      mem_783_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16375) begin
      mem_782_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16374) begin
      mem_781_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16374) begin
      mem_780_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16373) begin
      mem_779_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16373) begin
      mem_778_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16372) begin
      mem_777_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16372) begin
      mem_776_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16371) begin
      mem_775_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16371) begin
      mem_774_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16370) begin
      mem_773_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16370) begin
      mem_772_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16369) begin
      mem_771_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16369) begin
      mem_770_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16368) begin
      mem_769_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16368) begin
      mem_768_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16367) begin
      mem_767_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16367) begin
      mem_766_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16366) begin
      mem_765_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16366) begin
      mem_764_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16365) begin
      mem_763_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16365) begin
      mem_762_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16364) begin
      mem_761_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16364) begin
      mem_760_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16363) begin
      mem_759_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16363) begin
      mem_758_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16362) begin
      mem_757_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16362) begin
      mem_756_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16361) begin
      mem_755_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16361) begin
      mem_754_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16360) begin
      mem_753_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16360) begin
      mem_752_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16359) begin
      mem_751_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16359) begin
      mem_750_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16358) begin
      mem_749_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16358) begin
      mem_748_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16357) begin
      mem_747_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16357) begin
      mem_746_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16356) begin
      mem_745_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16356) begin
      mem_744_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16355) begin
      mem_743_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16355) begin
      mem_742_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16354) begin
      mem_741_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16354) begin
      mem_740_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16353) begin
      mem_739_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16353) begin
      mem_738_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16352) begin
      mem_737_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16352) begin
      mem_736_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16351) begin
      mem_735_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16351) begin
      mem_734_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16350) begin
      mem_733_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16350) begin
      mem_732_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16349) begin
      mem_731_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16349) begin
      mem_730_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16348) begin
      mem_729_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16348) begin
      mem_728_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16347) begin
      mem_727_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16347) begin
      mem_726_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16346) begin
      mem_725_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16346) begin
      mem_724_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16345) begin
      mem_723_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16345) begin
      mem_722_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16344) begin
      mem_721_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16344) begin
      mem_720_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16343) begin
      mem_719_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16343) begin
      mem_718_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16342) begin
      mem_717_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16342) begin
      mem_716_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16341) begin
      mem_715_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16341) begin
      mem_714_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16340) begin
      mem_713_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16340) begin
      mem_712_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16339) begin
      mem_711_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16339) begin
      mem_710_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16338) begin
      mem_709_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16338) begin
      mem_708_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16337) begin
      mem_707_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16337) begin
      mem_706_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16336) begin
      mem_705_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16336) begin
      mem_704_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16335) begin
      mem_703_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16335) begin
      mem_702_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16334) begin
      mem_701_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16334) begin
      mem_700_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16333) begin
      mem_699_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16333) begin
      mem_698_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16332) begin
      mem_697_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16332) begin
      mem_696_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16331) begin
      mem_695_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16331) begin
      mem_694_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16330) begin
      mem_693_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16330) begin
      mem_692_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16329) begin
      mem_691_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16329) begin
      mem_690_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16328) begin
      mem_689_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16328) begin
      mem_688_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16327) begin
      mem_687_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16327) begin
      mem_686_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16326) begin
      mem_685_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16326) begin
      mem_684_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16325) begin
      mem_683_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16325) begin
      mem_682_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16324) begin
      mem_681_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16324) begin
      mem_680_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16323) begin
      mem_679_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16323) begin
      mem_678_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16322) begin
      mem_677_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16322) begin
      mem_676_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16321) begin
      mem_675_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16321) begin
      mem_674_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16320) begin
      mem_673_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16320) begin
      mem_672_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16319) begin
      mem_671_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16319) begin
      mem_670_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16318) begin
      mem_669_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16318) begin
      mem_668_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16317) begin
      mem_667_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16317) begin
      mem_666_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16316) begin
      mem_665_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16316) begin
      mem_664_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16315) begin
      mem_663_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16315) begin
      mem_662_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16314) begin
      mem_661_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16314) begin
      mem_660_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16313) begin
      mem_659_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16313) begin
      mem_658_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16312) begin
      mem_657_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16312) begin
      mem_656_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16311) begin
      mem_655_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16311) begin
      mem_654_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16310) begin
      mem_653_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16310) begin
      mem_652_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16309) begin
      mem_651_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16309) begin
      mem_650_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16308) begin
      mem_649_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16308) begin
      mem_648_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16307) begin
      mem_647_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16307) begin
      mem_646_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16306) begin
      mem_645_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16306) begin
      mem_644_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16305) begin
      mem_643_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16305) begin
      mem_642_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16304) begin
      mem_641_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16304) begin
      mem_640_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16303) begin
      mem_639_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16303) begin
      mem_638_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16302) begin
      mem_637_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16302) begin
      mem_636_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16301) begin
      mem_635_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16301) begin
      mem_634_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16300) begin
      mem_633_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16300) begin
      mem_632_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16299) begin
      mem_631_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16299) begin
      mem_630_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16298) begin
      mem_629_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N16298) begin
      mem_628_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N16297) begin
      mem_627_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16297) begin
      mem_626_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16296) begin
      mem_625_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16296) begin
      mem_624_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16295) begin
      mem_623_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16295) begin
      mem_622_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16294) begin
      mem_621_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16294) begin
      mem_620_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16293) begin
      mem_619_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16293) begin
      mem_618_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16292) begin
      mem_617_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16292) begin
      mem_616_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16291) begin
      mem_615_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16291) begin
      mem_614_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16290) begin
      mem_613_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16290) begin
      mem_612_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16289) begin
      mem_611_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16289) begin
      mem_610_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16288) begin
      mem_609_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16288) begin
      mem_608_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16287) begin
      mem_607_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16287) begin
      mem_606_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16286) begin
      mem_605_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16286) begin
      mem_604_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16285) begin
      mem_603_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16285) begin
      mem_602_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16284) begin
      mem_601_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16284) begin
      mem_600_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16283) begin
      mem_599_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16283) begin
      mem_598_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16282) begin
      mem_597_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16282) begin
      mem_596_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16281) begin
      mem_595_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16281) begin
      mem_594_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16280) begin
      mem_593_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16280) begin
      mem_592_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16279) begin
      mem_591_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16279) begin
      mem_590_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16278) begin
      mem_589_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16278) begin
      mem_588_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16277) begin
      mem_587_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16277) begin
      mem_586_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16276) begin
      mem_585_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16276) begin
      mem_584_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16275) begin
      mem_583_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16275) begin
      mem_582_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16274) begin
      mem_581_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16274) begin
      mem_580_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16273) begin
      mem_579_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16273) begin
      mem_578_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16272) begin
      mem_577_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16272) begin
      mem_576_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16271) begin
      mem_575_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16271) begin
      mem_574_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16270) begin
      mem_573_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16270) begin
      mem_572_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16269) begin
      mem_571_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16269) begin
      mem_570_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16268) begin
      mem_569_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16268) begin
      mem_568_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16267) begin
      mem_567_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16267) begin
      mem_566_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16266) begin
      mem_565_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16266) begin
      mem_564_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16265) begin
      mem_563_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16265) begin
      mem_562_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16264) begin
      mem_561_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16264) begin
      mem_560_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16263) begin
      mem_559_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16263) begin
      mem_558_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16262) begin
      mem_557_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16262) begin
      mem_556_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16261) begin
      mem_555_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16261) begin
      mem_554_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16260) begin
      mem_553_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16260) begin
      mem_552_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16259) begin
      mem_551_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16259) begin
      mem_550_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16258) begin
      mem_549_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16258) begin
      mem_548_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16257) begin
      mem_547_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16257) begin
      mem_546_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16256) begin
      mem_545_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16256) begin
      mem_544_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16255) begin
      mem_543_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16255) begin
      mem_542_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16254) begin
      mem_541_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16254) begin
      mem_540_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16253) begin
      mem_539_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16253) begin
      mem_538_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16252) begin
      mem_537_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16252) begin
      mem_536_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16251) begin
      mem_535_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16251) begin
      mem_534_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16250) begin
      mem_533_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16250) begin
      mem_532_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16249) begin
      mem_531_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16249) begin
      mem_530_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16248) begin
      mem_529_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16248) begin
      mem_528_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16247) begin
      mem_527_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16247) begin
      mem_526_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16246) begin
      mem_525_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16246) begin
      mem_524_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16245) begin
      mem_523_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16245) begin
      mem_522_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16244) begin
      mem_521_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16244) begin
      mem_520_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16243) begin
      mem_519_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16243) begin
      mem_518_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16242) begin
      mem_517_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16242) begin
      mem_516_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16241) begin
      mem_515_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16241) begin
      mem_514_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16240) begin
      mem_513_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16240) begin
      mem_512_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16239) begin
      mem_511_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16239) begin
      mem_510_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16238) begin
      mem_509_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16238) begin
      mem_508_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16237) begin
      mem_507_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16237) begin
      mem_506_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16236) begin
      mem_505_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16236) begin
      mem_504_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16235) begin
      mem_503_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16235) begin
      mem_502_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16234) begin
      mem_501_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16234) begin
      mem_500_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16233) begin
      mem_499_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16233) begin
      mem_498_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16232) begin
      mem_497_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16232) begin
      mem_496_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16231) begin
      mem_495_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16231) begin
      mem_494_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16230) begin
      mem_493_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16230) begin
      mem_492_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16229) begin
      mem_491_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16229) begin
      mem_490_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16228) begin
      mem_489_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16228) begin
      mem_488_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16227) begin
      mem_487_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16227) begin
      mem_486_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16226) begin
      mem_485_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16226) begin
      mem_484_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16225) begin
      mem_483_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16225) begin
      mem_482_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16224) begin
      mem_481_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16224) begin
      mem_480_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16223) begin
      mem_479_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16223) begin
      mem_478_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16222) begin
      mem_477_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16222) begin
      mem_476_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16221) begin
      mem_475_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16221) begin
      mem_474_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16220) begin
      mem_473_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16220) begin
      mem_472_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16219) begin
      mem_471_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16219) begin
      mem_470_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16218) begin
      mem_469_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16218) begin
      mem_468_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16217) begin
      mem_467_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16217) begin
      mem_466_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16216) begin
      mem_465_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16216) begin
      mem_464_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16215) begin
      mem_463_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16215) begin
      mem_462_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16214) begin
      mem_461_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16214) begin
      mem_460_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16213) begin
      mem_459_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16213) begin
      mem_458_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16212) begin
      mem_457_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16212) begin
      mem_456_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16211) begin
      mem_455_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16211) begin
      mem_454_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16210) begin
      mem_453_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16210) begin
      mem_452_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16209) begin
      mem_451_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16209) begin
      mem_450_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16208) begin
      mem_449_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16208) begin
      mem_448_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16207) begin
      mem_447_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16207) begin
      mem_446_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16206) begin
      mem_445_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16206) begin
      mem_444_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16205) begin
      mem_443_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16205) begin
      mem_442_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16204) begin
      mem_441_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16204) begin
      mem_440_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16203) begin
      mem_439_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16203) begin
      mem_438_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16202) begin
      mem_437_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16202) begin
      mem_436_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16201) begin
      mem_435_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16201) begin
      mem_434_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16200) begin
      mem_433_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16200) begin
      mem_432_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16199) begin
      mem_431_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N16199) begin
      mem_430_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N16198) begin
      mem_429_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16198) begin
      mem_428_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16197) begin
      mem_427_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16197) begin
      mem_426_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16196) begin
      mem_425_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16196) begin
      mem_424_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16195) begin
      mem_423_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16195) begin
      mem_422_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16194) begin
      mem_421_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16194) begin
      mem_420_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16193) begin
      mem_419_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16193) begin
      mem_418_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16192) begin
      mem_417_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16192) begin
      mem_416_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16191) begin
      mem_415_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16191) begin
      mem_414_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16190) begin
      mem_413_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16190) begin
      mem_412_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16189) begin
      mem_411_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16189) begin
      mem_410_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16188) begin
      mem_409_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16188) begin
      mem_408_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16187) begin
      mem_407_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16187) begin
      mem_406_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16186) begin
      mem_405_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16186) begin
      mem_404_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16185) begin
      mem_403_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16185) begin
      mem_402_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16184) begin
      mem_401_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16184) begin
      mem_400_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16183) begin
      mem_399_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16183) begin
      mem_398_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16182) begin
      mem_397_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16182) begin
      mem_396_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16181) begin
      mem_395_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16181) begin
      mem_394_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16180) begin
      mem_393_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16180) begin
      mem_392_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16179) begin
      mem_391_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16179) begin
      mem_390_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16178) begin
      mem_389_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16178) begin
      mem_388_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16177) begin
      mem_387_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16177) begin
      mem_386_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16176) begin
      mem_385_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16176) begin
      mem_384_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16175) begin
      mem_383_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16175) begin
      mem_382_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16174) begin
      mem_381_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16174) begin
      mem_380_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16173) begin
      mem_379_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16173) begin
      mem_378_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16172) begin
      mem_377_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16172) begin
      mem_376_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16171) begin
      mem_375_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16171) begin
      mem_374_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16170) begin
      mem_373_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16170) begin
      mem_372_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16169) begin
      mem_371_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16169) begin
      mem_370_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16168) begin
      mem_369_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16168) begin
      mem_368_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16167) begin
      mem_367_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16167) begin
      mem_366_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16166) begin
      mem_365_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16166) begin
      mem_364_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16165) begin
      mem_363_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16165) begin
      mem_362_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16164) begin
      mem_361_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16164) begin
      mem_360_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16163) begin
      mem_359_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16163) begin
      mem_358_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16162) begin
      mem_357_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16162) begin
      mem_356_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16161) begin
      mem_355_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16161) begin
      mem_354_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16160) begin
      mem_353_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16160) begin
      mem_352_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16159) begin
      mem_351_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16159) begin
      mem_350_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16158) begin
      mem_349_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16158) begin
      mem_348_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16157) begin
      mem_347_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16157) begin
      mem_346_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16156) begin
      mem_345_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16156) begin
      mem_344_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16155) begin
      mem_343_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16155) begin
      mem_342_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16154) begin
      mem_341_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16154) begin
      mem_340_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16153) begin
      mem_339_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16153) begin
      mem_338_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16152) begin
      mem_337_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16152) begin
      mem_336_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16151) begin
      mem_335_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16151) begin
      mem_334_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16150) begin
      mem_333_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16150) begin
      mem_332_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16149) begin
      mem_331_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16149) begin
      mem_330_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16148) begin
      mem_329_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16148) begin
      mem_328_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16147) begin
      mem_327_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16147) begin
      mem_326_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16146) begin
      mem_325_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16146) begin
      mem_324_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16145) begin
      mem_323_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16145) begin
      mem_322_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16144) begin
      mem_321_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16144) begin
      mem_320_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16143) begin
      mem_319_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16143) begin
      mem_318_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16142) begin
      mem_317_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16142) begin
      mem_316_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16141) begin
      mem_315_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16141) begin
      mem_314_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16140) begin
      mem_313_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16140) begin
      mem_312_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16139) begin
      mem_311_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16139) begin
      mem_310_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16138) begin
      mem_309_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16138) begin
      mem_308_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16137) begin
      mem_307_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16137) begin
      mem_306_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16136) begin
      mem_305_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16136) begin
      mem_304_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16135) begin
      mem_303_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16135) begin
      mem_302_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16134) begin
      mem_301_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16134) begin
      mem_300_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16133) begin
      mem_299_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16133) begin
      mem_298_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16132) begin
      mem_297_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16132) begin
      mem_296_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16131) begin
      mem_295_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16131) begin
      mem_294_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16130) begin
      mem_293_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16130) begin
      mem_292_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16129) begin
      mem_291_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16129) begin
      mem_290_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16128) begin
      mem_289_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16128) begin
      mem_288_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16127) begin
      mem_287_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16127) begin
      mem_286_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16126) begin
      mem_285_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16126) begin
      mem_284_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16125) begin
      mem_283_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16125) begin
      mem_282_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16124) begin
      mem_281_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16124) begin
      mem_280_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16123) begin
      mem_279_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16123) begin
      mem_278_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16122) begin
      mem_277_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16122) begin
      mem_276_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16121) begin
      mem_275_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16121) begin
      mem_274_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16120) begin
      mem_273_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16120) begin
      mem_272_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16119) begin
      mem_271_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16119) begin
      mem_270_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16118) begin
      mem_269_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16118) begin
      mem_268_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16117) begin
      mem_267_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16117) begin
      mem_266_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16116) begin
      mem_265_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16116) begin
      mem_264_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16115) begin
      mem_263_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16115) begin
      mem_262_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16114) begin
      mem_261_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16114) begin
      mem_260_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16113) begin
      mem_259_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16113) begin
      mem_258_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16112) begin
      mem_257_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16112) begin
      mem_256_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16111) begin
      mem_255_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16111) begin
      mem_254_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16110) begin
      mem_253_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16110) begin
      mem_252_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16109) begin
      mem_251_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16109) begin
      mem_250_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16108) begin
      mem_249_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16108) begin
      mem_248_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16107) begin
      mem_247_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16107) begin
      mem_246_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16106) begin
      mem_245_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16106) begin
      mem_244_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16105) begin
      mem_243_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16105) begin
      mem_242_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16104) begin
      mem_241_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16104) begin
      mem_240_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16103) begin
      mem_239_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16103) begin
      mem_238_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16102) begin
      mem_237_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16102) begin
      mem_236_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16101) begin
      mem_235_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16101) begin
      mem_234_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16100) begin
      mem_233_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N16100) begin
      mem_232_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N16099) begin
      mem_231_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16099) begin
      mem_230_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16098) begin
      mem_229_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16098) begin
      mem_228_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16097) begin
      mem_227_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16097) begin
      mem_226_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16096) begin
      mem_225_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16096) begin
      mem_224_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16095) begin
      mem_223_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16095) begin
      mem_222_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16094) begin
      mem_221_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16094) begin
      mem_220_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16093) begin
      mem_219_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16093) begin
      mem_218_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16092) begin
      mem_217_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16092) begin
      mem_216_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16091) begin
      mem_215_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16091) begin
      mem_214_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16090) begin
      mem_213_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16090) begin
      mem_212_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16089) begin
      mem_211_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16089) begin
      mem_210_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16088) begin
      mem_209_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16088) begin
      mem_208_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16087) begin
      mem_207_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16087) begin
      mem_206_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16086) begin
      mem_205_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16086) begin
      mem_204_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16085) begin
      mem_203_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16085) begin
      mem_202_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16084) begin
      mem_201_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16084) begin
      mem_200_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16083) begin
      mem_199_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16083) begin
      mem_198_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16082) begin
      mem_197_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16082) begin
      mem_196_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16081) begin
      mem_195_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16081) begin
      mem_194_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16080) begin
      mem_193_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16080) begin
      mem_192_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16079) begin
      mem_191_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16079) begin
      mem_190_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16078) begin
      mem_189_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16078) begin
      mem_188_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16077) begin
      mem_187_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16077) begin
      mem_186_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16076) begin
      mem_185_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16076) begin
      mem_184_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16075) begin
      mem_183_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16075) begin
      mem_182_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16074) begin
      mem_181_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16074) begin
      mem_180_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16073) begin
      mem_179_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16073) begin
      mem_178_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16072) begin
      mem_177_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16072) begin
      mem_176_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16071) begin
      mem_175_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16071) begin
      mem_174_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16070) begin
      mem_173_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16070) begin
      mem_172_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16069) begin
      mem_171_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16069) begin
      mem_170_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16068) begin
      mem_169_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16068) begin
      mem_168_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16067) begin
      mem_167_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16067) begin
      mem_166_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16066) begin
      mem_165_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16066) begin
      mem_164_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16065) begin
      mem_163_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16065) begin
      mem_162_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16064) begin
      mem_161_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16064) begin
      mem_160_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16063) begin
      mem_159_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16063) begin
      mem_158_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16062) begin
      mem_157_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16062) begin
      mem_156_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16061) begin
      mem_155_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16061) begin
      mem_154_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16060) begin
      mem_153_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16060) begin
      mem_152_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16059) begin
      mem_151_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16059) begin
      mem_150_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16058) begin
      mem_149_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16058) begin
      mem_148_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16057) begin
      mem_147_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16057) begin
      mem_146_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16056) begin
      mem_145_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16056) begin
      mem_144_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16055) begin
      mem_143_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16055) begin
      mem_142_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16054) begin
      mem_141_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16054) begin
      mem_140_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16053) begin
      mem_139_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16053) begin
      mem_138_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16052) begin
      mem_137_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16052) begin
      mem_136_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16051) begin
      mem_135_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16051) begin
      mem_134_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16050) begin
      mem_133_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16050) begin
      mem_132_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16049) begin
      mem_131_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16049) begin
      mem_130_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16048) begin
      mem_129_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16048) begin
      mem_128_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16047) begin
      mem_127_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16047) begin
      mem_126_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16046) begin
      mem_125_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16046) begin
      mem_124_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16045) begin
      mem_123_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16045) begin
      mem_122_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16044) begin
      mem_121_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16044) begin
      mem_120_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16043) begin
      mem_119_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16043) begin
      mem_118_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16042) begin
      mem_117_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16042) begin
      mem_116_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16041) begin
      mem_115_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16041) begin
      mem_114_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16040) begin
      mem_113_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16040) begin
      mem_112_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16039) begin
      mem_111_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16039) begin
      mem_110_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16038) begin
      mem_109_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16038) begin
      mem_108_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16037) begin
      mem_107_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16037) begin
      mem_106_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16036) begin
      mem_105_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16036) begin
      mem_104_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16035) begin
      mem_103_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16035) begin
      mem_102_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16034) begin
      mem_101_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16034) begin
      mem_100_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16033) begin
      mem_99_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16033) begin
      mem_98_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16032) begin
      mem_97_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16032) begin
      mem_96_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16031) begin
      mem_95_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16031) begin
      mem_94_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16030) begin
      mem_93_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16030) begin
      mem_92_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16029) begin
      mem_91_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16029) begin
      mem_90_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16028) begin
      mem_89_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16028) begin
      mem_88_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16027) begin
      mem_87_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16027) begin
      mem_86_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16026) begin
      mem_85_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16026) begin
      mem_84_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16025) begin
      mem_83_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16025) begin
      mem_82_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16024) begin
      mem_81_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16024) begin
      mem_80_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16023) begin
      mem_79_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16023) begin
      mem_78_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16022) begin
      mem_77_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16022) begin
      mem_76_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16021) begin
      mem_75_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16021) begin
      mem_74_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16020) begin
      mem_73_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16020) begin
      mem_72_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16019) begin
      mem_71_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16019) begin
      mem_70_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16018) begin
      mem_69_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16018) begin
      mem_68_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16017) begin
      mem_67_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16017) begin
      mem_66_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16016) begin
      mem_65_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16016) begin
      mem_64_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16015) begin
      mem_63_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16015) begin
      mem_62_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16014) begin
      mem_61_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16014) begin
      mem_60_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16013) begin
      mem_59_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16013) begin
      mem_58_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16012) begin
      mem_57_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16012) begin
      mem_56_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16011) begin
      mem_55_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16011) begin
      mem_54_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16010) begin
      mem_53_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16010) begin
      mem_52_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16009) begin
      mem_51_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16009) begin
      mem_50_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16008) begin
      mem_49_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16008) begin
      mem_48_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16007) begin
      mem_47_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16007) begin
      mem_46_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16006) begin
      mem_45_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16006) begin
      mem_44_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16005) begin
      mem_43_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16005) begin
      mem_42_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16004) begin
      mem_41_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16004) begin
      mem_40_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16003) begin
      mem_39_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16003) begin
      mem_38_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16002) begin
      mem_37_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16002) begin
      mem_36_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16001) begin
      mem_35_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N16001) begin
      mem_34_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N16000) begin
      mem_33_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N16000) begin
      mem_32_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15999) begin
      mem_31_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15999) begin
      mem_30_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15998) begin
      mem_29_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15998) begin
      mem_28_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15997) begin
      mem_27_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15997) begin
      mem_26_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15996) begin
      mem_25_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15996) begin
      mem_24_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15995) begin
      mem_23_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15995) begin
      mem_22_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15994) begin
      mem_21_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15994) begin
      mem_20_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15993) begin
      mem_19_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15993) begin
      mem_18_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15992) begin
      mem_17_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15992) begin
      mem_16_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15991) begin
      mem_15_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15991) begin
      mem_14_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15990) begin
      mem_13_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15990) begin
      mem_12_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15987) begin
      mem_11_sv2v_reg <= N15989;
    end 
  end


  always @(posedge clk_i) begin
    if(N15987) begin
      mem_10_sv2v_reg <= N15988;
    end 
  end


  always @(posedge clk_i) begin
    if(N15984) begin
      mem_9_sv2v_reg <= N15986;
    end 
  end


  always @(posedge clk_i) begin
    if(N15984) begin
      mem_8_sv2v_reg <= N15985;
    end 
  end


  always @(posedge clk_i) begin
    if(N15981) begin
      mem_7_sv2v_reg <= N15983;
    end 
  end


  always @(posedge clk_i) begin
    if(N15981) begin
      mem_6_sv2v_reg <= N15982;
    end 
  end


  always @(posedge clk_i) begin
    if(N15978) begin
      mem_5_sv2v_reg <= N15980;
    end 
  end


  always @(posedge clk_i) begin
    if(N15978) begin
      mem_4_sv2v_reg <= N15979;
    end 
  end


  always @(posedge clk_i) begin
    if(N15975) begin
      mem_3_sv2v_reg <= N15977;
    end 
  end


  always @(posedge clk_i) begin
    if(N15975) begin
      mem_2_sv2v_reg <= N15976;
    end 
  end


  always @(posedge clk_i) begin
    if(N15972) begin
      mem_1_sv2v_reg <= N15974;
    end 
  end


  always @(posedge clk_i) begin
    if(N15972) begin
      mem_0_sv2v_reg <= N15973;
    end 
  end

  assign N16498 = idx_w_i[7] & idx_w_i[8];
  assign N16499 = N0 & idx_w_i[8];
  assign N0 = ~idx_w_i[7];
  assign N16500 = idx_w_i[7] & N1;
  assign N1 = ~idx_w_i[8];
  assign N16501 = N2 & N3;
  assign N2 = ~idx_w_i[7];
  assign N3 = ~idx_w_i[8];
  assign N16502 = idx_w_i[5] & idx_w_i[6];
  assign N16503 = N4 & idx_w_i[6];
  assign N4 = ~idx_w_i[5];
  assign N16504 = idx_w_i[5] & N5;
  assign N5 = ~idx_w_i[6];
  assign N16505 = N6 & N7;
  assign N6 = ~idx_w_i[5];
  assign N7 = ~idx_w_i[6];
  assign N16506 = N16498 & N16502;
  assign N16507 = N16498 & N16503;
  assign N16508 = N16498 & N16504;
  assign N16509 = N16498 & N16505;
  assign N16510 = N16499 & N16502;
  assign N16511 = N16499 & N16503;
  assign N16512 = N16499 & N16504;
  assign N16513 = N16499 & N16505;
  assign N16514 = N16500 & N16502;
  assign N16515 = N16500 & N16503;
  assign N16516 = N16500 & N16504;
  assign N16517 = N16500 & N16505;
  assign N16518 = N16501 & N16502;
  assign N16519 = N16501 & N16503;
  assign N16520 = N16501 & N16504;
  assign N16521 = N16501 & N16505;
  assign N16522 = idx_w_i[3] & idx_w_i[4];
  assign N16523 = N8 & idx_w_i[4];
  assign N8 = ~idx_w_i[3];
  assign N16524 = idx_w_i[3] & N9;
  assign N9 = ~idx_w_i[4];
  assign N16525 = N10 & N11;
  assign N10 = ~idx_w_i[3];
  assign N11 = ~idx_w_i[4];
  assign N16526 = ~idx_w_i[2];
  assign N16527 = idx_w_i[0] & idx_w_i[1];
  assign N16528 = N12 & idx_w_i[1];
  assign N12 = ~idx_w_i[0];
  assign N16529 = idx_w_i[0] & N13;
  assign N13 = ~idx_w_i[1];
  assign N16530 = N14 & N15;
  assign N14 = ~idx_w_i[0];
  assign N15 = ~idx_w_i[1];
  assign N16531 = idx_w_i[2] & N16527;
  assign N16532 = idx_w_i[2] & N16528;
  assign N16533 = idx_w_i[2] & N16529;
  assign N16534 = idx_w_i[2] & N16530;
  assign N16535 = N16526 & N16527;
  assign N16536 = N16526 & N16528;
  assign N16537 = N16526 & N16529;
  assign N16538 = N16526 & N16530;
  assign N16539 = N16522 & N16531;
  assign N16540 = N16522 & N16532;
  assign N16541 = N16522 & N16533;
  assign N16542 = N16522 & N16534;
  assign N16543 = N16522 & N16535;
  assign N16544 = N16522 & N16536;
  assign N16545 = N16522 & N16537;
  assign N16546 = N16522 & N16538;
  assign N16547 = N16523 & N16531;
  assign N16548 = N16523 & N16532;
  assign N16549 = N16523 & N16533;
  assign N16550 = N16523 & N16534;
  assign N16551 = N16523 & N16535;
  assign N16552 = N16523 & N16536;
  assign N16553 = N16523 & N16537;
  assign N16554 = N16523 & N16538;
  assign N16555 = N16524 & N16531;
  assign N16556 = N16524 & N16532;
  assign N16557 = N16524 & N16533;
  assign N16558 = N16524 & N16534;
  assign N16559 = N16524 & N16535;
  assign N16560 = N16524 & N16536;
  assign N16561 = N16524 & N16537;
  assign N16562 = N16524 & N16538;
  assign N16563 = N16525 & N16531;
  assign N16564 = N16525 & N16532;
  assign N16565 = N16525 & N16533;
  assign N16566 = N16525 & N16534;
  assign N16567 = N16525 & N16535;
  assign N16568 = N16525 & N16536;
  assign N16569 = N16525 & N16537;
  assign N16570 = N16525 & N16538;
  assign N5076 = N16506 & N16539;
  assign N5075 = N16506 & N16540;
  assign N5074 = N16506 & N16541;
  assign N5073 = N16506 & N16542;
  assign N5072 = N16506 & N16543;
  assign N5071 = N16506 & N16544;
  assign N5070 = N16506 & N16545;
  assign N5069 = N16506 & N16546;
  assign N5068 = N16506 & N16547;
  assign N5067 = N16506 & N16548;
  assign N5066 = N16506 & N16549;
  assign N5065 = N16506 & N16550;
  assign N5064 = N16506 & N16551;
  assign N5063 = N16506 & N16552;
  assign N5062 = N16506 & N16553;
  assign N5061 = N16506 & N16554;
  assign N5060 = N16506 & N16555;
  assign N5059 = N16506 & N16556;
  assign N5058 = N16506 & N16557;
  assign N5057 = N16506 & N16558;
  assign N5056 = N16506 & N16559;
  assign N5055 = N16506 & N16560;
  assign N5054 = N16506 & N16561;
  assign N5053 = N16506 & N16562;
  assign N5052 = N16506 & N16563;
  assign N5051 = N16506 & N16564;
  assign N5050 = N16506 & N16565;
  assign N5049 = N16506 & N16566;
  assign N5048 = N16506 & N16567;
  assign N5047 = N16506 & N16568;
  assign N5046 = N16506 & N16569;
  assign N5045 = N16506 & N16570;
  assign N5044 = N16507 & N16539;
  assign N5043 = N16507 & N16540;
  assign N5042 = N16507 & N16541;
  assign N5041 = N16507 & N16542;
  assign N5040 = N16507 & N16543;
  assign N5039 = N16507 & N16544;
  assign N5038 = N16507 & N16545;
  assign N5037 = N16507 & N16546;
  assign N5036 = N16507 & N16547;
  assign N5035 = N16507 & N16548;
  assign N5034 = N16507 & N16549;
  assign N5033 = N16507 & N16550;
  assign N5032 = N16507 & N16551;
  assign N5031 = N16507 & N16552;
  assign N5030 = N16507 & N16553;
  assign N5029 = N16507 & N16554;
  assign N5028 = N16507 & N16555;
  assign N5027 = N16507 & N16556;
  assign N5026 = N16507 & N16557;
  assign N5025 = N16507 & N16558;
  assign N5024 = N16507 & N16559;
  assign N5023 = N16507 & N16560;
  assign N5022 = N16507 & N16561;
  assign N5021 = N16507 & N16562;
  assign N5020 = N16507 & N16563;
  assign N5019 = N16507 & N16564;
  assign N5018 = N16507 & N16565;
  assign N5017 = N16507 & N16566;
  assign N5016 = N16507 & N16567;
  assign N5015 = N16507 & N16568;
  assign N5014 = N16507 & N16569;
  assign N5013 = N16507 & N16570;
  assign N5012 = N16508 & N16539;
  assign N5011 = N16508 & N16540;
  assign N5010 = N16508 & N16541;
  assign N5009 = N16508 & N16542;
  assign N5008 = N16508 & N16543;
  assign N5007 = N16508 & N16544;
  assign N5006 = N16508 & N16545;
  assign N5005 = N16508 & N16546;
  assign N5004 = N16508 & N16547;
  assign N5003 = N16508 & N16548;
  assign N5002 = N16508 & N16549;
  assign N5001 = N16508 & N16550;
  assign N5000 = N16508 & N16551;
  assign N4999 = N16508 & N16552;
  assign N4998 = N16508 & N16553;
  assign N4997 = N16508 & N16554;
  assign N4996 = N16508 & N16555;
  assign N4995 = N16508 & N16556;
  assign N4994 = N16508 & N16557;
  assign N4993 = N16508 & N16558;
  assign N4992 = N16508 & N16559;
  assign N4991 = N16508 & N16560;
  assign N4990 = N16508 & N16561;
  assign N4989 = N16508 & N16562;
  assign N4988 = N16508 & N16563;
  assign N4987 = N16508 & N16564;
  assign N4986 = N16508 & N16565;
  assign N4985 = N16508 & N16566;
  assign N4984 = N16508 & N16567;
  assign N4983 = N16508 & N16568;
  assign N4982 = N16508 & N16569;
  assign N4981 = N16508 & N16570;
  assign N4980 = N16509 & N16539;
  assign N4979 = N16509 & N16540;
  assign N4978 = N16509 & N16541;
  assign N4977 = N16509 & N16542;
  assign N4976 = N16509 & N16543;
  assign N4975 = N16509 & N16544;
  assign N4974 = N16509 & N16545;
  assign N4973 = N16509 & N16546;
  assign N4972 = N16509 & N16547;
  assign N4971 = N16509 & N16548;
  assign N4970 = N16509 & N16549;
  assign N4969 = N16509 & N16550;
  assign N4968 = N16509 & N16551;
  assign N4967 = N16509 & N16552;
  assign N4966 = N16509 & N16553;
  assign N4965 = N16509 & N16554;
  assign N4964 = N16509 & N16555;
  assign N4963 = N16509 & N16556;
  assign N4962 = N16509 & N16557;
  assign N4961 = N16509 & N16558;
  assign N4960 = N16509 & N16559;
  assign N4959 = N16509 & N16560;
  assign N4958 = N16509 & N16561;
  assign N4957 = N16509 & N16562;
  assign N4956 = N16509 & N16563;
  assign N4955 = N16509 & N16564;
  assign N4954 = N16509 & N16565;
  assign N4953 = N16509 & N16566;
  assign N4952 = N16509 & N16567;
  assign N4951 = N16509 & N16568;
  assign N4950 = N16509 & N16569;
  assign N4949 = N16509 & N16570;
  assign N4948 = N16510 & N16539;
  assign N4947 = N16510 & N16540;
  assign N4946 = N16510 & N16541;
  assign N4945 = N16510 & N16542;
  assign N4944 = N16510 & N16543;
  assign N4943 = N16510 & N16544;
  assign N4942 = N16510 & N16545;
  assign N4941 = N16510 & N16546;
  assign N4940 = N16510 & N16547;
  assign N4939 = N16510 & N16548;
  assign N4938 = N16510 & N16549;
  assign N4937 = N16510 & N16550;
  assign N4936 = N16510 & N16551;
  assign N4935 = N16510 & N16552;
  assign N4934 = N16510 & N16553;
  assign N4933 = N16510 & N16554;
  assign N4932 = N16510 & N16555;
  assign N4931 = N16510 & N16556;
  assign N4930 = N16510 & N16557;
  assign N4929 = N16510 & N16558;
  assign N4928 = N16510 & N16559;
  assign N4927 = N16510 & N16560;
  assign N4926 = N16510 & N16561;
  assign N4925 = N16510 & N16562;
  assign N4924 = N16510 & N16563;
  assign N4923 = N16510 & N16564;
  assign N4922 = N16510 & N16565;
  assign N4921 = N16510 & N16566;
  assign N4920 = N16510 & N16567;
  assign N4919 = N16510 & N16568;
  assign N4918 = N16510 & N16569;
  assign N4917 = N16510 & N16570;
  assign N4916 = N16511 & N16539;
  assign N4915 = N16511 & N16540;
  assign N4914 = N16511 & N16541;
  assign N4913 = N16511 & N16542;
  assign N4912 = N16511 & N16543;
  assign N4911 = N16511 & N16544;
  assign N4910 = N16511 & N16545;
  assign N4909 = N16511 & N16546;
  assign N4908 = N16511 & N16547;
  assign N4907 = N16511 & N16548;
  assign N4906 = N16511 & N16549;
  assign N4905 = N16511 & N16550;
  assign N4904 = N16511 & N16551;
  assign N4903 = N16511 & N16552;
  assign N4902 = N16511 & N16553;
  assign N4901 = N16511 & N16554;
  assign N4900 = N16511 & N16555;
  assign N4899 = N16511 & N16556;
  assign N4898 = N16511 & N16557;
  assign N4897 = N16511 & N16558;
  assign N4896 = N16511 & N16559;
  assign N4895 = N16511 & N16560;
  assign N4894 = N16511 & N16561;
  assign N4893 = N16511 & N16562;
  assign N4892 = N16511 & N16563;
  assign N4891 = N16511 & N16564;
  assign N4890 = N16511 & N16565;
  assign N4889 = N16511 & N16566;
  assign N4888 = N16511 & N16567;
  assign N4887 = N16511 & N16568;
  assign N4886 = N16511 & N16569;
  assign N4885 = N16511 & N16570;
  assign N4884 = N16512 & N16539;
  assign N4883 = N16512 & N16540;
  assign N4882 = N16512 & N16541;
  assign N4881 = N16512 & N16542;
  assign N4880 = N16512 & N16543;
  assign N4879 = N16512 & N16544;
  assign N4878 = N16512 & N16545;
  assign N4877 = N16512 & N16546;
  assign N4876 = N16512 & N16547;
  assign N4875 = N16512 & N16548;
  assign N4874 = N16512 & N16549;
  assign N4873 = N16512 & N16550;
  assign N4872 = N16512 & N16551;
  assign N4871 = N16512 & N16552;
  assign N4870 = N16512 & N16553;
  assign N4869 = N16512 & N16554;
  assign N4868 = N16512 & N16555;
  assign N4867 = N16512 & N16556;
  assign N4866 = N16512 & N16557;
  assign N4865 = N16512 & N16558;
  assign N4864 = N16512 & N16559;
  assign N4863 = N16512 & N16560;
  assign N4862 = N16512 & N16561;
  assign N4861 = N16512 & N16562;
  assign N4860 = N16512 & N16563;
  assign N4859 = N16512 & N16564;
  assign N4858 = N16512 & N16565;
  assign N4857 = N16512 & N16566;
  assign N4856 = N16512 & N16567;
  assign N4855 = N16512 & N16568;
  assign N4854 = N16512 & N16569;
  assign N4853 = N16512 & N16570;
  assign N4852 = N16513 & N16539;
  assign N4851 = N16513 & N16540;
  assign N4850 = N16513 & N16541;
  assign N4849 = N16513 & N16542;
  assign N4848 = N16513 & N16543;
  assign N4847 = N16513 & N16544;
  assign N4846 = N16513 & N16545;
  assign N4845 = N16513 & N16546;
  assign N4844 = N16513 & N16547;
  assign N4843 = N16513 & N16548;
  assign N4842 = N16513 & N16549;
  assign N4841 = N16513 & N16550;
  assign N4840 = N16513 & N16551;
  assign N4839 = N16513 & N16552;
  assign N4838 = N16513 & N16553;
  assign N4837 = N16513 & N16554;
  assign N4836 = N16513 & N16555;
  assign N4835 = N16513 & N16556;
  assign N4834 = N16513 & N16557;
  assign N4833 = N16513 & N16558;
  assign N4832 = N16513 & N16559;
  assign N4831 = N16513 & N16560;
  assign N4830 = N16513 & N16561;
  assign N4829 = N16513 & N16562;
  assign N4828 = N16513 & N16563;
  assign N4827 = N16513 & N16564;
  assign N4826 = N16513 & N16565;
  assign N4825 = N16513 & N16566;
  assign N4824 = N16513 & N16567;
  assign N4823 = N16513 & N16568;
  assign N4822 = N16513 & N16569;
  assign N4821 = N16513 & N16570;
  assign N4820 = N16514 & N16539;
  assign N4819 = N16514 & N16540;
  assign N4818 = N16514 & N16541;
  assign N4817 = N16514 & N16542;
  assign N4816 = N16514 & N16543;
  assign N4815 = N16514 & N16544;
  assign N4814 = N16514 & N16545;
  assign N4813 = N16514 & N16546;
  assign N4812 = N16514 & N16547;
  assign N4811 = N16514 & N16548;
  assign N4810 = N16514 & N16549;
  assign N4809 = N16514 & N16550;
  assign N4808 = N16514 & N16551;
  assign N4807 = N16514 & N16552;
  assign N4806 = N16514 & N16553;
  assign N4805 = N16514 & N16554;
  assign N4804 = N16514 & N16555;
  assign N4803 = N16514 & N16556;
  assign N4802 = N16514 & N16557;
  assign N4801 = N16514 & N16558;
  assign N4800 = N16514 & N16559;
  assign N4799 = N16514 & N16560;
  assign N4798 = N16514 & N16561;
  assign N4797 = N16514 & N16562;
  assign N4796 = N16514 & N16563;
  assign N4795 = N16514 & N16564;
  assign N4794 = N16514 & N16565;
  assign N4793 = N16514 & N16566;
  assign N4792 = N16514 & N16567;
  assign N4791 = N16514 & N16568;
  assign N4790 = N16514 & N16569;
  assign N4789 = N16514 & N16570;
  assign N4788 = N16515 & N16539;
  assign N4787 = N16515 & N16540;
  assign N4786 = N16515 & N16541;
  assign N4785 = N16515 & N16542;
  assign N4784 = N16515 & N16543;
  assign N4783 = N16515 & N16544;
  assign N4782 = N16515 & N16545;
  assign N4781 = N16515 & N16546;
  assign N4780 = N16515 & N16547;
  assign N4779 = N16515 & N16548;
  assign N4778 = N16515 & N16549;
  assign N4777 = N16515 & N16550;
  assign N4776 = N16515 & N16551;
  assign N4775 = N16515 & N16552;
  assign N4774 = N16515 & N16553;
  assign N4773 = N16515 & N16554;
  assign N4772 = N16515 & N16555;
  assign N4771 = N16515 & N16556;
  assign N4770 = N16515 & N16557;
  assign N4769 = N16515 & N16558;
  assign N4768 = N16515 & N16559;
  assign N4767 = N16515 & N16560;
  assign N4766 = N16515 & N16561;
  assign N4765 = N16515 & N16562;
  assign N4764 = N16515 & N16563;
  assign N4763 = N16515 & N16564;
  assign N4762 = N16515 & N16565;
  assign N4761 = N16515 & N16566;
  assign N4760 = N16515 & N16567;
  assign N4759 = N16515 & N16568;
  assign N4758 = N16515 & N16569;
  assign N4757 = N16515 & N16570;
  assign N4756 = N16516 & N16539;
  assign N4755 = N16516 & N16540;
  assign N4754 = N16516 & N16541;
  assign N4753 = N16516 & N16542;
  assign N4752 = N16516 & N16543;
  assign N4751 = N16516 & N16544;
  assign N4750 = N16516 & N16545;
  assign N4749 = N16516 & N16546;
  assign N4748 = N16516 & N16547;
  assign N4747 = N16516 & N16548;
  assign N4746 = N16516 & N16549;
  assign N4745 = N16516 & N16550;
  assign N4744 = N16516 & N16551;
  assign N4743 = N16516 & N16552;
  assign N4742 = N16516 & N16553;
  assign N4741 = N16516 & N16554;
  assign N4740 = N16516 & N16555;
  assign N4739 = N16516 & N16556;
  assign N4738 = N16516 & N16557;
  assign N4737 = N16516 & N16558;
  assign N4736 = N16516 & N16559;
  assign N4735 = N16516 & N16560;
  assign N4734 = N16516 & N16561;
  assign N4733 = N16516 & N16562;
  assign N4732 = N16516 & N16563;
  assign N4731 = N16516 & N16564;
  assign N4730 = N16516 & N16565;
  assign N4729 = N16516 & N16566;
  assign N4728 = N16516 & N16567;
  assign N4727 = N16516 & N16568;
  assign N4726 = N16516 & N16569;
  assign N4725 = N16516 & N16570;
  assign N4724 = N16517 & N16539;
  assign N4723 = N16517 & N16540;
  assign N4722 = N16517 & N16541;
  assign N4721 = N16517 & N16542;
  assign N4720 = N16517 & N16543;
  assign N4719 = N16517 & N16544;
  assign N4718 = N16517 & N16545;
  assign N4717 = N16517 & N16546;
  assign N4716 = N16517 & N16547;
  assign N4715 = N16517 & N16548;
  assign N4714 = N16517 & N16549;
  assign N4713 = N16517 & N16550;
  assign N4712 = N16517 & N16551;
  assign N4711 = N16517 & N16552;
  assign N4710 = N16517 & N16553;
  assign N4709 = N16517 & N16554;
  assign N4708 = N16517 & N16555;
  assign N4707 = N16517 & N16556;
  assign N4706 = N16517 & N16557;
  assign N4705 = N16517 & N16558;
  assign N4704 = N16517 & N16559;
  assign N4703 = N16517 & N16560;
  assign N4702 = N16517 & N16561;
  assign N4701 = N16517 & N16562;
  assign N4700 = N16517 & N16563;
  assign N4699 = N16517 & N16564;
  assign N4698 = N16517 & N16565;
  assign N4697 = N16517 & N16566;
  assign N4696 = N16517 & N16567;
  assign N4695 = N16517 & N16568;
  assign N4694 = N16517 & N16569;
  assign N4693 = N16517 & N16570;
  assign N4692 = N16518 & N16539;
  assign N4691 = N16518 & N16540;
  assign N4690 = N16518 & N16541;
  assign N4689 = N16518 & N16542;
  assign N4688 = N16518 & N16543;
  assign N4687 = N16518 & N16544;
  assign N4686 = N16518 & N16545;
  assign N4685 = N16518 & N16546;
  assign N4684 = N16518 & N16547;
  assign N4683 = N16518 & N16548;
  assign N4682 = N16518 & N16549;
  assign N4681 = N16518 & N16550;
  assign N4680 = N16518 & N16551;
  assign N4679 = N16518 & N16552;
  assign N4678 = N16518 & N16553;
  assign N4677 = N16518 & N16554;
  assign N4676 = N16518 & N16555;
  assign N4675 = N16518 & N16556;
  assign N4674 = N16518 & N16557;
  assign N4673 = N16518 & N16558;
  assign N4672 = N16518 & N16559;
  assign N4671 = N16518 & N16560;
  assign N4670 = N16518 & N16561;
  assign N4669 = N16518 & N16562;
  assign N4668 = N16518 & N16563;
  assign N4667 = N16518 & N16564;
  assign N4666 = N16518 & N16565;
  assign N4665 = N16518 & N16566;
  assign N4664 = N16518 & N16567;
  assign N4663 = N16518 & N16568;
  assign N4662 = N16518 & N16569;
  assign N4661 = N16518 & N16570;
  assign N4660 = N16519 & N16539;
  assign N4659 = N16519 & N16540;
  assign N4658 = N16519 & N16541;
  assign N4657 = N16519 & N16542;
  assign N4656 = N16519 & N16543;
  assign N4655 = N16519 & N16544;
  assign N4654 = N16519 & N16545;
  assign N4653 = N16519 & N16546;
  assign N4652 = N16519 & N16547;
  assign N4651 = N16519 & N16548;
  assign N4650 = N16519 & N16549;
  assign N4649 = N16519 & N16550;
  assign N4648 = N16519 & N16551;
  assign N4647 = N16519 & N16552;
  assign N4646 = N16519 & N16553;
  assign N4645 = N16519 & N16554;
  assign N4644 = N16519 & N16555;
  assign N4643 = N16519 & N16556;
  assign N4642 = N16519 & N16557;
  assign N4641 = N16519 & N16558;
  assign N4640 = N16519 & N16559;
  assign N4639 = N16519 & N16560;
  assign N4638 = N16519 & N16561;
  assign N4637 = N16519 & N16562;
  assign N4636 = N16519 & N16563;
  assign N4635 = N16519 & N16564;
  assign N4634 = N16519 & N16565;
  assign N4633 = N16519 & N16566;
  assign N4632 = N16519 & N16567;
  assign N4631 = N16519 & N16568;
  assign N4630 = N16519 & N16569;
  assign N4629 = N16519 & N16570;
  assign N4628 = N16520 & N16539;
  assign N4627 = N16520 & N16540;
  assign N4626 = N16520 & N16541;
  assign N4625 = N16520 & N16542;
  assign N4624 = N16520 & N16543;
  assign N4623 = N16520 & N16544;
  assign N4622 = N16520 & N16545;
  assign N4621 = N16520 & N16546;
  assign N4620 = N16520 & N16547;
  assign N4619 = N16520 & N16548;
  assign N4618 = N16520 & N16549;
  assign N4617 = N16520 & N16550;
  assign N4616 = N16520 & N16551;
  assign N4615 = N16520 & N16552;
  assign N4614 = N16520 & N16553;
  assign N4613 = N16520 & N16554;
  assign N4612 = N16520 & N16555;
  assign N4611 = N16520 & N16556;
  assign N4610 = N16520 & N16557;
  assign N4609 = N16520 & N16558;
  assign N4608 = N16520 & N16559;
  assign N4607 = N16520 & N16560;
  assign N4606 = N16520 & N16561;
  assign N4605 = N16520 & N16562;
  assign N4604 = N16520 & N16563;
  assign N4603 = N16520 & N16564;
  assign N4602 = N16520 & N16565;
  assign N4601 = N16520 & N16566;
  assign N4600 = N16520 & N16567;
  assign N4599 = N16520 & N16568;
  assign N4598 = N16520 & N16569;
  assign N4597 = N16520 & N16570;
  assign N4596 = N16521 & N16539;
  assign N4595 = N16521 & N16540;
  assign N4594 = N16521 & N16541;
  assign N4593 = N16521 & N16542;
  assign N4592 = N16521 & N16543;
  assign N4591 = N16521 & N16544;
  assign N4590 = N16521 & N16545;
  assign N4589 = N16521 & N16546;
  assign N4588 = N16521 & N16547;
  assign N4587 = N16521 & N16548;
  assign N4586 = N16521 & N16549;
  assign N4585 = N16521 & N16550;
  assign N4584 = N16521 & N16551;
  assign N4583 = N16521 & N16552;
  assign N4582 = N16521 & N16553;
  assign N4581 = N16521 & N16554;
  assign N4580 = N16521 & N16555;
  assign N4579 = N16521 & N16556;
  assign N4578 = N16521 & N16557;
  assign N4577 = N16521 & N16558;
  assign N4576 = N16521 & N16559;
  assign N4575 = N16521 & N16560;
  assign N4574 = N16521 & N16561;
  assign N4573 = N16521 & N16562;
  assign N4572 = N16521 & N16563;
  assign N4571 = N16521 & N16564;
  assign N4570 = N16521 & N16565;
  assign N4569 = N16521 & N16566;
  assign N4568 = N16521 & N16567;
  assign N4567 = N16521 & N16568;
  assign N4566 = N16521 & N16569;
  assign N4565 = N16521 & N16570;
  assign N16571 = N16498 & N16502;
  assign N16572 = N16498 & N16503;
  assign N16573 = N16498 & N16504;
  assign N16574 = N16498 & N16505;
  assign N16575 = N16499 & N16502;
  assign N16576 = N16499 & N16503;
  assign N16577 = N16499 & N16504;
  assign N16578 = N16499 & N16505;
  assign N16579 = N16500 & N16502;
  assign N16580 = N16500 & N16503;
  assign N16581 = N16500 & N16504;
  assign N16582 = N16500 & N16505;
  assign N16583 = N16501 & N16502;
  assign N16584 = N16501 & N16503;
  assign N16585 = N16501 & N16504;
  assign N16586 = N16501 & N16505;
  assign N10253 = N16571 & N16539;
  assign N10252 = N16571 & N16540;
  assign N10251 = N16571 & N16541;
  assign N10250 = N16571 & N16542;
  assign N10249 = N16571 & N16543;
  assign N10248 = N16571 & N16544;
  assign N10247 = N16571 & N16545;
  assign N10246 = N16571 & N16546;
  assign N10245 = N16571 & N16547;
  assign N10244 = N16571 & N16548;
  assign N10243 = N16571 & N16549;
  assign N10242 = N16571 & N16550;
  assign N10241 = N16571 & N16551;
  assign N10240 = N16571 & N16552;
  assign N10239 = N16571 & N16553;
  assign N10238 = N16571 & N16554;
  assign N10237 = N16571 & N16555;
  assign N10236 = N16571 & N16556;
  assign N10235 = N16571 & N16557;
  assign N10234 = N16571 & N16558;
  assign N10233 = N16571 & N16559;
  assign N10232 = N16571 & N16560;
  assign N10231 = N16571 & N16561;
  assign N10230 = N16571 & N16562;
  assign N10229 = N16571 & N16563;
  assign N10228 = N16571 & N16564;
  assign N10227 = N16571 & N16565;
  assign N10226 = N16571 & N16566;
  assign N10225 = N16571 & N16567;
  assign N10224 = N16571 & N16568;
  assign N10223 = N16571 & N16569;
  assign N10222 = N16571 & N16570;
  assign N10221 = N16572 & N16539;
  assign N10220 = N16572 & N16540;
  assign N10219 = N16572 & N16541;
  assign N10218 = N16572 & N16542;
  assign N10217 = N16572 & N16543;
  assign N10216 = N16572 & N16544;
  assign N10215 = N16572 & N16545;
  assign N10214 = N16572 & N16546;
  assign N10213 = N16572 & N16547;
  assign N10212 = N16572 & N16548;
  assign N10211 = N16572 & N16549;
  assign N10210 = N16572 & N16550;
  assign N10209 = N16572 & N16551;
  assign N10208 = N16572 & N16552;
  assign N10207 = N16572 & N16553;
  assign N10206 = N16572 & N16554;
  assign N10205 = N16572 & N16555;
  assign N10204 = N16572 & N16556;
  assign N10203 = N16572 & N16557;
  assign N10202 = N16572 & N16558;
  assign N10201 = N16572 & N16559;
  assign N10200 = N16572 & N16560;
  assign N10199 = N16572 & N16561;
  assign N10198 = N16572 & N16562;
  assign N10197 = N16572 & N16563;
  assign N10196 = N16572 & N16564;
  assign N10195 = N16572 & N16565;
  assign N10194 = N16572 & N16566;
  assign N10193 = N16572 & N16567;
  assign N10192 = N16572 & N16568;
  assign N10191 = N16572 & N16569;
  assign N10190 = N16572 & N16570;
  assign N10189 = N16573 & N16539;
  assign N10188 = N16573 & N16540;
  assign N10187 = N16573 & N16541;
  assign N10186 = N16573 & N16542;
  assign N10185 = N16573 & N16543;
  assign N10184 = N16573 & N16544;
  assign N10183 = N16573 & N16545;
  assign N10182 = N16573 & N16546;
  assign N10181 = N16573 & N16547;
  assign N10180 = N16573 & N16548;
  assign N10179 = N16573 & N16549;
  assign N10178 = N16573 & N16550;
  assign N10177 = N16573 & N16551;
  assign N10176 = N16573 & N16552;
  assign N10175 = N16573 & N16553;
  assign N10174 = N16573 & N16554;
  assign N10173 = N16573 & N16555;
  assign N10172 = N16573 & N16556;
  assign N10171 = N16573 & N16557;
  assign N10170 = N16573 & N16558;
  assign N10169 = N16573 & N16559;
  assign N10168 = N16573 & N16560;
  assign N10167 = N16573 & N16561;
  assign N10166 = N16573 & N16562;
  assign N10165 = N16573 & N16563;
  assign N10164 = N16573 & N16564;
  assign N10163 = N16573 & N16565;
  assign N10162 = N16573 & N16566;
  assign N10161 = N16573 & N16567;
  assign N10160 = N16573 & N16568;
  assign N10159 = N16573 & N16569;
  assign N10158 = N16573 & N16570;
  assign N10157 = N16574 & N16539;
  assign N10156 = N16574 & N16540;
  assign N10155 = N16574 & N16541;
  assign N10154 = N16574 & N16542;
  assign N10153 = N16574 & N16543;
  assign N10152 = N16574 & N16544;
  assign N10151 = N16574 & N16545;
  assign N10150 = N16574 & N16546;
  assign N10149 = N16574 & N16547;
  assign N10148 = N16574 & N16548;
  assign N10147 = N16574 & N16549;
  assign N10146 = N16574 & N16550;
  assign N10145 = N16574 & N16551;
  assign N10144 = N16574 & N16552;
  assign N10143 = N16574 & N16553;
  assign N10142 = N16574 & N16554;
  assign N10141 = N16574 & N16555;
  assign N10140 = N16574 & N16556;
  assign N10139 = N16574 & N16557;
  assign N10138 = N16574 & N16558;
  assign N10137 = N16574 & N16559;
  assign N10136 = N16574 & N16560;
  assign N10135 = N16574 & N16561;
  assign N10134 = N16574 & N16562;
  assign N10133 = N16574 & N16563;
  assign N10132 = N16574 & N16564;
  assign N10131 = N16574 & N16565;
  assign N10130 = N16574 & N16566;
  assign N10129 = N16574 & N16567;
  assign N10128 = N16574 & N16568;
  assign N10127 = N16574 & N16569;
  assign N10126 = N16574 & N16570;
  assign N10125 = N16575 & N16539;
  assign N10124 = N16575 & N16540;
  assign N10123 = N16575 & N16541;
  assign N10122 = N16575 & N16542;
  assign N10121 = N16575 & N16543;
  assign N10120 = N16575 & N16544;
  assign N10119 = N16575 & N16545;
  assign N10118 = N16575 & N16546;
  assign N10117 = N16575 & N16547;
  assign N10116 = N16575 & N16548;
  assign N10115 = N16575 & N16549;
  assign N10114 = N16575 & N16550;
  assign N10113 = N16575 & N16551;
  assign N10112 = N16575 & N16552;
  assign N10111 = N16575 & N16553;
  assign N10110 = N16575 & N16554;
  assign N10109 = N16575 & N16555;
  assign N10108 = N16575 & N16556;
  assign N10107 = N16575 & N16557;
  assign N10106 = N16575 & N16558;
  assign N10105 = N16575 & N16559;
  assign N10104 = N16575 & N16560;
  assign N10103 = N16575 & N16561;
  assign N10102 = N16575 & N16562;
  assign N10101 = N16575 & N16563;
  assign N10100 = N16575 & N16564;
  assign N10099 = N16575 & N16565;
  assign N10098 = N16575 & N16566;
  assign N10097 = N16575 & N16567;
  assign N10096 = N16575 & N16568;
  assign N10095 = N16575 & N16569;
  assign N10094 = N16575 & N16570;
  assign N10093 = N16576 & N16539;
  assign N10092 = N16576 & N16540;
  assign N10091 = N16576 & N16541;
  assign N10090 = N16576 & N16542;
  assign N10089 = N16576 & N16543;
  assign N10088 = N16576 & N16544;
  assign N10087 = N16576 & N16545;
  assign N10086 = N16576 & N16546;
  assign N10085 = N16576 & N16547;
  assign N10084 = N16576 & N16548;
  assign N10083 = N16576 & N16549;
  assign N10082 = N16576 & N16550;
  assign N10081 = N16576 & N16551;
  assign N10080 = N16576 & N16552;
  assign N10079 = N16576 & N16553;
  assign N10078 = N16576 & N16554;
  assign N10077 = N16576 & N16555;
  assign N10076 = N16576 & N16556;
  assign N10075 = N16576 & N16557;
  assign N10074 = N16576 & N16558;
  assign N10073 = N16576 & N16559;
  assign N10072 = N16576 & N16560;
  assign N10071 = N16576 & N16561;
  assign N10070 = N16576 & N16562;
  assign N10069 = N16576 & N16563;
  assign N10068 = N16576 & N16564;
  assign N10067 = N16576 & N16565;
  assign N10066 = N16576 & N16566;
  assign N10065 = N16576 & N16567;
  assign N10064 = N16576 & N16568;
  assign N10063 = N16576 & N16569;
  assign N10062 = N16576 & N16570;
  assign N10061 = N16577 & N16539;
  assign N10060 = N16577 & N16540;
  assign N10059 = N16577 & N16541;
  assign N10058 = N16577 & N16542;
  assign N10057 = N16577 & N16543;
  assign N10056 = N16577 & N16544;
  assign N10055 = N16577 & N16545;
  assign N10054 = N16577 & N16546;
  assign N10053 = N16577 & N16547;
  assign N10052 = N16577 & N16548;
  assign N10051 = N16577 & N16549;
  assign N10050 = N16577 & N16550;
  assign N10049 = N16577 & N16551;
  assign N10048 = N16577 & N16552;
  assign N10047 = N16577 & N16553;
  assign N10046 = N16577 & N16554;
  assign N10045 = N16577 & N16555;
  assign N10044 = N16577 & N16556;
  assign N10043 = N16577 & N16557;
  assign N10042 = N16577 & N16558;
  assign N10041 = N16577 & N16559;
  assign N10040 = N16577 & N16560;
  assign N10039 = N16577 & N16561;
  assign N10038 = N16577 & N16562;
  assign N10037 = N16577 & N16563;
  assign N10036 = N16577 & N16564;
  assign N10035 = N16577 & N16565;
  assign N10034 = N16577 & N16566;
  assign N10033 = N16577 & N16567;
  assign N10032 = N16577 & N16568;
  assign N10031 = N16577 & N16569;
  assign N10030 = N16577 & N16570;
  assign N10029 = N16578 & N16539;
  assign N10028 = N16578 & N16540;
  assign N10027 = N16578 & N16541;
  assign N10026 = N16578 & N16542;
  assign N10025 = N16578 & N16543;
  assign N10024 = N16578 & N16544;
  assign N10023 = N16578 & N16545;
  assign N10022 = N16578 & N16546;
  assign N10021 = N16578 & N16547;
  assign N10020 = N16578 & N16548;
  assign N10019 = N16578 & N16549;
  assign N10018 = N16578 & N16550;
  assign N10017 = N16578 & N16551;
  assign N10016 = N16578 & N16552;
  assign N10015 = N16578 & N16553;
  assign N10014 = N16578 & N16554;
  assign N10013 = N16578 & N16555;
  assign N10012 = N16578 & N16556;
  assign N10011 = N16578 & N16557;
  assign N10010 = N16578 & N16558;
  assign N10009 = N16578 & N16559;
  assign N10008 = N16578 & N16560;
  assign N10007 = N16578 & N16561;
  assign N10006 = N16578 & N16562;
  assign N10005 = N16578 & N16563;
  assign N10004 = N16578 & N16564;
  assign N10003 = N16578 & N16565;
  assign N10002 = N16578 & N16566;
  assign N10001 = N16578 & N16567;
  assign N10000 = N16578 & N16568;
  assign N9999 = N16578 & N16569;
  assign N9998 = N16578 & N16570;
  assign N9997 = N16579 & N16539;
  assign N9996 = N16579 & N16540;
  assign N9995 = N16579 & N16541;
  assign N9994 = N16579 & N16542;
  assign N9993 = N16579 & N16543;
  assign N9992 = N16579 & N16544;
  assign N9991 = N16579 & N16545;
  assign N9990 = N16579 & N16546;
  assign N9989 = N16579 & N16547;
  assign N9988 = N16579 & N16548;
  assign N9987 = N16579 & N16549;
  assign N9986 = N16579 & N16550;
  assign N9985 = N16579 & N16551;
  assign N9984 = N16579 & N16552;
  assign N9983 = N16579 & N16553;
  assign N9982 = N16579 & N16554;
  assign N9981 = N16579 & N16555;
  assign N9980 = N16579 & N16556;
  assign N9979 = N16579 & N16557;
  assign N9978 = N16579 & N16558;
  assign N9977 = N16579 & N16559;
  assign N9976 = N16579 & N16560;
  assign N9975 = N16579 & N16561;
  assign N9974 = N16579 & N16562;
  assign N9973 = N16579 & N16563;
  assign N9972 = N16579 & N16564;
  assign N9971 = N16579 & N16565;
  assign N9970 = N16579 & N16566;
  assign N9969 = N16579 & N16567;
  assign N9968 = N16579 & N16568;
  assign N9967 = N16579 & N16569;
  assign N9966 = N16579 & N16570;
  assign N9965 = N16580 & N16539;
  assign N9964 = N16580 & N16540;
  assign N9963 = N16580 & N16541;
  assign N9962 = N16580 & N16542;
  assign N9961 = N16580 & N16543;
  assign N9960 = N16580 & N16544;
  assign N9959 = N16580 & N16545;
  assign N9958 = N16580 & N16546;
  assign N9957 = N16580 & N16547;
  assign N9956 = N16580 & N16548;
  assign N9955 = N16580 & N16549;
  assign N9954 = N16580 & N16550;
  assign N9953 = N16580 & N16551;
  assign N9952 = N16580 & N16552;
  assign N9951 = N16580 & N16553;
  assign N9950 = N16580 & N16554;
  assign N9949 = N16580 & N16555;
  assign N9948 = N16580 & N16556;
  assign N9947 = N16580 & N16557;
  assign N9946 = N16580 & N16558;
  assign N9945 = N16580 & N16559;
  assign N9944 = N16580 & N16560;
  assign N9943 = N16580 & N16561;
  assign N9942 = N16580 & N16562;
  assign N9941 = N16580 & N16563;
  assign N9940 = N16580 & N16564;
  assign N9939 = N16580 & N16565;
  assign N9938 = N16580 & N16566;
  assign N9937 = N16580 & N16567;
  assign N9936 = N16580 & N16568;
  assign N9935 = N16580 & N16569;
  assign N9934 = N16580 & N16570;
  assign N9933 = N16581 & N16539;
  assign N9932 = N16581 & N16540;
  assign N9931 = N16581 & N16541;
  assign N9930 = N16581 & N16542;
  assign N9929 = N16581 & N16543;
  assign N9928 = N16581 & N16544;
  assign N9927 = N16581 & N16545;
  assign N9926 = N16581 & N16546;
  assign N9925 = N16581 & N16547;
  assign N9924 = N16581 & N16548;
  assign N9923 = N16581 & N16549;
  assign N9922 = N16581 & N16550;
  assign N9921 = N16581 & N16551;
  assign N9920 = N16581 & N16552;
  assign N9919 = N16581 & N16553;
  assign N9918 = N16581 & N16554;
  assign N9917 = N16581 & N16555;
  assign N9916 = N16581 & N16556;
  assign N9915 = N16581 & N16557;
  assign N9914 = N16581 & N16558;
  assign N9913 = N16581 & N16559;
  assign N9912 = N16581 & N16560;
  assign N9911 = N16581 & N16561;
  assign N9910 = N16581 & N16562;
  assign N9909 = N16581 & N16563;
  assign N9908 = N16581 & N16564;
  assign N9907 = N16581 & N16565;
  assign N9906 = N16581 & N16566;
  assign N9905 = N16581 & N16567;
  assign N9904 = N16581 & N16568;
  assign N9903 = N16581 & N16569;
  assign N9902 = N16581 & N16570;
  assign N9901 = N16582 & N16539;
  assign N9900 = N16582 & N16540;
  assign N9899 = N16582 & N16541;
  assign N9898 = N16582 & N16542;
  assign N9897 = N16582 & N16543;
  assign N9896 = N16582 & N16544;
  assign N9895 = N16582 & N16545;
  assign N9894 = N16582 & N16546;
  assign N9893 = N16582 & N16547;
  assign N9892 = N16582 & N16548;
  assign N9891 = N16582 & N16549;
  assign N9890 = N16582 & N16550;
  assign N9889 = N16582 & N16551;
  assign N9888 = N16582 & N16552;
  assign N9887 = N16582 & N16553;
  assign N9886 = N16582 & N16554;
  assign N9885 = N16582 & N16555;
  assign N9884 = N16582 & N16556;
  assign N9883 = N16582 & N16557;
  assign N9882 = N16582 & N16558;
  assign N9881 = N16582 & N16559;
  assign N9880 = N16582 & N16560;
  assign N9879 = N16582 & N16561;
  assign N9878 = N16582 & N16562;
  assign N9877 = N16582 & N16563;
  assign N9876 = N16582 & N16564;
  assign N9875 = N16582 & N16565;
  assign N9874 = N16582 & N16566;
  assign N9873 = N16582 & N16567;
  assign N9872 = N16582 & N16568;
  assign N9871 = N16582 & N16569;
  assign N9870 = N16582 & N16570;
  assign N9869 = N16583 & N16539;
  assign N9868 = N16583 & N16540;
  assign N9867 = N16583 & N16541;
  assign N9866 = N16583 & N16542;
  assign N9865 = N16583 & N16543;
  assign N9864 = N16583 & N16544;
  assign N9863 = N16583 & N16545;
  assign N9862 = N16583 & N16546;
  assign N9861 = N16583 & N16547;
  assign N9860 = N16583 & N16548;
  assign N9859 = N16583 & N16549;
  assign N9858 = N16583 & N16550;
  assign N9857 = N16583 & N16551;
  assign N9856 = N16583 & N16552;
  assign N9855 = N16583 & N16553;
  assign N9854 = N16583 & N16554;
  assign N9853 = N16583 & N16555;
  assign N9852 = N16583 & N16556;
  assign N9851 = N16583 & N16557;
  assign N9850 = N16583 & N16558;
  assign N9849 = N16583 & N16559;
  assign N9848 = N16583 & N16560;
  assign N9847 = N16583 & N16561;
  assign N9846 = N16583 & N16562;
  assign N9845 = N16583 & N16563;
  assign N9844 = N16583 & N16564;
  assign N9843 = N16583 & N16565;
  assign N9842 = N16583 & N16566;
  assign N9841 = N16583 & N16567;
  assign N9840 = N16583 & N16568;
  assign N9839 = N16583 & N16569;
  assign N9838 = N16583 & N16570;
  assign N9837 = N16584 & N16539;
  assign N9836 = N16584 & N16540;
  assign N9835 = N16584 & N16541;
  assign N9834 = N16584 & N16542;
  assign N9833 = N16584 & N16543;
  assign N9832 = N16584 & N16544;
  assign N9831 = N16584 & N16545;
  assign N9830 = N16584 & N16546;
  assign N9829 = N16584 & N16547;
  assign N9828 = N16584 & N16548;
  assign N9827 = N16584 & N16549;
  assign N9826 = N16584 & N16550;
  assign N9825 = N16584 & N16551;
  assign N9824 = N16584 & N16552;
  assign N9823 = N16584 & N16553;
  assign N9822 = N16584 & N16554;
  assign N9821 = N16584 & N16555;
  assign N9820 = N16584 & N16556;
  assign N9819 = N16584 & N16557;
  assign N9818 = N16584 & N16558;
  assign N9817 = N16584 & N16559;
  assign N9816 = N16584 & N16560;
  assign N9815 = N16584 & N16561;
  assign N9814 = N16584 & N16562;
  assign N9813 = N16584 & N16563;
  assign N9812 = N16584 & N16564;
  assign N9811 = N16584 & N16565;
  assign N9810 = N16584 & N16566;
  assign N9809 = N16584 & N16567;
  assign N9808 = N16584 & N16568;
  assign N9807 = N16584 & N16569;
  assign N9806 = N16584 & N16570;
  assign N9805 = N16585 & N16539;
  assign N9804 = N16585 & N16540;
  assign N9803 = N16585 & N16541;
  assign N9802 = N16585 & N16542;
  assign N9801 = N16585 & N16543;
  assign N9800 = N16585 & N16544;
  assign N9799 = N16585 & N16545;
  assign N9798 = N16585 & N16546;
  assign N9797 = N16585 & N16547;
  assign N9796 = N16585 & N16548;
  assign N9795 = N16585 & N16549;
  assign N9794 = N16585 & N16550;
  assign N9793 = N16585 & N16551;
  assign N9792 = N16585 & N16552;
  assign N9791 = N16585 & N16553;
  assign N9790 = N16585 & N16554;
  assign N9789 = N16585 & N16555;
  assign N9788 = N16585 & N16556;
  assign N9787 = N16585 & N16557;
  assign N9786 = N16585 & N16558;
  assign N9785 = N16585 & N16559;
  assign N9784 = N16585 & N16560;
  assign N9783 = N16585 & N16561;
  assign N9782 = N16585 & N16562;
  assign N9781 = N16585 & N16563;
  assign N9780 = N16585 & N16564;
  assign N9779 = N16585 & N16565;
  assign N9778 = N16585 & N16566;
  assign N9777 = N16585 & N16567;
  assign N9776 = N16585 & N16568;
  assign N9775 = N16585 & N16569;
  assign N9774 = N16585 & N16570;
  assign N9773 = N16586 & N16539;
  assign N9772 = N16586 & N16540;
  assign N9771 = N16586 & N16541;
  assign N9770 = N16586 & N16542;
  assign N9769 = N16586 & N16543;
  assign N9768 = N16586 & N16544;
  assign N9767 = N16586 & N16545;
  assign N9766 = N16586 & N16546;
  assign N9765 = N16586 & N16547;
  assign N9764 = N16586 & N16548;
  assign N9763 = N16586 & N16549;
  assign N9762 = N16586 & N16550;
  assign N9761 = N16586 & N16551;
  assign N9760 = N16586 & N16552;
  assign N9759 = N16586 & N16553;
  assign N9758 = N16586 & N16554;
  assign N9757 = N16586 & N16555;
  assign N9756 = N16586 & N16556;
  assign N9755 = N16586 & N16557;
  assign N9754 = N16586 & N16558;
  assign N9753 = N16586 & N16559;
  assign N9752 = N16586 & N16560;
  assign N9751 = N16586 & N16561;
  assign N9750 = N16586 & N16562;
  assign N9749 = N16586 & N16563;
  assign N9748 = N16586 & N16564;
  assign N9747 = N16586 & N16565;
  assign N9746 = N16586 & N16566;
  assign N9745 = N16586 & N16567;
  assign N9744 = N16586 & N16568;
  assign N9743 = N16586 & N16569;
  assign N9742 = N16586 & N16570;
  assign N16587 = N16498 & N16502;
  assign N16588 = N16498 & N16503;
  assign N16589 = N16498 & N16504;
  assign N16590 = N16498 & N16505;
  assign N16591 = N16499 & N16502;
  assign N16592 = N16499 & N16503;
  assign N16593 = N16499 & N16504;
  assign N16594 = N16499 & N16505;
  assign N16595 = N16500 & N16502;
  assign N16596 = N16500 & N16503;
  assign N16597 = N16500 & N16504;
  assign N16598 = N16500 & N16505;
  assign N16599 = N16501 & N16502;
  assign N16600 = N16501 & N16503;
  assign N16601 = N16501 & N16504;
  assign N16602 = N16501 & N16505;
  assign N16603 = N16522 & N16531;
  assign N16604 = N16522 & N16532;
  assign N16605 = N16522 & N16533;
  assign N16606 = N16522 & N16534;
  assign N16607 = N16522 & N16535;
  assign N16608 = N16522 & N16536;
  assign N16609 = N16522 & N16537;
  assign N16610 = N16522 & N16538;
  assign N16611 = N16523 & N16531;
  assign N16612 = N16523 & N16532;
  assign N16613 = N16523 & N16533;
  assign N16614 = N16523 & N16534;
  assign N16615 = N16523 & N16535;
  assign N16616 = N16523 & N16536;
  assign N16617 = N16523 & N16537;
  assign N16618 = N16523 & N16538;
  assign N16619 = N16524 & N16531;
  assign N16620 = N16524 & N16532;
  assign N16621 = N16524 & N16533;
  assign N16622 = N16524 & N16534;
  assign N16623 = N16524 & N16535;
  assign N16624 = N16524 & N16536;
  assign N16625 = N16524 & N16537;
  assign N16626 = N16524 & N16538;
  assign N16627 = N16525 & N16531;
  assign N16628 = N16525 & N16532;
  assign N16629 = N16525 & N16533;
  assign N16630 = N16525 & N16534;
  assign N16631 = N16525 & N16535;
  assign N16632 = N16525 & N16536;
  assign N16633 = N16525 & N16537;
  assign N16634 = N16525 & N16538;
  assign N14036 = N16587 & N16603;
  assign N14035 = N16587 & N16604;
  assign N14034 = N16587 & N16605;
  assign N14033 = N16587 & N16606;
  assign N14032 = N16587 & N16607;
  assign N14031 = N16587 & N16608;
  assign N14030 = N16587 & N16609;
  assign N14029 = N16587 & N16610;
  assign N14028 = N16587 & N16611;
  assign N14027 = N16587 & N16612;
  assign N14026 = N16587 & N16613;
  assign N14025 = N16587 & N16614;
  assign N14024 = N16587 & N16615;
  assign N14023 = N16587 & N16616;
  assign N14022 = N16587 & N16617;
  assign N14021 = N16587 & N16618;
  assign N14020 = N16587 & N16619;
  assign N14019 = N16587 & N16620;
  assign N14018 = N16587 & N16621;
  assign N14017 = N16587 & N16622;
  assign N14016 = N16587 & N16623;
  assign N14015 = N16587 & N16624;
  assign N14014 = N16587 & N16625;
  assign N14013 = N16587 & N16626;
  assign N14012 = N16587 & N16627;
  assign N14011 = N16587 & N16628;
  assign N14010 = N16587 & N16629;
  assign N14009 = N16587 & N16630;
  assign N14008 = N16587 & N16631;
  assign N14007 = N16587 & N16632;
  assign N14006 = N16587 & N16633;
  assign N14005 = N16587 & N16634;
  assign N14004 = N16588 & N16603;
  assign N14003 = N16588 & N16604;
  assign N14002 = N16588 & N16605;
  assign N14001 = N16588 & N16606;
  assign N14000 = N16588 & N16607;
  assign N13999 = N16588 & N16608;
  assign N13998 = N16588 & N16609;
  assign N13997 = N16588 & N16610;
  assign N13996 = N16588 & N16611;
  assign N13995 = N16588 & N16612;
  assign N13994 = N16588 & N16613;
  assign N13993 = N16588 & N16614;
  assign N13992 = N16588 & N16615;
  assign N13991 = N16588 & N16616;
  assign N13990 = N16588 & N16617;
  assign N13989 = N16588 & N16618;
  assign N13988 = N16588 & N16619;
  assign N13987 = N16588 & N16620;
  assign N13986 = N16588 & N16621;
  assign N13985 = N16588 & N16622;
  assign N13984 = N16588 & N16623;
  assign N13983 = N16588 & N16624;
  assign N13982 = N16588 & N16625;
  assign N13981 = N16588 & N16626;
  assign N13980 = N16588 & N16627;
  assign N13979 = N16588 & N16628;
  assign N13978 = N16588 & N16629;
  assign N13977 = N16588 & N16630;
  assign N13976 = N16588 & N16631;
  assign N13975 = N16588 & N16632;
  assign N13974 = N16588 & N16633;
  assign N13973 = N16588 & N16634;
  assign N13972 = N16589 & N16603;
  assign N13971 = N16589 & N16604;
  assign N13970 = N16589 & N16605;
  assign N13969 = N16589 & N16606;
  assign N13968 = N16589 & N16607;
  assign N13967 = N16589 & N16608;
  assign N13966 = N16589 & N16609;
  assign N13965 = N16589 & N16610;
  assign N13964 = N16589 & N16611;
  assign N13963 = N16589 & N16612;
  assign N13962 = N16589 & N16613;
  assign N13961 = N16589 & N16614;
  assign N13960 = N16589 & N16615;
  assign N13959 = N16589 & N16616;
  assign N13958 = N16589 & N16617;
  assign N13957 = N16589 & N16618;
  assign N13956 = N16589 & N16619;
  assign N13955 = N16589 & N16620;
  assign N13954 = N16589 & N16621;
  assign N13953 = N16589 & N16622;
  assign N13952 = N16589 & N16623;
  assign N13951 = N16589 & N16624;
  assign N13950 = N16589 & N16625;
  assign N13949 = N16589 & N16626;
  assign N13948 = N16589 & N16627;
  assign N13947 = N16589 & N16628;
  assign N13946 = N16589 & N16629;
  assign N13945 = N16589 & N16630;
  assign N13944 = N16589 & N16631;
  assign N13943 = N16589 & N16632;
  assign N13942 = N16589 & N16633;
  assign N13941 = N16589 & N16634;
  assign N13940 = N16590 & N16603;
  assign N13939 = N16590 & N16604;
  assign N13938 = N16590 & N16605;
  assign N13937 = N16590 & N16606;
  assign N13936 = N16590 & N16607;
  assign N13935 = N16590 & N16608;
  assign N13934 = N16590 & N16609;
  assign N13933 = N16590 & N16610;
  assign N13932 = N16590 & N16611;
  assign N13931 = N16590 & N16612;
  assign N13930 = N16590 & N16613;
  assign N13929 = N16590 & N16614;
  assign N13928 = N16590 & N16615;
  assign N13927 = N16590 & N16616;
  assign N13926 = N16590 & N16617;
  assign N13925 = N16590 & N16618;
  assign N13924 = N16590 & N16619;
  assign N13923 = N16590 & N16620;
  assign N13922 = N16590 & N16621;
  assign N13921 = N16590 & N16622;
  assign N13920 = N16590 & N16623;
  assign N13919 = N16590 & N16624;
  assign N13918 = N16590 & N16625;
  assign N13917 = N16590 & N16626;
  assign N13916 = N16590 & N16627;
  assign N13915 = N16590 & N16628;
  assign N13914 = N16590 & N16629;
  assign N13913 = N16590 & N16630;
  assign N13912 = N16590 & N16631;
  assign N13911 = N16590 & N16632;
  assign N13910 = N16590 & N16633;
  assign N13909 = N16590 & N16634;
  assign N13908 = N16591 & N16603;
  assign N13907 = N16591 & N16604;
  assign N13906 = N16591 & N16605;
  assign N13905 = N16591 & N16606;
  assign N13904 = N16591 & N16607;
  assign N13903 = N16591 & N16608;
  assign N13902 = N16591 & N16609;
  assign N13901 = N16591 & N16610;
  assign N13900 = N16591 & N16611;
  assign N13899 = N16591 & N16612;
  assign N13898 = N16591 & N16613;
  assign N13897 = N16591 & N16614;
  assign N13896 = N16591 & N16615;
  assign N13895 = N16591 & N16616;
  assign N13894 = N16591 & N16617;
  assign N13893 = N16591 & N16618;
  assign N13892 = N16591 & N16619;
  assign N13891 = N16591 & N16620;
  assign N13890 = N16591 & N16621;
  assign N13889 = N16591 & N16622;
  assign N13888 = N16591 & N16623;
  assign N13887 = N16591 & N16624;
  assign N13886 = N16591 & N16625;
  assign N13885 = N16591 & N16626;
  assign N13884 = N16591 & N16627;
  assign N13883 = N16591 & N16628;
  assign N13882 = N16591 & N16629;
  assign N13881 = N16591 & N16630;
  assign N13880 = N16591 & N16631;
  assign N13879 = N16591 & N16632;
  assign N13878 = N16591 & N16633;
  assign N13877 = N16591 & N16634;
  assign N13876 = N16592 & N16603;
  assign N13875 = N16592 & N16604;
  assign N13874 = N16592 & N16605;
  assign N13873 = N16592 & N16606;
  assign N13872 = N16592 & N16607;
  assign N13871 = N16592 & N16608;
  assign N13870 = N16592 & N16609;
  assign N13869 = N16592 & N16610;
  assign N13868 = N16592 & N16611;
  assign N13867 = N16592 & N16612;
  assign N13866 = N16592 & N16613;
  assign N13865 = N16592 & N16614;
  assign N13864 = N16592 & N16615;
  assign N13863 = N16592 & N16616;
  assign N13862 = N16592 & N16617;
  assign N13861 = N16592 & N16618;
  assign N13860 = N16592 & N16619;
  assign N13859 = N16592 & N16620;
  assign N13858 = N16592 & N16621;
  assign N13857 = N16592 & N16622;
  assign N13856 = N16592 & N16623;
  assign N13855 = N16592 & N16624;
  assign N13854 = N16592 & N16625;
  assign N13853 = N16592 & N16626;
  assign N13852 = N16592 & N16627;
  assign N13851 = N16592 & N16628;
  assign N13850 = N16592 & N16629;
  assign N13849 = N16592 & N16630;
  assign N13848 = N16592 & N16631;
  assign N13847 = N16592 & N16632;
  assign N13846 = N16592 & N16633;
  assign N13845 = N16592 & N16634;
  assign N13844 = N16593 & N16603;
  assign N13843 = N16593 & N16604;
  assign N13842 = N16593 & N16605;
  assign N13841 = N16593 & N16606;
  assign N13840 = N16593 & N16607;
  assign N13839 = N16593 & N16608;
  assign N13838 = N16593 & N16609;
  assign N13837 = N16593 & N16610;
  assign N13836 = N16593 & N16611;
  assign N13835 = N16593 & N16612;
  assign N13834 = N16593 & N16613;
  assign N13833 = N16593 & N16614;
  assign N13832 = N16593 & N16615;
  assign N13831 = N16593 & N16616;
  assign N13830 = N16593 & N16617;
  assign N13829 = N16593 & N16618;
  assign N13828 = N16593 & N16619;
  assign N13827 = N16593 & N16620;
  assign N13826 = N16593 & N16621;
  assign N13825 = N16593 & N16622;
  assign N13824 = N16593 & N16623;
  assign N13823 = N16593 & N16624;
  assign N13822 = N16593 & N16625;
  assign N13821 = N16593 & N16626;
  assign N13820 = N16593 & N16627;
  assign N13819 = N16593 & N16628;
  assign N13818 = N16593 & N16629;
  assign N13817 = N16593 & N16630;
  assign N13816 = N16593 & N16631;
  assign N13815 = N16593 & N16632;
  assign N13814 = N16593 & N16633;
  assign N13813 = N16593 & N16634;
  assign N13812 = N16594 & N16603;
  assign N13811 = N16594 & N16604;
  assign N13810 = N16594 & N16605;
  assign N13809 = N16594 & N16606;
  assign N13808 = N16594 & N16607;
  assign N13807 = N16594 & N16608;
  assign N13806 = N16594 & N16609;
  assign N13805 = N16594 & N16610;
  assign N13804 = N16594 & N16611;
  assign N13803 = N16594 & N16612;
  assign N13802 = N16594 & N16613;
  assign N13801 = N16594 & N16614;
  assign N13800 = N16594 & N16615;
  assign N13799 = N16594 & N16616;
  assign N13798 = N16594 & N16617;
  assign N13797 = N16594 & N16618;
  assign N13796 = N16594 & N16619;
  assign N13795 = N16594 & N16620;
  assign N13794 = N16594 & N16621;
  assign N13793 = N16594 & N16622;
  assign N13792 = N16594 & N16623;
  assign N13791 = N16594 & N16624;
  assign N13790 = N16594 & N16625;
  assign N13789 = N16594 & N16626;
  assign N13788 = N16594 & N16627;
  assign N13787 = N16594 & N16628;
  assign N13786 = N16594 & N16629;
  assign N13785 = N16594 & N16630;
  assign N13784 = N16594 & N16631;
  assign N13783 = N16594 & N16632;
  assign N13782 = N16594 & N16633;
  assign N13781 = N16594 & N16634;
  assign N13780 = N16595 & N16603;
  assign N13779 = N16595 & N16604;
  assign N13778 = N16595 & N16605;
  assign N13777 = N16595 & N16606;
  assign N13776 = N16595 & N16607;
  assign N13775 = N16595 & N16608;
  assign N13774 = N16595 & N16609;
  assign N13773 = N16595 & N16610;
  assign N13772 = N16595 & N16611;
  assign N13771 = N16595 & N16612;
  assign N13770 = N16595 & N16613;
  assign N13769 = N16595 & N16614;
  assign N13768 = N16595 & N16615;
  assign N13767 = N16595 & N16616;
  assign N13766 = N16595 & N16617;
  assign N13765 = N16595 & N16618;
  assign N13764 = N16595 & N16619;
  assign N13763 = N16595 & N16620;
  assign N13762 = N16595 & N16621;
  assign N13761 = N16595 & N16622;
  assign N13760 = N16595 & N16623;
  assign N13759 = N16595 & N16624;
  assign N13758 = N16595 & N16625;
  assign N13757 = N16595 & N16626;
  assign N13756 = N16595 & N16627;
  assign N13755 = N16595 & N16628;
  assign N13754 = N16595 & N16629;
  assign N13753 = N16595 & N16630;
  assign N13752 = N16595 & N16631;
  assign N13751 = N16595 & N16632;
  assign N13750 = N16595 & N16633;
  assign N13749 = N16595 & N16634;
  assign N13748 = N16596 & N16603;
  assign N13747 = N16596 & N16604;
  assign N13746 = N16596 & N16605;
  assign N13745 = N16596 & N16606;
  assign N13744 = N16596 & N16607;
  assign N13743 = N16596 & N16608;
  assign N13742 = N16596 & N16609;
  assign N13741 = N16596 & N16610;
  assign N13740 = N16596 & N16611;
  assign N13739 = N16596 & N16612;
  assign N13738 = N16596 & N16613;
  assign N13737 = N16596 & N16614;
  assign N13736 = N16596 & N16615;
  assign N13735 = N16596 & N16616;
  assign N13734 = N16596 & N16617;
  assign N13733 = N16596 & N16618;
  assign N13732 = N16596 & N16619;
  assign N13731 = N16596 & N16620;
  assign N13730 = N16596 & N16621;
  assign N13729 = N16596 & N16622;
  assign N13728 = N16596 & N16623;
  assign N13727 = N16596 & N16624;
  assign N13726 = N16596 & N16625;
  assign N13725 = N16596 & N16626;
  assign N13724 = N16596 & N16627;
  assign N13723 = N16596 & N16628;
  assign N13722 = N16596 & N16629;
  assign N13721 = N16596 & N16630;
  assign N13720 = N16596 & N16631;
  assign N13719 = N16596 & N16632;
  assign N13718 = N16596 & N16633;
  assign N13717 = N16596 & N16634;
  assign N13716 = N16597 & N16603;
  assign N13715 = N16597 & N16604;
  assign N13714 = N16597 & N16605;
  assign N13713 = N16597 & N16606;
  assign N13712 = N16597 & N16607;
  assign N13711 = N16597 & N16608;
  assign N13710 = N16597 & N16609;
  assign N13709 = N16597 & N16610;
  assign N13708 = N16597 & N16611;
  assign N13707 = N16597 & N16612;
  assign N13706 = N16597 & N16613;
  assign N13705 = N16597 & N16614;
  assign N13704 = N16597 & N16615;
  assign N13703 = N16597 & N16616;
  assign N13702 = N16597 & N16617;
  assign N13701 = N16597 & N16618;
  assign N13700 = N16597 & N16619;
  assign N13699 = N16597 & N16620;
  assign N13698 = N16597 & N16621;
  assign N13697 = N16597 & N16622;
  assign N13696 = N16597 & N16623;
  assign N13695 = N16597 & N16624;
  assign N13694 = N16597 & N16625;
  assign N13693 = N16597 & N16626;
  assign N13692 = N16597 & N16627;
  assign N13691 = N16597 & N16628;
  assign N13690 = N16597 & N16629;
  assign N13689 = N16597 & N16630;
  assign N13688 = N16597 & N16631;
  assign N13687 = N16597 & N16632;
  assign N13686 = N16597 & N16633;
  assign N13685 = N16597 & N16634;
  assign N13684 = N16598 & N16603;
  assign N13683 = N16598 & N16604;
  assign N13682 = N16598 & N16605;
  assign N13681 = N16598 & N16606;
  assign N13680 = N16598 & N16607;
  assign N13679 = N16598 & N16608;
  assign N13678 = N16598 & N16609;
  assign N13677 = N16598 & N16610;
  assign N13676 = N16598 & N16611;
  assign N13675 = N16598 & N16612;
  assign N13674 = N16598 & N16613;
  assign N13673 = N16598 & N16614;
  assign N13672 = N16598 & N16615;
  assign N13671 = N16598 & N16616;
  assign N13670 = N16598 & N16617;
  assign N13669 = N16598 & N16618;
  assign N13668 = N16598 & N16619;
  assign N13667 = N16598 & N16620;
  assign N13666 = N16598 & N16621;
  assign N13665 = N16598 & N16622;
  assign N13664 = N16598 & N16623;
  assign N13663 = N16598 & N16624;
  assign N13662 = N16598 & N16625;
  assign N13661 = N16598 & N16626;
  assign N13660 = N16598 & N16627;
  assign N13659 = N16598 & N16628;
  assign N13658 = N16598 & N16629;
  assign N13657 = N16598 & N16630;
  assign N13656 = N16598 & N16631;
  assign N13655 = N16598 & N16632;
  assign N13654 = N16598 & N16633;
  assign N13653 = N16598 & N16634;
  assign N13652 = N16599 & N16603;
  assign N13651 = N16599 & N16604;
  assign N13650 = N16599 & N16605;
  assign N13649 = N16599 & N16606;
  assign N13648 = N16599 & N16607;
  assign N13647 = N16599 & N16608;
  assign N13646 = N16599 & N16609;
  assign N13645 = N16599 & N16610;
  assign N13644 = N16599 & N16611;
  assign N13643 = N16599 & N16612;
  assign N13642 = N16599 & N16613;
  assign N13641 = N16599 & N16614;
  assign N13640 = N16599 & N16615;
  assign N13639 = N16599 & N16616;
  assign N13638 = N16599 & N16617;
  assign N13637 = N16599 & N16618;
  assign N13636 = N16599 & N16619;
  assign N13635 = N16599 & N16620;
  assign N13634 = N16599 & N16621;
  assign N13633 = N16599 & N16622;
  assign N13632 = N16599 & N16623;
  assign N13631 = N16599 & N16624;
  assign N13630 = N16599 & N16625;
  assign N13629 = N16599 & N16626;
  assign N13628 = N16599 & N16627;
  assign N13627 = N16599 & N16628;
  assign N13626 = N16599 & N16629;
  assign N13625 = N16599 & N16630;
  assign N13624 = N16599 & N16631;
  assign N13623 = N16599 & N16632;
  assign N13622 = N16599 & N16633;
  assign N13621 = N16599 & N16634;
  assign N13620 = N16600 & N16603;
  assign N13619 = N16600 & N16604;
  assign N13618 = N16600 & N16605;
  assign N13617 = N16600 & N16606;
  assign N13616 = N16600 & N16607;
  assign N13615 = N16600 & N16608;
  assign N13614 = N16600 & N16609;
  assign N13613 = N16600 & N16610;
  assign N13612 = N16600 & N16611;
  assign N13611 = N16600 & N16612;
  assign N13610 = N16600 & N16613;
  assign N13609 = N16600 & N16614;
  assign N13608 = N16600 & N16615;
  assign N13607 = N16600 & N16616;
  assign N13606 = N16600 & N16617;
  assign N13605 = N16600 & N16618;
  assign N13604 = N16600 & N16619;
  assign N13603 = N16600 & N16620;
  assign N13602 = N16600 & N16621;
  assign N13601 = N16600 & N16622;
  assign N13600 = N16600 & N16623;
  assign N13599 = N16600 & N16624;
  assign N13598 = N16600 & N16625;
  assign N13597 = N16600 & N16626;
  assign N13596 = N16600 & N16627;
  assign N13595 = N16600 & N16628;
  assign N13594 = N16600 & N16629;
  assign N13593 = N16600 & N16630;
  assign N13592 = N16600 & N16631;
  assign N13591 = N16600 & N16632;
  assign N13590 = N16600 & N16633;
  assign N13589 = N16600 & N16634;
  assign N13588 = N16601 & N16603;
  assign N13587 = N16601 & N16604;
  assign N13586 = N16601 & N16605;
  assign N13585 = N16601 & N16606;
  assign N13584 = N16601 & N16607;
  assign N13583 = N16601 & N16608;
  assign N13582 = N16601 & N16609;
  assign N13581 = N16601 & N16610;
  assign N13580 = N16601 & N16611;
  assign N13579 = N16601 & N16612;
  assign N13578 = N16601 & N16613;
  assign N13577 = N16601 & N16614;
  assign N13576 = N16601 & N16615;
  assign N13575 = N16601 & N16616;
  assign N13574 = N16601 & N16617;
  assign N13573 = N16601 & N16618;
  assign N13572 = N16601 & N16619;
  assign N13571 = N16601 & N16620;
  assign N13570 = N16601 & N16621;
  assign N13569 = N16601 & N16622;
  assign N13568 = N16601 & N16623;
  assign N13567 = N16601 & N16624;
  assign N13566 = N16601 & N16625;
  assign N13565 = N16601 & N16626;
  assign N13564 = N16601 & N16627;
  assign N13563 = N16601 & N16628;
  assign N13562 = N16601 & N16629;
  assign N13561 = N16601 & N16630;
  assign N13560 = N16601 & N16631;
  assign N13559 = N16601 & N16632;
  assign N13558 = N16601 & N16633;
  assign N13557 = N16601 & N16634;
  assign N13556 = N16602 & N16603;
  assign N13555 = N16602 & N16604;
  assign N13554 = N16602 & N16605;
  assign N13553 = N16602 & N16606;
  assign N13552 = N16602 & N16607;
  assign N13551 = N16602 & N16608;
  assign N13550 = N16602 & N16609;
  assign N13549 = N16602 & N16610;
  assign N13548 = N16602 & N16611;
  assign N13547 = N16602 & N16612;
  assign N13546 = N16602 & N16613;
  assign N13545 = N16602 & N16614;
  assign N13544 = N16602 & N16615;
  assign N13543 = N16602 & N16616;
  assign N13542 = N16602 & N16617;
  assign N13541 = N16602 & N16618;
  assign N13540 = N16602 & N16619;
  assign N13539 = N16602 & N16620;
  assign N13538 = N16602 & N16621;
  assign N13537 = N16602 & N16622;
  assign N13536 = N16602 & N16623;
  assign N13535 = N16602 & N16624;
  assign N13534 = N16602 & N16625;
  assign N13533 = N16602 & N16626;
  assign N13532 = N16602 & N16627;
  assign N13531 = N16602 & N16628;
  assign N13530 = N16602 & N16629;
  assign N13529 = N16602 & N16630;
  assign N13528 = N16602 & N16631;
  assign N13527 = N16602 & N16632;
  assign N13526 = N16602 & N16633;
  assign N13525 = N16602 & N16634;
  assign predict_o = (N16)? N1057 : 
                     (N17)? 1'b0 : 1'b0;
  assign N16 = r_v_i;
  assign N17 = N27;
  assign { N15971, N15970, N15969, N15968, N15967, N15966, N15965, N15964, N15963, N15962, N15961, N15960, N15959, N15958, N15957, N15956, N15955, N15954, N15953, N15952, N15951, N15950, N15949, N15948, N15947, N15946, N15945, N15944, N15943, N15942, N15941, N15940, N15939, N15938, N15937, N15936, N15935, N15934, N15933, N15932, N15931, N15930, N15929, N15928, N15927, N15926, N15925, N15924, N15923, N15922, N15921, N15920, N15919, N15918, N15917, N15916, N15915, N15914, N15913, N15912, N15911, N15910, N15909, N15908, N15907, N15906, N15905, N15904, N15903, N15902, N15901, N15900, N15899, N15898, N15897, N15896, N15895, N15894, N15893, N15892, N15891, N15890, N15889, N15888, N15887, N15886, N15885, N15884, N15883, N15882, N15881, N15880, N15879, N15878, N15877, N15876, N15875, N15874, N15873, N15872, N15871, N15870, N15869, N15868, N15867, N15866, N15865, N15864, N15863, N15862, N15861, N15860, N15859, N15858, N15857, N15856, N15855, N15854, N15853, N15852, N15851, N15850, N15849, N15848, N15847, N15846, N15845, N15844, N15843, N15842, N15841, N15840, N15839, N15838, N15837, N15836, N15835, N15834, N15833, N15832, N15831, N15830, N15829, N15828, N15827, N15826, N15825, N15824, N15823, N15822, N15821, N15820, N15819, N15818, N15817, N15816, N15815, N15814, N15813, N15812, N15811, N15810, N15809, N15808, N15807, N15806, N15805, N15804, N15803, N15802, N15801, N15800, N15799, N15798, N15797, N15796, N15795, N15794, N15793, N15792, N15791, N15790, N15789, N15788, N15787, N15786, N15785, N15784, N15783, N15782, N15781, N15780, N15779, N15778, N15777, N15776, N15775, N15774, N15773, N15772, N15771, N15770, N15769, N15768, N15767, N15766, N15765, N15764, N15763, N15762, N15761, N15760, N15759, N15758, N15757, N15756, N15755, N15754, N15753, N15752, N15751, N15750, N15749, N15748, N15747, N15746, N15745, N15744, N15743, N15742, N15741, N15740, N15739, N15738, N15737, N15736, N15735, N15734, N15733, N15732, N15731, N15730, N15729, N15728, N15727, N15726, N15725, N15724, N15723, N15722, N15721, N15720, N15719, N15718, N15717, N15716, N15715, N15714, N15713, N15712, N15711, N15710, N15709, N15708, N15707, N15706, N15705, N15704, N15703, N15702, N15701, N15700, N15699, N15698, N15697, N15696, N15695, N15694, N15693, N15692, N15691, N15690, N15689, N15688, N15687, N15686, N15685, N15684, N15683, N15682, N15681, N15680, N15679, N15678, N15677, N15676, N15675, N15674, N15673, N15672, N15671, N15670, N15669, N15668, N15667, N15666, N15665, N15664, N15663, N15662, N15661, N15660, N15659, N15658, N15657, N15656, N15655, N15654, N15653, N15652, N15651, N15650, N15649, N15648, N15647, N15646, N15645, N15644, N15643, N15642, N15641, N15640, N15639, N15638, N15637, N15636, N15635, N15634, N15633, N15632, N15631, N15630, N15629, N15628, N15627, N15626, N15625, N15624, N15623, N15622, N15621, N15620, N15619, N15618, N15617, N15616, N15615, N15614, N15613, N15612, N15611, N15610, N15609, N15608, N15607, N15606, N15605, N15604, N15603, N15602, N15601, N15600, N15599, N15598, N15597, N15596, N15595, N15594, N15593, N15592, N15591, N15590, N15589, N15588, N15587, N15586, N15585, N15584, N15583, N15582, N15581, N15580, N15579, N15578, N15577, N15576, N15575, N15574, N15573, N15572, N15571, N15570, N15569, N15568, N15567, N15566, N15565, N15564, N15563, N15562, N15561, N15560, N15559, N15558, N15557, N15556, N15555, N15554, N15553, N15552, N15551, N15550, N15549, N15548, N15547, N15546, N15545, N15544, N15543, N15542, N15541, N15540, N15539, N15538, N15537, N15536, N15535, N15534, N15533, N15532, N15531, N15530, N15529, N15528, N15527, N15526, N15525, N15524, N15523, N15522, N15521, N15520, N15519, N15518, N15517, N15516, N15515, N15514, N15513, N15512, N15511, N15510, N15509, N15508, N15507, N15506, N15505, N15504, N15503, N15502, N15501, N15500, N15499, N15498, N15497, N15496, N15495, N15494, N15493, N15492, N15491, N15490, N15489, N15488, N15487, N15486, N15485, N15484, N15483, N15482, N15481, N15480, N15479, N15478, N15477, N15476, N15475, N15474, N15473, N15472, N15471, N15470, N15469, N15468, N15467, N15466, N15463, N15460, N15457, N15454, N15451, N15448 } = (N18)? { N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N20)? { N5076, N5075, N5074, N5073, N5072, N5071, N5070, N5069, N5068, N5067, N5066, N5065, N5064, N5063, N5062, N5061, N5060, N5059, N5058, N5057, N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043, N5042, N5041, N5040, N5039, N5038, N5037, N5036, N5035, N5034, N5033, N5032, N5031, N5030, N5029, N5028, N5027, N5026, N5025, N5024, N5023, N5022, N5021, N5020, N5019, N5018, N5017, N5016, N5015, N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, N4995, N4994, N4993, N4992, N4991, N4990, N4989, N4988, N4987, N4986, N4985, N4984, N4983, N4982, N4981, N4980, N4979, N4978, N4977, N4976, N4975, N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961, N4960, N4959, N4958, N4957, N4956, N4955, N4954, N4953, N4952, N4951, N4950, N4949, N4948, N4947, N4946, N4945, N4944, N4943, N4942, N4941, N4940, N4939, N4938, N4937, N4936, N4935, N4934, N4933, N4932, N4931, N4930, N4929, N4928, N4927, N4926, N4925, N4924, N4923, N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, N4903, N4902, N4901, N4900, N4899, N4898, N4897, N4896, N4895, N4894, N4893, N4892, N4891, N4890, N4889, N4888, N4887, N4886, N4885, N4884, N4883, N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869, N4868, N4867, N4866, N4865, N4864, N4863, N4862, N4861, N4860, N4859, N4858, N4857, N4856, N4855, N4854, N4853, N4852, N4851, N4850, N4849, N4848, N4847, N4846, N4845, N4844, N4843, N4842, N4841, N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, N4820, N4819, N4818, N4817, N4816, N4815, N4814, N4813, N4812, N4811, N4810, N4809, N4808, N4807, N4806, N4805, N4804, N4803, N4802, N4801, N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787, N4786, N4785, N4784, N4783, N4782, N4781, N4780, N4779, N4778, N4777, N4776, N4775, N4774, N4773, N4772, N4771, N4770, N4769, N4768, N4767, N4766, N4765, N4764, N4763, N4762, N4761, N4760, N4759, N4758, N4757, N4756, N4755, N4754, N4753, N4752, N4751, N4750, N4749, N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, N4728, N4727, N4726, N4725, N4724, N4723, N4722, N4721, N4720, N4719, N4718, N4717, N4716, N4715, N4714, N4713, N4712, N4711, N4710, N4709, N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695, N4694, N4693, N4692, N4691, N4690, N4689, N4688, N4687, N4686, N4685, N4684, N4683, N4682, N4681, N4680, N4679, N4678, N4677, N4676, N4675, N4674, N4673, N4672, N4671, N4670, N4669, N4668, N4667, N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, N4646, N4645, N4644, N4643, N4642, N4641, N4640, N4639, N4638, N4637, N4636, N4635, N4634, N4633, N4632, N4631, N4630, N4629, N4628, N4627, N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613, N4612, N4611, N4610, N4609, N4608, N4607, N4606, N4605, N4604, N4603, N4602, N4601, N4600, N4599, N4598, N4597, N4596, N4595, N4594, N4593, N4592, N4591, N4590, N4589, N4588, N4587, N4586, N4585, N4584, N4583, N4582, N4581, N4580, N4579, N4578, N4577, N4576, N4575, N4574, N4573, N4572, N4571, N4570, N4569, N4568, N4567, N4566, N4565 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N21)? { N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N22)? { N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N23)? { N10253, N10252, N10251, N10250, N10249, N10248, N10247, N10246, N10245, N10244, N10243, N10242, N10241, N10240, N10239, N10238, N10237, N10236, N10235, N10234, N10233, N10232, N10231, N10230, N10229, N10228, N10227, N10226, N10225, N10224, N10223, N10222, N10221, N10220, N10219, N10218, N10217, N10216, N10215, N10214, N10213, N10212, N10211, N10210, N10209, N10208, N10207, N10206, N10205, N10204, N10203, N10202, N10201, N10200, N10199, N10198, N10197, N10196, N10195, N10194, N10193, N10192, N10191, N10190, N10189, N10188, N10187, N10186, N10185, N10184, N10183, N10182, N10181, N10180, N10179, N10178, N10177, N10176, N10175, N10174, N10173, N10172, N10171, N10170, N10169, N10168, N10167, N10166, N10165, N10164, N10163, N10162, N10161, N10160, N10159, N10158, N10157, N10156, N10155, N10154, N10153, N10152, N10151, N10150, N10149, N10148, N10147, N10146, N10145, N10144, N10143, N10142, N10141, N10140, N10139, N10138, N10137, N10136, N10135, N10134, N10133, N10132, N10131, N10130, N10129, N10128, N10127, N10126, N10125, N10124, N10123, N10122, N10121, N10120, N10119, N10118, N10117, N10116, N10115, N10114, N10113, N10112, N10111, N10110, N10109, N10108, N10107, N10106, N10105, N10104, N10103, N10102, N10101, N10100, N10099, N10098, N10097, N10096, N10095, N10094, N10093, N10092, N10091, N10090, N10089, N10088, N10087, N10086, N10085, N10084, N10083, N10082, N10081, N10080, N10079, N10078, N10077, N10076, N10075, N10074, N10073, N10072, N10071, N10070, N10069, N10068, N10067, N10066, N10065, N10064, N10063, N10062, N10061, N10060, N10059, N10058, N10057, N10056, N10055, N10054, N10053, N10052, N10051, N10050, N10049, N10048, N10047, N10046, N10045, N10044, N10043, N10042, N10041, N10040, N10039, N10038, N10037, N10036, N10035, N10034, N10033, N10032, N10031, N10030, N10029, N10028, N10027, N10026, N10025, N10024, N10023, N10022, N10021, N10020, N10019, N10018, N10017, N10016, N10015, N10014, N10013, N10012, N10011, N10010, N10009, N10008, N10007, N10006, N10005, N10004, N10003, N10002, N10001, N10000, N9999, N9998, N9997, N9996, N9995, N9994, N9993, N9992, N9991, N9990, N9989, N9988, N9987, N9986, N9985, N9984, N9983, N9982, N9981, N9980, N9979, N9978, N9977, N9976, N9975, N9974, N9973, N9972, N9971, N9970, N9969, N9968, N9967, N9966, N9965, N9964, N9963, N9962, N9961, N9960, N9959, N9958, N9957, N9956, N9955, N9954, N9953, N9952, N9951, N9950, N9949, N9948, N9947, N9946, N9945, N9944, N9943, N9942, N9941, N9940, N9939, N9938, N9937, N9936, N9935, N9934, N9933, N9932, N9931, N9930, N9929, N9928, N9927, N9926, N9925, N9924, N9923, N9922, N9921, N9920, N9919, N9918, N9917, N9916, N9915, N9914, N9913, N9912, N9911, N9910, N9909, N9908, N9907, N9906, N9905, N9904, N9903, N9902, N9901, N9900, N9899, N9898, N9897, N9896, N9895, N9894, N9893, N9892, N9891, N9890, N9889, N9888, N9887, N9886, N9885, N9884, N9883, N9882, N9881, N9880, N9879, N9878, N9877, N9876, N9875, N9874, N9873, N9872, N9871, N9870, N9869, N9868, N9867, N9866, N9865, N9864, N9863, N9862, N9861, N9860, N9859, N9858, N9857, N9856, N9855, N9854, N9853, N9852, N9851, N9850, N9849, N9848, N9847, N9846, N9845, N9844, N9843, N9842, N9841, N9840, N9839, N9838, N9837, N9836, N9835, N9834, N9833, N9832, N9831, N9830, N9829, N9828, N9827, N9826, N9825, N9824, N9823, N9822, N9821, N9820, N9819, N9818, N9817, N9816, N9815, N9814, N9813, N9812, N9811, N9810, N9809, N9808, N9807, N9806, N9805, N9804, N9803, N9802, N9801, N9800, N9799, N9798, N9797, N9796, N9795, N9794, N9793, N9792, N9791, N9790, N9789, N9788, N9787, N9786, N9785, N9784, N9783, N9782, N9781, N9780, N9779, N9778, N9777, N9776, N9775, N9774, N9773, N9772, N9771, N9770, N9769, N9768, N9767, N9766, N9765, N9764, N9763, N9762, N9761, N9760, N9759, N9758, N9757, N9756, N9755, N9754, N9753, N9752, N9751, N9750, N9749, N9748, N9747, N9746, N9745, N9744, N9743, N9742 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N24)? { N14036, N14035, N14034, N14033, N14032, N14031, N14030, N14029, N14028, N14027, N14026, N14025, N14024, N14023, N14022, N14021, N14020, N14019, N14018, N14017, N14016, N14015, N14014, N14013, N14012, N14011, N14010, N14009, N14008, N14007, N14006, N14005, N14004, N14003, N14002, N14001, N14000, N13999, N13998, N13997, N13996, N13995, N13994, N13993, N13992, N13991, N13990, N13989, N13988, N13987, N13986, N13985, N13984, N13983, N13982, N13981, N13980, N13979, N13978, N13977, N13976, N13975, N13974, N13973, N13972, N13971, N13970, N13969, N13968, N13967, N13966, N13965, N13964, N13963, N13962, N13961, N13960, N13959, N13958, N13957, N13956, N13955, N13954, N13953, N13952, N13951, N13950, N13949, N13948, N13947, N13946, N13945, N13944, N13943, N13942, N13941, N13940, N13939, N13938, N13937, N13936, N13935, N13934, N13933, N13932, N13931, N13930, N13929, N13928, N13927, N13926, N13925, N13924, N13923, N13922, N13921, N13920, N13919, N13918, N13917, N13916, N13915, N13914, N13913, N13912, N13911, N13910, N13909, N13908, N13907, N13906, N13905, N13904, N13903, N13902, N13901, N13900, N13899, N13898, N13897, N13896, N13895, N13894, N13893, N13892, N13891, N13890, N13889, N13888, N13887, N13886, N13885, N13884, N13883, N13882, N13881, N13880, N13879, N13878, N13877, N13876, N13875, N13874, N13873, N13872, N13871, N13870, N13869, N13868, N13867, N13866, N13865, N13864, N13863, N13862, N13861, N13860, N13859, N13858, N13857, N13856, N13855, N13854, N13853, N13852, N13851, N13850, N13849, N13848, N13847, N13846, N13845, N13844, N13843, N13842, N13841, N13840, N13839, N13838, N13837, N13836, N13835, N13834, N13833, N13832, N13831, N13830, N13829, N13828, N13827, N13826, N13825, N13824, N13823, N13822, N13821, N13820, N13819, N13818, N13817, N13816, N13815, N13814, N13813, N13812, N13811, N13810, N13809, N13808, N13807, N13806, N13805, N13804, N13803, N13802, N13801, N13800, N13799, N13798, N13797, N13796, N13795, N13794, N13793, N13792, N13791, N13790, N13789, N13788, N13787, N13786, N13785, N13784, N13783, N13782, N13781, N13780, N13779, N13778, N13777, N13776, N13775, N13774, N13773, N13772, N13771, N13770, N13769, N13768, N13767, N13766, N13765, N13764, N13763, N13762, N13761, N13760, N13759, N13758, N13757, N13756, N13755, N13754, N13753, N13752, N13751, N13750, N13749, N13748, N13747, N13746, N13745, N13744, N13743, N13742, N13741, N13740, N13739, N13738, N13737, N13736, N13735, N13734, N13733, N13732, N13731, N13730, N13729, N13728, N13727, N13726, N13725, N13724, N13723, N13722, N13721, N13720, N13719, N13718, N13717, N13716, N13715, N13714, N13713, N13712, N13711, N13710, N13709, N13708, N13707, N13706, N13705, N13704, N13703, N13702, N13701, N13700, N13699, N13698, N13697, N13696, N13695, N13694, N13693, N13692, N13691, N13690, N13689, N13688, N13687, N13686, N13685, N13684, N13683, N13682, N13681, N13680, N13679, N13678, N13677, N13676, N13675, N13674, N13673, N13672, N13671, N13670, N13669, N13668, N13667, N13666, N13665, N13664, N13663, N13662, N13661, N13660, N13659, N13658, N13657, N13656, N13655, N13654, N13653, N13652, N13651, N13650, N13649, N13648, N13647, N13646, N13645, N13644, N13643, N13642, N13641, N13640, N13639, N13638, N13637, N13636, N13635, N13634, N13633, N13632, N13631, N13630, N13629, N13628, N13627, N13626, N13625, N13624, N13623, N13622, N13621, N13620, N13619, N13618, N13617, N13616, N13615, N13614, N13613, N13612, N13611, N13610, N13609, N13608, N13607, N13606, N13605, N13604, N13603, N13602, N13601, N13600, N13599, N13598, N13597, N13596, N13595, N13594, N13593, N13592, N13591, N13590, N13589, N13588, N13587, N13586, N13585, N13584, N13583, N13582, N13581, N13580, N13579, N13578, N13577, N13576, N13575, N13574, N13573, N13572, N13571, N13570, N13569, N13568, N13567, N13566, N13565, N13564, N13563, N13562, N13561, N13560, N13559, N13558, N13557, N13556, N13555, N13554, N13553, N13552, N13551, N13550, N13549, N13548, N13547, N13546, N13545, N13544, N13543, N13542, N13541, N13540, N13539, N13538, N13537, N13536, N13535, N13534, N13533, N13532, N13531, N13530, N13529, N13528, N13527, N13526, N13525 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N25)? { N14036, N14035, N14034, N14033, N14032, N14031, N14030, N14029, N14028, N14027, N14026, N14025, N14024, N14023, N14022, N14021, N14020, N14019, N14018, N14017, N14016, N14015, N14014, N14013, N14012, N14011, N14010, N14009, N14008, N14007, N14006, N14005, N14004, N14003, N14002, N14001, N14000, N13999, N13998, N13997, N13996, N13995, N13994, N13993, N13992, N13991, N13990, N13989, N13988, N13987, N13986, N13985, N13984, N13983, N13982, N13981, N13980, N13979, N13978, N13977, N13976, N13975, N13974, N13973, N13972, N13971, N13970, N13969, N13968, N13967, N13966, N13965, N13964, N13963, N13962, N13961, N13960, N13959, N13958, N13957, N13956, N13955, N13954, N13953, N13952, N13951, N13950, N13949, N13948, N13947, N13946, N13945, N13944, N13943, N13942, N13941, N13940, N13939, N13938, N13937, N13936, N13935, N13934, N13933, N13932, N13931, N13930, N13929, N13928, N13927, N13926, N13925, N13924, N13923, N13922, N13921, N13920, N13919, N13918, N13917, N13916, N13915, N13914, N13913, N13912, N13911, N13910, N13909, N13908, N13907, N13906, N13905, N13904, N13903, N13902, N13901, N13900, N13899, N13898, N13897, N13896, N13895, N13894, N13893, N13892, N13891, N13890, N13889, N13888, N13887, N13886, N13885, N13884, N13883, N13882, N13881, N13880, N13879, N13878, N13877, N13876, N13875, N13874, N13873, N13872, N13871, N13870, N13869, N13868, N13867, N13866, N13865, N13864, N13863, N13862, N13861, N13860, N13859, N13858, N13857, N13856, N13855, N13854, N13853, N13852, N13851, N13850, N13849, N13848, N13847, N13846, N13845, N13844, N13843, N13842, N13841, N13840, N13839, N13838, N13837, N13836, N13835, N13834, N13833, N13832, N13831, N13830, N13829, N13828, N13827, N13826, N13825, N13824, N13823, N13822, N13821, N13820, N13819, N13818, N13817, N13816, N13815, N13814, N13813, N13812, N13811, N13810, N13809, N13808, N13807, N13806, N13805, N13804, N13803, N13802, N13801, N13800, N13799, N13798, N13797, N13796, N13795, N13794, N13793, N13792, N13791, N13790, N13789, N13788, N13787, N13786, N13785, N13784, N13783, N13782, N13781, N13780, N13779, N13778, N13777, N13776, N13775, N13774, N13773, N13772, N13771, N13770, N13769, N13768, N13767, N13766, N13765, N13764, N13763, N13762, N13761, N13760, N13759, N13758, N13757, N13756, N13755, N13754, N13753, N13752, N13751, N13750, N13749, N13748, N13747, N13746, N13745, N13744, N13743, N13742, N13741, N13740, N13739, N13738, N13737, N13736, N13735, N13734, N13733, N13732, N13731, N13730, N13729, N13728, N13727, N13726, N13725, N13724, N13723, N13722, N13721, N13720, N13719, N13718, N13717, N13716, N13715, N13714, N13713, N13712, N13711, N13710, N13709, N13708, N13707, N13706, N13705, N13704, N13703, N13702, N13701, N13700, N13699, N13698, N13697, N13696, N13695, N13694, N13693, N13692, N13691, N13690, N13689, N13688, N13687, N13686, N13685, N13684, N13683, N13682, N13681, N13680, N13679, N13678, N13677, N13676, N13675, N13674, N13673, N13672, N13671, N13670, N13669, N13668, N13667, N13666, N13665, N13664, N13663, N13662, N13661, N13660, N13659, N13658, N13657, N13656, N13655, N13654, N13653, N13652, N13651, N13650, N13649, N13648, N13647, N13646, N13645, N13644, N13643, N13642, N13641, N13640, N13639, N13638, N13637, N13636, N13635, N13634, N13633, N13632, N13631, N13630, N13629, N13628, N13627, N13626, N13625, N13624, N13623, N13622, N13621, N13620, N13619, N13618, N13617, N13616, N13615, N13614, N13613, N13612, N13611, N13610, N13609, N13608, N13607, N13606, N13605, N13604, N13603, N13602, N13601, N13600, N13599, N13598, N13597, N13596, N13595, N13594, N13593, N13592, N13591, N13590, N13589, N13588, N13587, N13586, N13585, N13584, N13583, N13582, N13581, N13580, N13579, N13578, N13577, N13576, N13575, N13574, N13573, N13572, N13571, N13570, N13569, N13568, N13567, N13566, N13565, N13564, N13563, N13562, N13561, N13560, N13559, N13558, N13557, N13556, N13555, N13554, N13553, N13552, N13551, N13550, N13549, N13548, N13547, N13546, N13545, N13544, N13543, N13542, N13541, N13540, N13539, N13538, N13537, N13536, N13535, N13534, N13533, N13532, N13531, N13530, N13529, N13528, N13527, N13526, N13525 } : 1'b0;
  assign N18 = N2670;
  assign N19 = N2673;
  assign N20 = N2676;
  assign N21 = N2678;
  assign N22 = N2681;
  assign N23 = N2683;
  assign N24 = N2686;
  assign N25 = N2688;
  assign { N15465, N15464, N15462, N15461, N15459, N15458, N15456, N15455, N15453, N15452, N15450, N15449 } = (N18)? { N5077, 1'b1, N5077, 1'b1, N5077, 1'b1, N5077, 1'b1, N5077, 1'b1, N5077, 1'b1 } : 
                                                                                                              (N19)? { N6760, 1'b1, N6760, 1'b1, N6760, 1'b1, N6760, 1'b1, N6760, 1'b1, N6760, 1'b1 } : 
                                                                                                              (N20)? { N8267, 1'b1, N8267, 1'b1, N8267, 1'b1, N8267, 1'b1, N8267, 1'b1, N8267, 1'b1 } : 
                                                                                                              (N21)? { N10254, 1'b1, N10254, 1'b1, N10254, 1'b1, N10254, 1'b1, N10254, 1'b1, N10254, 1'b1 } : 
                                                                                                              (N22)? { N11087, N11088, N11087, N11088, N11087, N11088, N11087, N11088, N11087, N11088, N11087, N11088 } : 
                                                                                                              (N23)? { N12112, N12818, N12112, N12818, N12112, N12818, N12112, N12818, N12112, N12818, N12112, N12818 } : 
                                                                                                              (N24)? { N13523, N13524, N13523, N13524, N13523, N13524, N13523, N13524, N13523, N13524, N13523, N13524 } : 
                                                                                                              (N25)? { N14741, N15447, N14741, N15447, N14741, N15447, N14741, N15447, N14741, N15447, N14741, N15447 } : 1'b0;
  assign { N16495, N16494, N16493, N16492, N16491, N16490, N16489, N16488, N16487, N16486, N16485, N16484, N16483, N16482, N16481, N16480, N16479, N16478, N16477, N16476, N16475, N16474, N16473, N16472, N16471, N16470, N16469, N16468, N16467, N16466, N16465, N16464, N16463, N16462, N16461, N16460, N16459, N16458, N16457, N16456, N16455, N16454, N16453, N16452, N16451, N16450, N16449, N16448, N16447, N16446, N16445, N16444, N16443, N16442, N16441, N16440, N16439, N16438, N16437, N16436, N16435, N16434, N16433, N16432, N16431, N16430, N16429, N16428, N16427, N16426, N16425, N16424, N16423, N16422, N16421, N16420, N16419, N16418, N16417, N16416, N16415, N16414, N16413, N16412, N16411, N16410, N16409, N16408, N16407, N16406, N16405, N16404, N16403, N16402, N16401, N16400, N16399, N16398, N16397, N16396, N16395, N16394, N16393, N16392, N16391, N16390, N16389, N16388, N16387, N16386, N16385, N16384, N16383, N16382, N16381, N16380, N16379, N16378, N16377, N16376, N16375, N16374, N16373, N16372, N16371, N16370, N16369, N16368, N16367, N16366, N16365, N16364, N16363, N16362, N16361, N16360, N16359, N16358, N16357, N16356, N16355, N16354, N16353, N16352, N16351, N16350, N16349, N16348, N16347, N16346, N16345, N16344, N16343, N16342, N16341, N16340, N16339, N16338, N16337, N16336, N16335, N16334, N16333, N16332, N16331, N16330, N16329, N16328, N16327, N16326, N16325, N16324, N16323, N16322, N16321, N16320, N16319, N16318, N16317, N16316, N16315, N16314, N16313, N16312, N16311, N16310, N16309, N16308, N16307, N16306, N16305, N16304, N16303, N16302, N16301, N16300, N16299, N16298, N16297, N16296, N16295, N16294, N16293, N16292, N16291, N16290, N16289, N16288, N16287, N16286, N16285, N16284, N16283, N16282, N16281, N16280, N16279, N16278, N16277, N16276, N16275, N16274, N16273, N16272, N16271, N16270, N16269, N16268, N16267, N16266, N16265, N16264, N16263, N16262, N16261, N16260, N16259, N16258, N16257, N16256, N16255, N16254, N16253, N16252, N16251, N16250, N16249, N16248, N16247, N16246, N16245, N16244, N16243, N16242, N16241, N16240, N16239, N16238, N16237, N16236, N16235, N16234, N16233, N16232, N16231, N16230, N16229, N16228, N16227, N16226, N16225, N16224, N16223, N16222, N16221, N16220, N16219, N16218, N16217, N16216, N16215, N16214, N16213, N16212, N16211, N16210, N16209, N16208, N16207, N16206, N16205, N16204, N16203, N16202, N16201, N16200, N16199, N16198, N16197, N16196, N16195, N16194, N16193, N16192, N16191, N16190, N16189, N16188, N16187, N16186, N16185, N16184, N16183, N16182, N16181, N16180, N16179, N16178, N16177, N16176, N16175, N16174, N16173, N16172, N16171, N16170, N16169, N16168, N16167, N16166, N16165, N16164, N16163, N16162, N16161, N16160, N16159, N16158, N16157, N16156, N16155, N16154, N16153, N16152, N16151, N16150, N16149, N16148, N16147, N16146, N16145, N16144, N16143, N16142, N16141, N16140, N16139, N16138, N16137, N16136, N16135, N16134, N16133, N16132, N16131, N16130, N16129, N16128, N16127, N16126, N16125, N16124, N16123, N16122, N16121, N16120, N16119, N16118, N16117, N16116, N16115, N16114, N16113, N16112, N16111, N16110, N16109, N16108, N16107, N16106, N16105, N16104, N16103, N16102, N16101, N16100, N16099, N16098, N16097, N16096, N16095, N16094, N16093, N16092, N16091, N16090, N16089, N16088, N16087, N16086, N16085, N16084, N16083, N16082, N16081, N16080, N16079, N16078, N16077, N16076, N16075, N16074, N16073, N16072, N16071, N16070, N16069, N16068, N16067, N16066, N16065, N16064, N16063, N16062, N16061, N16060, N16059, N16058, N16057, N16056, N16055, N16054, N16053, N16052, N16051, N16050, N16049, N16048, N16047, N16046, N16045, N16044, N16043, N16042, N16041, N16040, N16039, N16038, N16037, N16036, N16035, N16034, N16033, N16032, N16031, N16030, N16029, N16028, N16027, N16026, N16025, N16024, N16023, N16022, N16021, N16020, N16019, N16018, N16017, N16016, N16015, N16014, N16013, N16012, N16011, N16010, N16009, N16008, N16007, N16006, N16005, N16004, N16003, N16002, N16001, N16000, N15999, N15998, N15997, N15996, N15995, N15994, N15993, N15992, N15991, N15990, N15987, N15984, N15981, N15978, N15975, N15972 } = (N26)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N16497)? { N15971, N15970, N15969, N15968, N15967, N15966, N15965, N15964, N15963, N15962, N15961, N15960, N15959, N15958, N15957, N15956, N15955, N15954, N15953, N15952, N15951, N15950, N15949, N15948, N15947, N15946, N15945, N15944, N15943, N15942, N15941, N15940, N15939, N15938, N15937, N15936, N15935, N15934, N15933, N15932, N15931, N15930, N15929, N15928, N15927, N15926, N15925, N15924, N15923, N15922, N15921, N15920, N15919, N15918, N15917, N15916, N15915, N15914, N15913, N15912, N15911, N15910, N15909, N15908, N15907, N15906, N15905, N15904, N15903, N15902, N15901, N15900, N15899, N15898, N15897, N15896, N15895, N15894, N15893, N15892, N15891, N15890, N15889, N15888, N15887, N15886, N15885, N15884, N15883, N15882, N15881, N15880, N15879, N15878, N15877, N15876, N15875, N15874, N15873, N15872, N15871, N15870, N15869, N15868, N15867, N15866, N15865, N15864, N15863, N15862, N15861, N15860, N15859, N15858, N15857, N15856, N15855, N15854, N15853, N15852, N15851, N15850, N15849, N15848, N15847, N15846, N15845, N15844, N15843, N15842, N15841, N15840, N15839, N15838, N15837, N15836, N15835, N15834, N15833, N15832, N15831, N15830, N15829, N15828, N15827, N15826, N15825, N15824, N15823, N15822, N15821, N15820, N15819, N15818, N15817, N15816, N15815, N15814, N15813, N15812, N15811, N15810, N15809, N15808, N15807, N15806, N15805, N15804, N15803, N15802, N15801, N15800, N15799, N15798, N15797, N15796, N15795, N15794, N15793, N15792, N15791, N15790, N15789, N15788, N15787, N15786, N15785, N15784, N15783, N15782, N15781, N15780, N15779, N15778, N15777, N15776, N15775, N15774, N15773, N15772, N15771, N15770, N15769, N15768, N15767, N15766, N15765, N15764, N15763, N15762, N15761, N15760, N15759, N15758, N15757, N15756, N15755, N15754, N15753, N15752, N15751, N15750, N15749, N15748, N15747, N15746, N15745, N15744, N15743, N15742, N15741, N15740, N15739, N15738, N15737, N15736, N15735, N15734, N15733, N15732, N15731, N15730, N15729, N15728, N15727, N15726, N15725, N15724, N15723, N15722, N15721, N15720, N15719, N15718, N15717, N15716, N15715, N15714, N15713, N15712, N15711, N15710, N15709, N15708, N15707, N15706, N15705, N15704, N15703, N15702, N15701, N15700, N15699, N15698, N15697, N15696, N15695, N15694, N15693, N15692, N15691, N15690, N15689, N15688, N15687, N15686, N15685, N15684, N15683, N15682, N15681, N15680, N15679, N15678, N15677, N15676, N15675, N15674, N15673, N15672, N15671, N15670, N15669, N15668, N15667, N15666, N15665, N15664, N15663, N15662, N15661, N15660, N15659, N15658, N15657, N15656, N15655, N15654, N15653, N15652, N15651, N15650, N15649, N15648, N15647, N15646, N15645, N15644, N15643, N15642, N15641, N15640, N15639, N15638, N15637, N15636, N15635, N15634, N15633, N15632, N15631, N15630, N15629, N15628, N15627, N15626, N15625, N15624, N15623, N15622, N15621, N15620, N15619, N15618, N15617, N15616, N15615, N15614, N15613, N15612, N15611, N15610, N15609, N15608, N15607, N15606, N15605, N15604, N15603, N15602, N15601, N15600, N15599, N15598, N15597, N15596, N15595, N15594, N15593, N15592, N15591, N15590, N15589, N15588, N15587, N15586, N15585, N15584, N15583, N15582, N15581, N15580, N15579, N15578, N15577, N15576, N15575, N15574, N15573, N15572, N15571, N15570, N15569, N15568, N15567, N15566, N15565, N15564, N15563, N15562, N15561, N15560, N15559, N15558, N15557, N15556, N15555, N15554, N15553, N15552, N15551, N15550, N15549, N15548, N15547, N15546, N15545, N15544, N15543, N15542, N15541, N15540, N15539, N15538, N15537, N15536, N15535, N15534, N15533, N15532, N15531, N15530, N15529, N15528, N15527, N15526, N15525, N15524, N15523, N15522, N15521, N15520, N15519, N15518, N15517, N15516, N15515, N15514, N15513, N15512, N15511, N15510, N15509, N15508, N15507, N15506, N15505, N15504, N15503, N15502, N15501, N15500, N15499, N15498, N15497, N15496, N15495, N15494, N15493, N15492, N15491, N15490, N15489, N15488, N15487, N15486, N15485, N15484, N15483, N15482, N15481, N15480, N15479, N15478, N15477, N15476, N15475, N15474, N15473, N15472, N15471, N15470, N15469, N15468, N15467, N15466, N15463, N15460, N15457, N15454, N15451, N15448 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1059)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N26 = reset_i;
  assign { N15989, N15988, N15986, N15985, N15983, N15982, N15980, N15979, N15977, N15976, N15974, N15973 } = (N26)? { 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                                                                                                              (N16497)? { N15465, N15464, N15462, N15461, N15459, N15458, N15456, N15455, N15453, N15452, N15450, N15449 } : 1'b0;
  assign N27 = ~r_v_i;
  assign N28 = ~idx_r_i[0];
  assign N29 = ~idx_r_i[1];
  assign N30 = N28 & N29;
  assign N31 = N28 & idx_r_i[1];
  assign N32 = idx_r_i[0] & N29;
  assign N33 = idx_r_i[0] & idx_r_i[1];
  assign N34 = ~idx_r_i[2];
  assign N35 = N30 & N34;
  assign N36 = N30 & idx_r_i[2];
  assign N37 = N32 & N34;
  assign N38 = N32 & idx_r_i[2];
  assign N39 = N31 & N34;
  assign N40 = N31 & idx_r_i[2];
  assign N41 = N33 & N34;
  assign N42 = N33 & idx_r_i[2];
  assign N43 = ~idx_r_i[3];
  assign N44 = N35 & N43;
  assign N45 = N35 & idx_r_i[3];
  assign N46 = N37 & N43;
  assign N47 = N37 & idx_r_i[3];
  assign N48 = N39 & N43;
  assign N49 = N39 & idx_r_i[3];
  assign N50 = N41 & N43;
  assign N51 = N41 & idx_r_i[3];
  assign N52 = N36 & N43;
  assign N53 = N36 & idx_r_i[3];
  assign N54 = N38 & N43;
  assign N55 = N38 & idx_r_i[3];
  assign N56 = N40 & N43;
  assign N57 = N40 & idx_r_i[3];
  assign N58 = N42 & N43;
  assign N59 = N42 & idx_r_i[3];
  assign N60 = ~idx_r_i[4];
  assign N61 = N44 & N60;
  assign N62 = N44 & idx_r_i[4];
  assign N63 = N46 & N60;
  assign N64 = N46 & idx_r_i[4];
  assign N65 = N48 & N60;
  assign N66 = N48 & idx_r_i[4];
  assign N67 = N50 & N60;
  assign N68 = N50 & idx_r_i[4];
  assign N69 = N52 & N60;
  assign N70 = N52 & idx_r_i[4];
  assign N71 = N54 & N60;
  assign N72 = N54 & idx_r_i[4];
  assign N73 = N56 & N60;
  assign N74 = N56 & idx_r_i[4];
  assign N75 = N58 & N60;
  assign N76 = N58 & idx_r_i[4];
  assign N77 = N45 & N60;
  assign N78 = N45 & idx_r_i[4];
  assign N79 = N47 & N60;
  assign N80 = N47 & idx_r_i[4];
  assign N81 = N49 & N60;
  assign N82 = N49 & idx_r_i[4];
  assign N83 = N51 & N60;
  assign N84 = N51 & idx_r_i[4];
  assign N85 = N53 & N60;
  assign N86 = N53 & idx_r_i[4];
  assign N87 = N55 & N60;
  assign N88 = N55 & idx_r_i[4];
  assign N89 = N57 & N60;
  assign N90 = N57 & idx_r_i[4];
  assign N91 = N59 & N60;
  assign N92 = N59 & idx_r_i[4];
  assign N93 = ~idx_r_i[5];
  assign N94 = N61 & N93;
  assign N95 = N61 & idx_r_i[5];
  assign N96 = N63 & N93;
  assign N97 = N63 & idx_r_i[5];
  assign N98 = N65 & N93;
  assign N99 = N65 & idx_r_i[5];
  assign N100 = N67 & N93;
  assign N101 = N67 & idx_r_i[5];
  assign N102 = N69 & N93;
  assign N103 = N69 & idx_r_i[5];
  assign N104 = N71 & N93;
  assign N105 = N71 & idx_r_i[5];
  assign N106 = N73 & N93;
  assign N107 = N73 & idx_r_i[5];
  assign N108 = N75 & N93;
  assign N109 = N75 & idx_r_i[5];
  assign N110 = N77 & N93;
  assign N111 = N77 & idx_r_i[5];
  assign N112 = N79 & N93;
  assign N113 = N79 & idx_r_i[5];
  assign N114 = N81 & N93;
  assign N115 = N81 & idx_r_i[5];
  assign N116 = N83 & N93;
  assign N117 = N83 & idx_r_i[5];
  assign N118 = N85 & N93;
  assign N119 = N85 & idx_r_i[5];
  assign N120 = N87 & N93;
  assign N121 = N87 & idx_r_i[5];
  assign N122 = N89 & N93;
  assign N123 = N89 & idx_r_i[5];
  assign N124 = N91 & N93;
  assign N125 = N91 & idx_r_i[5];
  assign N126 = N62 & N93;
  assign N127 = N62 & idx_r_i[5];
  assign N128 = N64 & N93;
  assign N129 = N64 & idx_r_i[5];
  assign N130 = N66 & N93;
  assign N131 = N66 & idx_r_i[5];
  assign N132 = N68 & N93;
  assign N133 = N68 & idx_r_i[5];
  assign N134 = N70 & N93;
  assign N135 = N70 & idx_r_i[5];
  assign N136 = N72 & N93;
  assign N137 = N72 & idx_r_i[5];
  assign N138 = N74 & N93;
  assign N139 = N74 & idx_r_i[5];
  assign N140 = N76 & N93;
  assign N141 = N76 & idx_r_i[5];
  assign N142 = N78 & N93;
  assign N143 = N78 & idx_r_i[5];
  assign N144 = N80 & N93;
  assign N145 = N80 & idx_r_i[5];
  assign N146 = N82 & N93;
  assign N147 = N82 & idx_r_i[5];
  assign N148 = N84 & N93;
  assign N149 = N84 & idx_r_i[5];
  assign N150 = N86 & N93;
  assign N151 = N86 & idx_r_i[5];
  assign N152 = N88 & N93;
  assign N153 = N88 & idx_r_i[5];
  assign N154 = N90 & N93;
  assign N155 = N90 & idx_r_i[5];
  assign N156 = N92 & N93;
  assign N157 = N92 & idx_r_i[5];
  assign N158 = ~idx_r_i[6];
  assign N159 = N94 & N158;
  assign N160 = N94 & idx_r_i[6];
  assign N161 = N96 & N158;
  assign N162 = N96 & idx_r_i[6];
  assign N163 = N98 & N158;
  assign N164 = N98 & idx_r_i[6];
  assign N165 = N100 & N158;
  assign N166 = N100 & idx_r_i[6];
  assign N167 = N102 & N158;
  assign N168 = N102 & idx_r_i[6];
  assign N169 = N104 & N158;
  assign N170 = N104 & idx_r_i[6];
  assign N171 = N106 & N158;
  assign N172 = N106 & idx_r_i[6];
  assign N173 = N108 & N158;
  assign N174 = N108 & idx_r_i[6];
  assign N175 = N110 & N158;
  assign N176 = N110 & idx_r_i[6];
  assign N177 = N112 & N158;
  assign N178 = N112 & idx_r_i[6];
  assign N179 = N114 & N158;
  assign N180 = N114 & idx_r_i[6];
  assign N181 = N116 & N158;
  assign N182 = N116 & idx_r_i[6];
  assign N183 = N118 & N158;
  assign N184 = N118 & idx_r_i[6];
  assign N185 = N120 & N158;
  assign N186 = N120 & idx_r_i[6];
  assign N187 = N122 & N158;
  assign N188 = N122 & idx_r_i[6];
  assign N189 = N124 & N158;
  assign N190 = N124 & idx_r_i[6];
  assign N191 = N126 & N158;
  assign N192 = N126 & idx_r_i[6];
  assign N193 = N128 & N158;
  assign N194 = N128 & idx_r_i[6];
  assign N195 = N130 & N158;
  assign N196 = N130 & idx_r_i[6];
  assign N197 = N132 & N158;
  assign N198 = N132 & idx_r_i[6];
  assign N199 = N134 & N158;
  assign N200 = N134 & idx_r_i[6];
  assign N201 = N136 & N158;
  assign N202 = N136 & idx_r_i[6];
  assign N203 = N138 & N158;
  assign N204 = N138 & idx_r_i[6];
  assign N205 = N140 & N158;
  assign N206 = N140 & idx_r_i[6];
  assign N207 = N142 & N158;
  assign N208 = N142 & idx_r_i[6];
  assign N209 = N144 & N158;
  assign N210 = N144 & idx_r_i[6];
  assign N211 = N146 & N158;
  assign N212 = N146 & idx_r_i[6];
  assign N213 = N148 & N158;
  assign N214 = N148 & idx_r_i[6];
  assign N215 = N150 & N158;
  assign N216 = N150 & idx_r_i[6];
  assign N217 = N152 & N158;
  assign N218 = N152 & idx_r_i[6];
  assign N219 = N154 & N158;
  assign N220 = N154 & idx_r_i[6];
  assign N221 = N156 & N158;
  assign N222 = N156 & idx_r_i[6];
  assign N223 = N95 & N158;
  assign N224 = N95 & idx_r_i[6];
  assign N225 = N97 & N158;
  assign N226 = N97 & idx_r_i[6];
  assign N227 = N99 & N158;
  assign N228 = N99 & idx_r_i[6];
  assign N229 = N101 & N158;
  assign N230 = N101 & idx_r_i[6];
  assign N231 = N103 & N158;
  assign N232 = N103 & idx_r_i[6];
  assign N233 = N105 & N158;
  assign N234 = N105 & idx_r_i[6];
  assign N235 = N107 & N158;
  assign N236 = N107 & idx_r_i[6];
  assign N237 = N109 & N158;
  assign N238 = N109 & idx_r_i[6];
  assign N239 = N111 & N158;
  assign N240 = N111 & idx_r_i[6];
  assign N241 = N113 & N158;
  assign N242 = N113 & idx_r_i[6];
  assign N243 = N115 & N158;
  assign N244 = N115 & idx_r_i[6];
  assign N245 = N117 & N158;
  assign N246 = N117 & idx_r_i[6];
  assign N247 = N119 & N158;
  assign N248 = N119 & idx_r_i[6];
  assign N249 = N121 & N158;
  assign N250 = N121 & idx_r_i[6];
  assign N251 = N123 & N158;
  assign N252 = N123 & idx_r_i[6];
  assign N253 = N125 & N158;
  assign N254 = N125 & idx_r_i[6];
  assign N255 = N127 & N158;
  assign N256 = N127 & idx_r_i[6];
  assign N257 = N129 & N158;
  assign N258 = N129 & idx_r_i[6];
  assign N259 = N131 & N158;
  assign N260 = N131 & idx_r_i[6];
  assign N261 = N133 & N158;
  assign N262 = N133 & idx_r_i[6];
  assign N263 = N135 & N158;
  assign N264 = N135 & idx_r_i[6];
  assign N265 = N137 & N158;
  assign N266 = N137 & idx_r_i[6];
  assign N267 = N139 & N158;
  assign N268 = N139 & idx_r_i[6];
  assign N269 = N141 & N158;
  assign N270 = N141 & idx_r_i[6];
  assign N271 = N143 & N158;
  assign N272 = N143 & idx_r_i[6];
  assign N273 = N145 & N158;
  assign N274 = N145 & idx_r_i[6];
  assign N275 = N147 & N158;
  assign N276 = N147 & idx_r_i[6];
  assign N277 = N149 & N158;
  assign N278 = N149 & idx_r_i[6];
  assign N279 = N151 & N158;
  assign N280 = N151 & idx_r_i[6];
  assign N281 = N153 & N158;
  assign N282 = N153 & idx_r_i[6];
  assign N283 = N155 & N158;
  assign N284 = N155 & idx_r_i[6];
  assign N285 = N157 & N158;
  assign N286 = N157 & idx_r_i[6];
  assign N287 = ~idx_r_i[7];
  assign N288 = N159 & N287;
  assign N289 = N159 & idx_r_i[7];
  assign N290 = N161 & N287;
  assign N291 = N161 & idx_r_i[7];
  assign N292 = N163 & N287;
  assign N293 = N163 & idx_r_i[7];
  assign N294 = N165 & N287;
  assign N295 = N165 & idx_r_i[7];
  assign N296 = N167 & N287;
  assign N297 = N167 & idx_r_i[7];
  assign N298 = N169 & N287;
  assign N299 = N169 & idx_r_i[7];
  assign N300 = N171 & N287;
  assign N301 = N171 & idx_r_i[7];
  assign N302 = N173 & N287;
  assign N303 = N173 & idx_r_i[7];
  assign N304 = N175 & N287;
  assign N305 = N175 & idx_r_i[7];
  assign N306 = N177 & N287;
  assign N307 = N177 & idx_r_i[7];
  assign N308 = N179 & N287;
  assign N309 = N179 & idx_r_i[7];
  assign N310 = N181 & N287;
  assign N311 = N181 & idx_r_i[7];
  assign N312 = N183 & N287;
  assign N313 = N183 & idx_r_i[7];
  assign N314 = N185 & N287;
  assign N315 = N185 & idx_r_i[7];
  assign N316 = N187 & N287;
  assign N317 = N187 & idx_r_i[7];
  assign N318 = N189 & N287;
  assign N319 = N189 & idx_r_i[7];
  assign N320 = N191 & N287;
  assign N321 = N191 & idx_r_i[7];
  assign N322 = N193 & N287;
  assign N323 = N193 & idx_r_i[7];
  assign N324 = N195 & N287;
  assign N325 = N195 & idx_r_i[7];
  assign N326 = N197 & N287;
  assign N327 = N197 & idx_r_i[7];
  assign N328 = N199 & N287;
  assign N329 = N199 & idx_r_i[7];
  assign N330 = N201 & N287;
  assign N331 = N201 & idx_r_i[7];
  assign N332 = N203 & N287;
  assign N333 = N203 & idx_r_i[7];
  assign N334 = N205 & N287;
  assign N335 = N205 & idx_r_i[7];
  assign N336 = N207 & N287;
  assign N337 = N207 & idx_r_i[7];
  assign N338 = N209 & N287;
  assign N339 = N209 & idx_r_i[7];
  assign N340 = N211 & N287;
  assign N341 = N211 & idx_r_i[7];
  assign N342 = N213 & N287;
  assign N343 = N213 & idx_r_i[7];
  assign N344 = N215 & N287;
  assign N345 = N215 & idx_r_i[7];
  assign N346 = N217 & N287;
  assign N347 = N217 & idx_r_i[7];
  assign N348 = N219 & N287;
  assign N349 = N219 & idx_r_i[7];
  assign N350 = N221 & N287;
  assign N351 = N221 & idx_r_i[7];
  assign N352 = N223 & N287;
  assign N353 = N223 & idx_r_i[7];
  assign N354 = N225 & N287;
  assign N355 = N225 & idx_r_i[7];
  assign N356 = N227 & N287;
  assign N357 = N227 & idx_r_i[7];
  assign N358 = N229 & N287;
  assign N359 = N229 & idx_r_i[7];
  assign N360 = N231 & N287;
  assign N361 = N231 & idx_r_i[7];
  assign N362 = N233 & N287;
  assign N363 = N233 & idx_r_i[7];
  assign N364 = N235 & N287;
  assign N365 = N235 & idx_r_i[7];
  assign N366 = N237 & N287;
  assign N367 = N237 & idx_r_i[7];
  assign N368 = N239 & N287;
  assign N369 = N239 & idx_r_i[7];
  assign N370 = N241 & N287;
  assign N371 = N241 & idx_r_i[7];
  assign N372 = N243 & N287;
  assign N373 = N243 & idx_r_i[7];
  assign N374 = N245 & N287;
  assign N375 = N245 & idx_r_i[7];
  assign N376 = N247 & N287;
  assign N377 = N247 & idx_r_i[7];
  assign N378 = N249 & N287;
  assign N379 = N249 & idx_r_i[7];
  assign N380 = N251 & N287;
  assign N381 = N251 & idx_r_i[7];
  assign N382 = N253 & N287;
  assign N383 = N253 & idx_r_i[7];
  assign N384 = N255 & N287;
  assign N385 = N255 & idx_r_i[7];
  assign N386 = N257 & N287;
  assign N387 = N257 & idx_r_i[7];
  assign N388 = N259 & N287;
  assign N389 = N259 & idx_r_i[7];
  assign N390 = N261 & N287;
  assign N391 = N261 & idx_r_i[7];
  assign N392 = N263 & N287;
  assign N393 = N263 & idx_r_i[7];
  assign N394 = N265 & N287;
  assign N395 = N265 & idx_r_i[7];
  assign N396 = N267 & N287;
  assign N397 = N267 & idx_r_i[7];
  assign N398 = N269 & N287;
  assign N399 = N269 & idx_r_i[7];
  assign N400 = N271 & N287;
  assign N401 = N271 & idx_r_i[7];
  assign N402 = N273 & N287;
  assign N403 = N273 & idx_r_i[7];
  assign N404 = N275 & N287;
  assign N405 = N275 & idx_r_i[7];
  assign N406 = N277 & N287;
  assign N407 = N277 & idx_r_i[7];
  assign N408 = N279 & N287;
  assign N409 = N279 & idx_r_i[7];
  assign N410 = N281 & N287;
  assign N411 = N281 & idx_r_i[7];
  assign N412 = N283 & N287;
  assign N413 = N283 & idx_r_i[7];
  assign N414 = N285 & N287;
  assign N415 = N285 & idx_r_i[7];
  assign N416 = N160 & N287;
  assign N417 = N160 & idx_r_i[7];
  assign N418 = N162 & N287;
  assign N419 = N162 & idx_r_i[7];
  assign N420 = N164 & N287;
  assign N421 = N164 & idx_r_i[7];
  assign N422 = N166 & N287;
  assign N423 = N166 & idx_r_i[7];
  assign N424 = N168 & N287;
  assign N425 = N168 & idx_r_i[7];
  assign N426 = N170 & N287;
  assign N427 = N170 & idx_r_i[7];
  assign N428 = N172 & N287;
  assign N429 = N172 & idx_r_i[7];
  assign N430 = N174 & N287;
  assign N431 = N174 & idx_r_i[7];
  assign N432 = N176 & N287;
  assign N433 = N176 & idx_r_i[7];
  assign N434 = N178 & N287;
  assign N435 = N178 & idx_r_i[7];
  assign N436 = N180 & N287;
  assign N437 = N180 & idx_r_i[7];
  assign N438 = N182 & N287;
  assign N439 = N182 & idx_r_i[7];
  assign N440 = N184 & N287;
  assign N441 = N184 & idx_r_i[7];
  assign N442 = N186 & N287;
  assign N443 = N186 & idx_r_i[7];
  assign N444 = N188 & N287;
  assign N445 = N188 & idx_r_i[7];
  assign N446 = N190 & N287;
  assign N447 = N190 & idx_r_i[7];
  assign N448 = N192 & N287;
  assign N449 = N192 & idx_r_i[7];
  assign N450 = N194 & N287;
  assign N451 = N194 & idx_r_i[7];
  assign N452 = N196 & N287;
  assign N453 = N196 & idx_r_i[7];
  assign N454 = N198 & N287;
  assign N455 = N198 & idx_r_i[7];
  assign N456 = N200 & N287;
  assign N457 = N200 & idx_r_i[7];
  assign N458 = N202 & N287;
  assign N459 = N202 & idx_r_i[7];
  assign N460 = N204 & N287;
  assign N461 = N204 & idx_r_i[7];
  assign N462 = N206 & N287;
  assign N463 = N206 & idx_r_i[7];
  assign N464 = N208 & N287;
  assign N465 = N208 & idx_r_i[7];
  assign N466 = N210 & N287;
  assign N467 = N210 & idx_r_i[7];
  assign N468 = N212 & N287;
  assign N469 = N212 & idx_r_i[7];
  assign N470 = N214 & N287;
  assign N471 = N214 & idx_r_i[7];
  assign N472 = N216 & N287;
  assign N473 = N216 & idx_r_i[7];
  assign N474 = N218 & N287;
  assign N475 = N218 & idx_r_i[7];
  assign N476 = N220 & N287;
  assign N477 = N220 & idx_r_i[7];
  assign N478 = N222 & N287;
  assign N479 = N222 & idx_r_i[7];
  assign N480 = N224 & N287;
  assign N481 = N224 & idx_r_i[7];
  assign N482 = N226 & N287;
  assign N483 = N226 & idx_r_i[7];
  assign N484 = N228 & N287;
  assign N485 = N228 & idx_r_i[7];
  assign N486 = N230 & N287;
  assign N487 = N230 & idx_r_i[7];
  assign N488 = N232 & N287;
  assign N489 = N232 & idx_r_i[7];
  assign N490 = N234 & N287;
  assign N491 = N234 & idx_r_i[7];
  assign N492 = N236 & N287;
  assign N493 = N236 & idx_r_i[7];
  assign N494 = N238 & N287;
  assign N495 = N238 & idx_r_i[7];
  assign N496 = N240 & N287;
  assign N497 = N240 & idx_r_i[7];
  assign N498 = N242 & N287;
  assign N499 = N242 & idx_r_i[7];
  assign N500 = N244 & N287;
  assign N501 = N244 & idx_r_i[7];
  assign N502 = N246 & N287;
  assign N503 = N246 & idx_r_i[7];
  assign N504 = N248 & N287;
  assign N505 = N248 & idx_r_i[7];
  assign N506 = N250 & N287;
  assign N507 = N250 & idx_r_i[7];
  assign N508 = N252 & N287;
  assign N509 = N252 & idx_r_i[7];
  assign N510 = N254 & N287;
  assign N511 = N254 & idx_r_i[7];
  assign N512 = N256 & N287;
  assign N513 = N256 & idx_r_i[7];
  assign N514 = N258 & N287;
  assign N515 = N258 & idx_r_i[7];
  assign N516 = N260 & N287;
  assign N517 = N260 & idx_r_i[7];
  assign N518 = N262 & N287;
  assign N519 = N262 & idx_r_i[7];
  assign N520 = N264 & N287;
  assign N521 = N264 & idx_r_i[7];
  assign N522 = N266 & N287;
  assign N523 = N266 & idx_r_i[7];
  assign N524 = N268 & N287;
  assign N525 = N268 & idx_r_i[7];
  assign N526 = N270 & N287;
  assign N527 = N270 & idx_r_i[7];
  assign N528 = N272 & N287;
  assign N529 = N272 & idx_r_i[7];
  assign N530 = N274 & N287;
  assign N531 = N274 & idx_r_i[7];
  assign N532 = N276 & N287;
  assign N533 = N276 & idx_r_i[7];
  assign N534 = N278 & N287;
  assign N535 = N278 & idx_r_i[7];
  assign N536 = N280 & N287;
  assign N537 = N280 & idx_r_i[7];
  assign N538 = N282 & N287;
  assign N539 = N282 & idx_r_i[7];
  assign N540 = N284 & N287;
  assign N541 = N284 & idx_r_i[7];
  assign N542 = N286 & N287;
  assign N543 = N286 & idx_r_i[7];
  assign N544 = ~idx_r_i[8];
  assign N545 = N288 & N544;
  assign N546 = N288 & idx_r_i[8];
  assign N547 = N290 & N544;
  assign N548 = N290 & idx_r_i[8];
  assign N549 = N292 & N544;
  assign N550 = N292 & idx_r_i[8];
  assign N551 = N294 & N544;
  assign N552 = N294 & idx_r_i[8];
  assign N553 = N296 & N544;
  assign N554 = N296 & idx_r_i[8];
  assign N555 = N298 & N544;
  assign N556 = N298 & idx_r_i[8];
  assign N557 = N300 & N544;
  assign N558 = N300 & idx_r_i[8];
  assign N559 = N302 & N544;
  assign N560 = N302 & idx_r_i[8];
  assign N561 = N304 & N544;
  assign N562 = N304 & idx_r_i[8];
  assign N563 = N306 & N544;
  assign N564 = N306 & idx_r_i[8];
  assign N565 = N308 & N544;
  assign N566 = N308 & idx_r_i[8];
  assign N567 = N310 & N544;
  assign N568 = N310 & idx_r_i[8];
  assign N569 = N312 & N544;
  assign N570 = N312 & idx_r_i[8];
  assign N571 = N314 & N544;
  assign N572 = N314 & idx_r_i[8];
  assign N573 = N316 & N544;
  assign N574 = N316 & idx_r_i[8];
  assign N575 = N318 & N544;
  assign N576 = N318 & idx_r_i[8];
  assign N577 = N320 & N544;
  assign N578 = N320 & idx_r_i[8];
  assign N579 = N322 & N544;
  assign N580 = N322 & idx_r_i[8];
  assign N581 = N324 & N544;
  assign N582 = N324 & idx_r_i[8];
  assign N583 = N326 & N544;
  assign N584 = N326 & idx_r_i[8];
  assign N585 = N328 & N544;
  assign N586 = N328 & idx_r_i[8];
  assign N587 = N330 & N544;
  assign N588 = N330 & idx_r_i[8];
  assign N589 = N332 & N544;
  assign N590 = N332 & idx_r_i[8];
  assign N591 = N334 & N544;
  assign N592 = N334 & idx_r_i[8];
  assign N593 = N336 & N544;
  assign N594 = N336 & idx_r_i[8];
  assign N595 = N338 & N544;
  assign N596 = N338 & idx_r_i[8];
  assign N597 = N340 & N544;
  assign N598 = N340 & idx_r_i[8];
  assign N599 = N342 & N544;
  assign N600 = N342 & idx_r_i[8];
  assign N601 = N344 & N544;
  assign N602 = N344 & idx_r_i[8];
  assign N603 = N346 & N544;
  assign N604 = N346 & idx_r_i[8];
  assign N605 = N348 & N544;
  assign N606 = N348 & idx_r_i[8];
  assign N607 = N350 & N544;
  assign N608 = N350 & idx_r_i[8];
  assign N609 = N352 & N544;
  assign N610 = N352 & idx_r_i[8];
  assign N611 = N354 & N544;
  assign N612 = N354 & idx_r_i[8];
  assign N613 = N356 & N544;
  assign N614 = N356 & idx_r_i[8];
  assign N615 = N358 & N544;
  assign N616 = N358 & idx_r_i[8];
  assign N617 = N360 & N544;
  assign N618 = N360 & idx_r_i[8];
  assign N619 = N362 & N544;
  assign N620 = N362 & idx_r_i[8];
  assign N621 = N364 & N544;
  assign N622 = N364 & idx_r_i[8];
  assign N623 = N366 & N544;
  assign N624 = N366 & idx_r_i[8];
  assign N625 = N368 & N544;
  assign N626 = N368 & idx_r_i[8];
  assign N627 = N370 & N544;
  assign N628 = N370 & idx_r_i[8];
  assign N629 = N372 & N544;
  assign N630 = N372 & idx_r_i[8];
  assign N631 = N374 & N544;
  assign N632 = N374 & idx_r_i[8];
  assign N633 = N376 & N544;
  assign N634 = N376 & idx_r_i[8];
  assign N635 = N378 & N544;
  assign N636 = N378 & idx_r_i[8];
  assign N637 = N380 & N544;
  assign N638 = N380 & idx_r_i[8];
  assign N639 = N382 & N544;
  assign N640 = N382 & idx_r_i[8];
  assign N641 = N384 & N544;
  assign N642 = N384 & idx_r_i[8];
  assign N643 = N386 & N544;
  assign N644 = N386 & idx_r_i[8];
  assign N645 = N388 & N544;
  assign N646 = N388 & idx_r_i[8];
  assign N647 = N390 & N544;
  assign N648 = N390 & idx_r_i[8];
  assign N649 = N392 & N544;
  assign N650 = N392 & idx_r_i[8];
  assign N651 = N394 & N544;
  assign N652 = N394 & idx_r_i[8];
  assign N653 = N396 & N544;
  assign N654 = N396 & idx_r_i[8];
  assign N655 = N398 & N544;
  assign N656 = N398 & idx_r_i[8];
  assign N657 = N400 & N544;
  assign N658 = N400 & idx_r_i[8];
  assign N659 = N402 & N544;
  assign N660 = N402 & idx_r_i[8];
  assign N661 = N404 & N544;
  assign N662 = N404 & idx_r_i[8];
  assign N663 = N406 & N544;
  assign N664 = N406 & idx_r_i[8];
  assign N665 = N408 & N544;
  assign N666 = N408 & idx_r_i[8];
  assign N667 = N410 & N544;
  assign N668 = N410 & idx_r_i[8];
  assign N669 = N412 & N544;
  assign N670 = N412 & idx_r_i[8];
  assign N671 = N414 & N544;
  assign N672 = N414 & idx_r_i[8];
  assign N673 = N416 & N544;
  assign N674 = N416 & idx_r_i[8];
  assign N675 = N418 & N544;
  assign N676 = N418 & idx_r_i[8];
  assign N677 = N420 & N544;
  assign N678 = N420 & idx_r_i[8];
  assign N679 = N422 & N544;
  assign N680 = N422 & idx_r_i[8];
  assign N681 = N424 & N544;
  assign N682 = N424 & idx_r_i[8];
  assign N683 = N426 & N544;
  assign N684 = N426 & idx_r_i[8];
  assign N685 = N428 & N544;
  assign N686 = N428 & idx_r_i[8];
  assign N687 = N430 & N544;
  assign N688 = N430 & idx_r_i[8];
  assign N689 = N432 & N544;
  assign N690 = N432 & idx_r_i[8];
  assign N691 = N434 & N544;
  assign N692 = N434 & idx_r_i[8];
  assign N693 = N436 & N544;
  assign N694 = N436 & idx_r_i[8];
  assign N695 = N438 & N544;
  assign N696 = N438 & idx_r_i[8];
  assign N697 = N440 & N544;
  assign N698 = N440 & idx_r_i[8];
  assign N699 = N442 & N544;
  assign N700 = N442 & idx_r_i[8];
  assign N701 = N444 & N544;
  assign N702 = N444 & idx_r_i[8];
  assign N703 = N446 & N544;
  assign N704 = N446 & idx_r_i[8];
  assign N705 = N448 & N544;
  assign N706 = N448 & idx_r_i[8];
  assign N707 = N450 & N544;
  assign N708 = N450 & idx_r_i[8];
  assign N709 = N452 & N544;
  assign N710 = N452 & idx_r_i[8];
  assign N711 = N454 & N544;
  assign N712 = N454 & idx_r_i[8];
  assign N713 = N456 & N544;
  assign N714 = N456 & idx_r_i[8];
  assign N715 = N458 & N544;
  assign N716 = N458 & idx_r_i[8];
  assign N717 = N460 & N544;
  assign N718 = N460 & idx_r_i[8];
  assign N719 = N462 & N544;
  assign N720 = N462 & idx_r_i[8];
  assign N721 = N464 & N544;
  assign N722 = N464 & idx_r_i[8];
  assign N723 = N466 & N544;
  assign N724 = N466 & idx_r_i[8];
  assign N725 = N468 & N544;
  assign N726 = N468 & idx_r_i[8];
  assign N727 = N470 & N544;
  assign N728 = N470 & idx_r_i[8];
  assign N729 = N472 & N544;
  assign N730 = N472 & idx_r_i[8];
  assign N731 = N474 & N544;
  assign N732 = N474 & idx_r_i[8];
  assign N733 = N476 & N544;
  assign N734 = N476 & idx_r_i[8];
  assign N735 = N478 & N544;
  assign N736 = N478 & idx_r_i[8];
  assign N737 = N480 & N544;
  assign N738 = N480 & idx_r_i[8];
  assign N739 = N482 & N544;
  assign N740 = N482 & idx_r_i[8];
  assign N741 = N484 & N544;
  assign N742 = N484 & idx_r_i[8];
  assign N743 = N486 & N544;
  assign N744 = N486 & idx_r_i[8];
  assign N745 = N488 & N544;
  assign N746 = N488 & idx_r_i[8];
  assign N747 = N490 & N544;
  assign N748 = N490 & idx_r_i[8];
  assign N749 = N492 & N544;
  assign N750 = N492 & idx_r_i[8];
  assign N751 = N494 & N544;
  assign N752 = N494 & idx_r_i[8];
  assign N753 = N496 & N544;
  assign N754 = N496 & idx_r_i[8];
  assign N755 = N498 & N544;
  assign N756 = N498 & idx_r_i[8];
  assign N757 = N500 & N544;
  assign N758 = N500 & idx_r_i[8];
  assign N759 = N502 & N544;
  assign N760 = N502 & idx_r_i[8];
  assign N761 = N504 & N544;
  assign N762 = N504 & idx_r_i[8];
  assign N763 = N506 & N544;
  assign N764 = N506 & idx_r_i[8];
  assign N765 = N508 & N544;
  assign N766 = N508 & idx_r_i[8];
  assign N767 = N510 & N544;
  assign N768 = N510 & idx_r_i[8];
  assign N769 = N512 & N544;
  assign N770 = N512 & idx_r_i[8];
  assign N771 = N514 & N544;
  assign N772 = N514 & idx_r_i[8];
  assign N773 = N516 & N544;
  assign N774 = N516 & idx_r_i[8];
  assign N775 = N518 & N544;
  assign N776 = N518 & idx_r_i[8];
  assign N777 = N520 & N544;
  assign N778 = N520 & idx_r_i[8];
  assign N779 = N522 & N544;
  assign N780 = N522 & idx_r_i[8];
  assign N781 = N524 & N544;
  assign N782 = N524 & idx_r_i[8];
  assign N783 = N526 & N544;
  assign N784 = N526 & idx_r_i[8];
  assign N785 = N528 & N544;
  assign N786 = N528 & idx_r_i[8];
  assign N787 = N530 & N544;
  assign N788 = N530 & idx_r_i[8];
  assign N789 = N532 & N544;
  assign N790 = N532 & idx_r_i[8];
  assign N791 = N534 & N544;
  assign N792 = N534 & idx_r_i[8];
  assign N793 = N536 & N544;
  assign N794 = N536 & idx_r_i[8];
  assign N795 = N538 & N544;
  assign N796 = N538 & idx_r_i[8];
  assign N797 = N540 & N544;
  assign N798 = N540 & idx_r_i[8];
  assign N799 = N542 & N544;
  assign N800 = N542 & idx_r_i[8];
  assign N801 = N289 & N544;
  assign N802 = N289 & idx_r_i[8];
  assign N803 = N291 & N544;
  assign N804 = N291 & idx_r_i[8];
  assign N805 = N293 & N544;
  assign N806 = N293 & idx_r_i[8];
  assign N807 = N295 & N544;
  assign N808 = N295 & idx_r_i[8];
  assign N809 = N297 & N544;
  assign N810 = N297 & idx_r_i[8];
  assign N811 = N299 & N544;
  assign N812 = N299 & idx_r_i[8];
  assign N813 = N301 & N544;
  assign N814 = N301 & idx_r_i[8];
  assign N815 = N303 & N544;
  assign N816 = N303 & idx_r_i[8];
  assign N817 = N305 & N544;
  assign N818 = N305 & idx_r_i[8];
  assign N819 = N307 & N544;
  assign N820 = N307 & idx_r_i[8];
  assign N821 = N309 & N544;
  assign N822 = N309 & idx_r_i[8];
  assign N823 = N311 & N544;
  assign N824 = N311 & idx_r_i[8];
  assign N825 = N313 & N544;
  assign N826 = N313 & idx_r_i[8];
  assign N827 = N315 & N544;
  assign N828 = N315 & idx_r_i[8];
  assign N829 = N317 & N544;
  assign N830 = N317 & idx_r_i[8];
  assign N831 = N319 & N544;
  assign N832 = N319 & idx_r_i[8];
  assign N833 = N321 & N544;
  assign N834 = N321 & idx_r_i[8];
  assign N835 = N323 & N544;
  assign N836 = N323 & idx_r_i[8];
  assign N837 = N325 & N544;
  assign N838 = N325 & idx_r_i[8];
  assign N839 = N327 & N544;
  assign N840 = N327 & idx_r_i[8];
  assign N841 = N329 & N544;
  assign N842 = N329 & idx_r_i[8];
  assign N843 = N331 & N544;
  assign N844 = N331 & idx_r_i[8];
  assign N845 = N333 & N544;
  assign N846 = N333 & idx_r_i[8];
  assign N847 = N335 & N544;
  assign N848 = N335 & idx_r_i[8];
  assign N849 = N337 & N544;
  assign N850 = N337 & idx_r_i[8];
  assign N851 = N339 & N544;
  assign N852 = N339 & idx_r_i[8];
  assign N853 = N341 & N544;
  assign N854 = N341 & idx_r_i[8];
  assign N855 = N343 & N544;
  assign N856 = N343 & idx_r_i[8];
  assign N857 = N345 & N544;
  assign N858 = N345 & idx_r_i[8];
  assign N859 = N347 & N544;
  assign N860 = N347 & idx_r_i[8];
  assign N861 = N349 & N544;
  assign N862 = N349 & idx_r_i[8];
  assign N863 = N351 & N544;
  assign N864 = N351 & idx_r_i[8];
  assign N865 = N353 & N544;
  assign N866 = N353 & idx_r_i[8];
  assign N867 = N355 & N544;
  assign N868 = N355 & idx_r_i[8];
  assign N869 = N357 & N544;
  assign N870 = N357 & idx_r_i[8];
  assign N871 = N359 & N544;
  assign N872 = N359 & idx_r_i[8];
  assign N873 = N361 & N544;
  assign N874 = N361 & idx_r_i[8];
  assign N875 = N363 & N544;
  assign N876 = N363 & idx_r_i[8];
  assign N877 = N365 & N544;
  assign N878 = N365 & idx_r_i[8];
  assign N879 = N367 & N544;
  assign N880 = N367 & idx_r_i[8];
  assign N881 = N369 & N544;
  assign N882 = N369 & idx_r_i[8];
  assign N883 = N371 & N544;
  assign N884 = N371 & idx_r_i[8];
  assign N885 = N373 & N544;
  assign N886 = N373 & idx_r_i[8];
  assign N887 = N375 & N544;
  assign N888 = N375 & idx_r_i[8];
  assign N889 = N377 & N544;
  assign N890 = N377 & idx_r_i[8];
  assign N891 = N379 & N544;
  assign N892 = N379 & idx_r_i[8];
  assign N893 = N381 & N544;
  assign N894 = N381 & idx_r_i[8];
  assign N895 = N383 & N544;
  assign N896 = N383 & idx_r_i[8];
  assign N897 = N385 & N544;
  assign N898 = N385 & idx_r_i[8];
  assign N899 = N387 & N544;
  assign N900 = N387 & idx_r_i[8];
  assign N901 = N389 & N544;
  assign N902 = N389 & idx_r_i[8];
  assign N903 = N391 & N544;
  assign N904 = N391 & idx_r_i[8];
  assign N905 = N393 & N544;
  assign N906 = N393 & idx_r_i[8];
  assign N907 = N395 & N544;
  assign N908 = N395 & idx_r_i[8];
  assign N909 = N397 & N544;
  assign N910 = N397 & idx_r_i[8];
  assign N911 = N399 & N544;
  assign N912 = N399 & idx_r_i[8];
  assign N913 = N401 & N544;
  assign N914 = N401 & idx_r_i[8];
  assign N915 = N403 & N544;
  assign N916 = N403 & idx_r_i[8];
  assign N917 = N405 & N544;
  assign N918 = N405 & idx_r_i[8];
  assign N919 = N407 & N544;
  assign N920 = N407 & idx_r_i[8];
  assign N921 = N409 & N544;
  assign N922 = N409 & idx_r_i[8];
  assign N923 = N411 & N544;
  assign N924 = N411 & idx_r_i[8];
  assign N925 = N413 & N544;
  assign N926 = N413 & idx_r_i[8];
  assign N927 = N415 & N544;
  assign N928 = N415 & idx_r_i[8];
  assign N929 = N417 & N544;
  assign N930 = N417 & idx_r_i[8];
  assign N931 = N419 & N544;
  assign N932 = N419 & idx_r_i[8];
  assign N933 = N421 & N544;
  assign N934 = N421 & idx_r_i[8];
  assign N935 = N423 & N544;
  assign N936 = N423 & idx_r_i[8];
  assign N937 = N425 & N544;
  assign N938 = N425 & idx_r_i[8];
  assign N939 = N427 & N544;
  assign N940 = N427 & idx_r_i[8];
  assign N941 = N429 & N544;
  assign N942 = N429 & idx_r_i[8];
  assign N943 = N431 & N544;
  assign N944 = N431 & idx_r_i[8];
  assign N945 = N433 & N544;
  assign N946 = N433 & idx_r_i[8];
  assign N947 = N435 & N544;
  assign N948 = N435 & idx_r_i[8];
  assign N949 = N437 & N544;
  assign N950 = N437 & idx_r_i[8];
  assign N951 = N439 & N544;
  assign N952 = N439 & idx_r_i[8];
  assign N953 = N441 & N544;
  assign N954 = N441 & idx_r_i[8];
  assign N955 = N443 & N544;
  assign N956 = N443 & idx_r_i[8];
  assign N957 = N445 & N544;
  assign N958 = N445 & idx_r_i[8];
  assign N959 = N447 & N544;
  assign N960 = N447 & idx_r_i[8];
  assign N961 = N449 & N544;
  assign N962 = N449 & idx_r_i[8];
  assign N963 = N451 & N544;
  assign N964 = N451 & idx_r_i[8];
  assign N965 = N453 & N544;
  assign N966 = N453 & idx_r_i[8];
  assign N967 = N455 & N544;
  assign N968 = N455 & idx_r_i[8];
  assign N969 = N457 & N544;
  assign N970 = N457 & idx_r_i[8];
  assign N971 = N459 & N544;
  assign N972 = N459 & idx_r_i[8];
  assign N973 = N461 & N544;
  assign N974 = N461 & idx_r_i[8];
  assign N975 = N463 & N544;
  assign N976 = N463 & idx_r_i[8];
  assign N977 = N465 & N544;
  assign N978 = N465 & idx_r_i[8];
  assign N979 = N467 & N544;
  assign N980 = N467 & idx_r_i[8];
  assign N981 = N469 & N544;
  assign N982 = N469 & idx_r_i[8];
  assign N983 = N471 & N544;
  assign N984 = N471 & idx_r_i[8];
  assign N985 = N473 & N544;
  assign N986 = N473 & idx_r_i[8];
  assign N987 = N475 & N544;
  assign N988 = N475 & idx_r_i[8];
  assign N989 = N477 & N544;
  assign N990 = N477 & idx_r_i[8];
  assign N991 = N479 & N544;
  assign N992 = N479 & idx_r_i[8];
  assign N993 = N481 & N544;
  assign N994 = N481 & idx_r_i[8];
  assign N995 = N483 & N544;
  assign N996 = N483 & idx_r_i[8];
  assign N997 = N485 & N544;
  assign N998 = N485 & idx_r_i[8];
  assign N999 = N487 & N544;
  assign N1000 = N487 & idx_r_i[8];
  assign N1001 = N489 & N544;
  assign N1002 = N489 & idx_r_i[8];
  assign N1003 = N491 & N544;
  assign N1004 = N491 & idx_r_i[8];
  assign N1005 = N493 & N544;
  assign N1006 = N493 & idx_r_i[8];
  assign N1007 = N495 & N544;
  assign N1008 = N495 & idx_r_i[8];
  assign N1009 = N497 & N544;
  assign N1010 = N497 & idx_r_i[8];
  assign N1011 = N499 & N544;
  assign N1012 = N499 & idx_r_i[8];
  assign N1013 = N501 & N544;
  assign N1014 = N501 & idx_r_i[8];
  assign N1015 = N503 & N544;
  assign N1016 = N503 & idx_r_i[8];
  assign N1017 = N505 & N544;
  assign N1018 = N505 & idx_r_i[8];
  assign N1019 = N507 & N544;
  assign N1020 = N507 & idx_r_i[8];
  assign N1021 = N509 & N544;
  assign N1022 = N509 & idx_r_i[8];
  assign N1023 = N511 & N544;
  assign N1024 = N511 & idx_r_i[8];
  assign N1025 = N513 & N544;
  assign N1026 = N513 & idx_r_i[8];
  assign N1027 = N515 & N544;
  assign N1028 = N515 & idx_r_i[8];
  assign N1029 = N517 & N544;
  assign N1030 = N517 & idx_r_i[8];
  assign N1031 = N519 & N544;
  assign N1032 = N519 & idx_r_i[8];
  assign N1033 = N521 & N544;
  assign N1034 = N521 & idx_r_i[8];
  assign N1035 = N523 & N544;
  assign N1036 = N523 & idx_r_i[8];
  assign N1037 = N525 & N544;
  assign N1038 = N525 & idx_r_i[8];
  assign N1039 = N527 & N544;
  assign N1040 = N527 & idx_r_i[8];
  assign N1041 = N529 & N544;
  assign N1042 = N529 & idx_r_i[8];
  assign N1043 = N531 & N544;
  assign N1044 = N531 & idx_r_i[8];
  assign N1045 = N533 & N544;
  assign N1046 = N533 & idx_r_i[8];
  assign N1047 = N535 & N544;
  assign N1048 = N535 & idx_r_i[8];
  assign N1049 = N537 & N544;
  assign N1050 = N537 & idx_r_i[8];
  assign N1051 = N539 & N544;
  assign N1052 = N539 & idx_r_i[8];
  assign N1053 = N541 & N544;
  assign N1054 = N541 & idx_r_i[8];
  assign N1055 = N543 & N544;
  assign N1056 = N543 & idx_r_i[8];
  assign N1058 = w_v_i | reset_i;
  assign N1059 = ~N1058;
  assign N1060 = ~idx_w_i[5];
  assign N1061 = N3652 & N1060;
  assign N1062 = N3653 & N1060;
  assign N1063 = N3654 & N1060;
  assign N1064 = N3655 & N1060;
  assign N1065 = N3656 & N1060;
  assign N1066 = N3657 & N1060;
  assign N1067 = N3658 & N1060;
  assign N1068 = N3659 & N1060;
  assign N1069 = N3660 & N1060;
  assign N1070 = N3661 & N1060;
  assign N1071 = N3662 & N1060;
  assign N1072 = N3663 & N1060;
  assign N1073 = N3664 & N1060;
  assign N1074 = N3665 & N1060;
  assign N1075 = N3666 & N1060;
  assign N1076 = N3667 & N1060;
  assign N1077 = N2700 & N1060;
  assign N1078 = N2702 & N1060;
  assign N1079 = N2704 & N1060;
  assign N1080 = N2706 & N1060;
  assign N1081 = N2708 & N1060;
  assign N1082 = N2710 & N1060;
  assign N1083 = N2712 & N1060;
  assign N1084 = N2714 & N1060;
  assign N1085 = N11137 & N1060;
  assign N1086 = N11139 & N1060;
  assign N1087 = N11141 & N1060;
  assign N1088 = N11143 & N1060;
  assign N1089 = N11145 & N1060;
  assign N1090 = N11147 & N1060;
  assign N1091 = N11149 & N1060;
  assign N1092 = N11151 & N1060;
  assign N1093 = ~idx_w_i[6];
  assign N1094 = N1061 & N1093;
  assign N1095 = N1061 & idx_w_i[6];
  assign N1096 = N1062 & N1093;
  assign N1097 = N1062 & idx_w_i[6];
  assign N1098 = N1063 & N1093;
  assign N1099 = N1063 & idx_w_i[6];
  assign N1100 = N1064 & N1093;
  assign N1101 = N1064 & idx_w_i[6];
  assign N1102 = N1065 & N1093;
  assign N1103 = N1065 & idx_w_i[6];
  assign N1104 = N1066 & N1093;
  assign N1105 = N1066 & idx_w_i[6];
  assign N1106 = N1067 & N1093;
  assign N1107 = N1067 & idx_w_i[6];
  assign N1108 = N1068 & N1093;
  assign N1109 = N1068 & idx_w_i[6];
  assign N1110 = N1069 & N1093;
  assign N1111 = N1069 & idx_w_i[6];
  assign N1112 = N1070 & N1093;
  assign N1113 = N1070 & idx_w_i[6];
  assign N1114 = N1071 & N1093;
  assign N1115 = N1071 & idx_w_i[6];
  assign N1116 = N1072 & N1093;
  assign N1117 = N1072 & idx_w_i[6];
  assign N1118 = N1073 & N1093;
  assign N1119 = N1073 & idx_w_i[6];
  assign N1120 = N1074 & N1093;
  assign N1121 = N1074 & idx_w_i[6];
  assign N1122 = N1075 & N1093;
  assign N1123 = N1075 & idx_w_i[6];
  assign N1124 = N1076 & N1093;
  assign N1125 = N1076 & idx_w_i[6];
  assign N1126 = N1077 & N1093;
  assign N1127 = N1077 & idx_w_i[6];
  assign N1128 = N1078 & N1093;
  assign N1129 = N1078 & idx_w_i[6];
  assign N1130 = N1079 & N1093;
  assign N1131 = N1079 & idx_w_i[6];
  assign N1132 = N1080 & N1093;
  assign N1133 = N1080 & idx_w_i[6];
  assign N1134 = N1081 & N1093;
  assign N1135 = N1081 & idx_w_i[6];
  assign N1136 = N1082 & N1093;
  assign N1137 = N1082 & idx_w_i[6];
  assign N1138 = N1083 & N1093;
  assign N1139 = N1083 & idx_w_i[6];
  assign N1140 = N1084 & N1093;
  assign N1141 = N1084 & idx_w_i[6];
  assign N1142 = N1085 & N1093;
  assign N1143 = N1085 & idx_w_i[6];
  assign N1144 = N1086 & N1093;
  assign N1145 = N1086 & idx_w_i[6];
  assign N1146 = N1087 & N1093;
  assign N1147 = N1087 & idx_w_i[6];
  assign N1148 = N1088 & N1093;
  assign N1149 = N1088 & idx_w_i[6];
  assign N1150 = N1089 & N1093;
  assign N1151 = N1089 & idx_w_i[6];
  assign N1152 = N1090 & N1093;
  assign N1153 = N1090 & idx_w_i[6];
  assign N1154 = N1091 & N1093;
  assign N1155 = N1091 & idx_w_i[6];
  assign N1156 = N1092 & N1093;
  assign N1157 = N1092 & idx_w_i[6];
  assign N1158 = N3669 & N1093;
  assign N1159 = N3671 & N1093;
  assign N1160 = N3673 & N1093;
  assign N1161 = N3675 & N1093;
  assign N1162 = N3677 & N1093;
  assign N1163 = N3679 & N1093;
  assign N1164 = N3681 & N1093;
  assign N1165 = N3683 & N1093;
  assign N1166 = N3685 & N1093;
  assign N1167 = N3687 & N1093;
  assign N1168 = N3689 & N1093;
  assign N1169 = N3691 & N1093;
  assign N1170 = N3693 & N1093;
  assign N1171 = N3695 & N1093;
  assign N1172 = N3697 & N1093;
  assign N1173 = N3699 & N1093;
  assign N1174 = N2756 & N1093;
  assign N1175 = N2758 & N1093;
  assign N1176 = N2760 & N1093;
  assign N1177 = N2762 & N1093;
  assign N1178 = N2764 & N1093;
  assign N1179 = N2766 & N1093;
  assign N1180 = N2768 & N1093;
  assign N1181 = N2770 & N1093;
  assign N1182 = N11201 & N1093;
  assign N1183 = N11203 & N1093;
  assign N1184 = N11205 & N1093;
  assign N1185 = N11207 & N1093;
  assign N1186 = N11209 & N1093;
  assign N1187 = N11211 & N1093;
  assign N1188 = N11213 & N1093;
  assign N1189 = N11215 & N1093;
  assign N1190 = ~idx_w_i[7];
  assign N1191 = N1094 & N1190;
  assign N1192 = N1094 & idx_w_i[7];
  assign N1193 = N1096 & N1190;
  assign N1194 = N1096 & idx_w_i[7];
  assign N1195 = N1098 & N1190;
  assign N1196 = N1098 & idx_w_i[7];
  assign N1197 = N1100 & N1190;
  assign N1198 = N1100 & idx_w_i[7];
  assign N1199 = N1102 & N1190;
  assign N1200 = N1102 & idx_w_i[7];
  assign N1201 = N1104 & N1190;
  assign N1202 = N1104 & idx_w_i[7];
  assign N1203 = N1106 & N1190;
  assign N1204 = N1106 & idx_w_i[7];
  assign N1205 = N1108 & N1190;
  assign N1206 = N1108 & idx_w_i[7];
  assign N1207 = N1110 & N1190;
  assign N1208 = N1110 & idx_w_i[7];
  assign N1209 = N1112 & N1190;
  assign N1210 = N1112 & idx_w_i[7];
  assign N1211 = N1114 & N1190;
  assign N1212 = N1114 & idx_w_i[7];
  assign N1213 = N1116 & N1190;
  assign N1214 = N1116 & idx_w_i[7];
  assign N1215 = N1118 & N1190;
  assign N1216 = N1118 & idx_w_i[7];
  assign N1217 = N1120 & N1190;
  assign N1218 = N1120 & idx_w_i[7];
  assign N1219 = N1122 & N1190;
  assign N1220 = N1122 & idx_w_i[7];
  assign N1221 = N1124 & N1190;
  assign N1222 = N1124 & idx_w_i[7];
  assign N1223 = N1126 & N1190;
  assign N1224 = N1126 & idx_w_i[7];
  assign N1225 = N1128 & N1190;
  assign N1226 = N1128 & idx_w_i[7];
  assign N1227 = N1130 & N1190;
  assign N1228 = N1130 & idx_w_i[7];
  assign N1229 = N1132 & N1190;
  assign N1230 = N1132 & idx_w_i[7];
  assign N1231 = N1134 & N1190;
  assign N1232 = N1134 & idx_w_i[7];
  assign N1233 = N1136 & N1190;
  assign N1234 = N1136 & idx_w_i[7];
  assign N1235 = N1138 & N1190;
  assign N1236 = N1138 & idx_w_i[7];
  assign N1237 = N1140 & N1190;
  assign N1238 = N1140 & idx_w_i[7];
  assign N1239 = N1142 & N1190;
  assign N1240 = N1142 & idx_w_i[7];
  assign N1241 = N1144 & N1190;
  assign N1242 = N1144 & idx_w_i[7];
  assign N1243 = N1146 & N1190;
  assign N1244 = N1146 & idx_w_i[7];
  assign N1245 = N1148 & N1190;
  assign N1246 = N1148 & idx_w_i[7];
  assign N1247 = N1150 & N1190;
  assign N1248 = N1150 & idx_w_i[7];
  assign N1249 = N1152 & N1190;
  assign N1250 = N1152 & idx_w_i[7];
  assign N1251 = N1154 & N1190;
  assign N1252 = N1154 & idx_w_i[7];
  assign N1253 = N1156 & N1190;
  assign N1254 = N1156 & idx_w_i[7];
  assign N1255 = N1158 & N1190;
  assign N1256 = N1158 & idx_w_i[7];
  assign N1257 = N1159 & N1190;
  assign N1258 = N1159 & idx_w_i[7];
  assign N1259 = N1160 & N1190;
  assign N1260 = N1160 & idx_w_i[7];
  assign N1261 = N1161 & N1190;
  assign N1262 = N1161 & idx_w_i[7];
  assign N1263 = N1162 & N1190;
  assign N1264 = N1162 & idx_w_i[7];
  assign N1265 = N1163 & N1190;
  assign N1266 = N1163 & idx_w_i[7];
  assign N1267 = N1164 & N1190;
  assign N1268 = N1164 & idx_w_i[7];
  assign N1269 = N1165 & N1190;
  assign N1270 = N1165 & idx_w_i[7];
  assign N1271 = N1166 & N1190;
  assign N1272 = N1166 & idx_w_i[7];
  assign N1273 = N1167 & N1190;
  assign N1274 = N1167 & idx_w_i[7];
  assign N1275 = N1168 & N1190;
  assign N1276 = N1168 & idx_w_i[7];
  assign N1277 = N1169 & N1190;
  assign N1278 = N1169 & idx_w_i[7];
  assign N1279 = N1170 & N1190;
  assign N1280 = N1170 & idx_w_i[7];
  assign N1281 = N1171 & N1190;
  assign N1282 = N1171 & idx_w_i[7];
  assign N1283 = N1172 & N1190;
  assign N1284 = N1172 & idx_w_i[7];
  assign N1285 = N1173 & N1190;
  assign N1286 = N1173 & idx_w_i[7];
  assign N1287 = N1174 & N1190;
  assign N1288 = N1174 & idx_w_i[7];
  assign N1289 = N1175 & N1190;
  assign N1290 = N1175 & idx_w_i[7];
  assign N1291 = N1176 & N1190;
  assign N1292 = N1176 & idx_w_i[7];
  assign N1293 = N1177 & N1190;
  assign N1294 = N1177 & idx_w_i[7];
  assign N1295 = N1178 & N1190;
  assign N1296 = N1178 & idx_w_i[7];
  assign N1297 = N1179 & N1190;
  assign N1298 = N1179 & idx_w_i[7];
  assign N1299 = N1180 & N1190;
  assign N1300 = N1180 & idx_w_i[7];
  assign N1301 = N1181 & N1190;
  assign N1302 = N1181 & idx_w_i[7];
  assign N1303 = N1182 & N1190;
  assign N1304 = N1182 & idx_w_i[7];
  assign N1305 = N1183 & N1190;
  assign N1306 = N1183 & idx_w_i[7];
  assign N1307 = N1184 & N1190;
  assign N1308 = N1184 & idx_w_i[7];
  assign N1309 = N1185 & N1190;
  assign N1310 = N1185 & idx_w_i[7];
  assign N1311 = N1186 & N1190;
  assign N1312 = N1186 & idx_w_i[7];
  assign N1313 = N1187 & N1190;
  assign N1314 = N1187 & idx_w_i[7];
  assign N1315 = N1188 & N1190;
  assign N1316 = N1188 & idx_w_i[7];
  assign N1317 = N1189 & N1190;
  assign N1318 = N1189 & idx_w_i[7];
  assign N1319 = N1095 & N1190;
  assign N1320 = N1095 & idx_w_i[7];
  assign N1321 = N1097 & N1190;
  assign N1322 = N1097 & idx_w_i[7];
  assign N1323 = N1099 & N1190;
  assign N1324 = N1099 & idx_w_i[7];
  assign N1325 = N1101 & N1190;
  assign N1326 = N1101 & idx_w_i[7];
  assign N1327 = N1103 & N1190;
  assign N1328 = N1103 & idx_w_i[7];
  assign N1329 = N1105 & N1190;
  assign N1330 = N1105 & idx_w_i[7];
  assign N1331 = N1107 & N1190;
  assign N1332 = N1107 & idx_w_i[7];
  assign N1333 = N1109 & N1190;
  assign N1334 = N1109 & idx_w_i[7];
  assign N1335 = N1111 & N1190;
  assign N1336 = N1111 & idx_w_i[7];
  assign N1337 = N1113 & N1190;
  assign N1338 = N1113 & idx_w_i[7];
  assign N1339 = N1115 & N1190;
  assign N1340 = N1115 & idx_w_i[7];
  assign N1341 = N1117 & N1190;
  assign N1342 = N1117 & idx_w_i[7];
  assign N1343 = N1119 & N1190;
  assign N1344 = N1119 & idx_w_i[7];
  assign N1345 = N1121 & N1190;
  assign N1346 = N1121 & idx_w_i[7];
  assign N1347 = N1123 & N1190;
  assign N1348 = N1123 & idx_w_i[7];
  assign N1349 = N1125 & N1190;
  assign N1350 = N1125 & idx_w_i[7];
  assign N1351 = N1127 & N1190;
  assign N1352 = N1127 & idx_w_i[7];
  assign N1353 = N1129 & N1190;
  assign N1354 = N1129 & idx_w_i[7];
  assign N1355 = N1131 & N1190;
  assign N1356 = N1131 & idx_w_i[7];
  assign N1357 = N1133 & N1190;
  assign N1358 = N1133 & idx_w_i[7];
  assign N1359 = N1135 & N1190;
  assign N1360 = N1135 & idx_w_i[7];
  assign N1361 = N1137 & N1190;
  assign N1362 = N1137 & idx_w_i[7];
  assign N1363 = N1139 & N1190;
  assign N1364 = N1139 & idx_w_i[7];
  assign N1365 = N1141 & N1190;
  assign N1366 = N1141 & idx_w_i[7];
  assign N1367 = N1143 & N1190;
  assign N1368 = N1143 & idx_w_i[7];
  assign N1369 = N1145 & N1190;
  assign N1370 = N1145 & idx_w_i[7];
  assign N1371 = N1147 & N1190;
  assign N1372 = N1147 & idx_w_i[7];
  assign N1373 = N1149 & N1190;
  assign N1374 = N1149 & idx_w_i[7];
  assign N1375 = N1151 & N1190;
  assign N1376 = N1151 & idx_w_i[7];
  assign N1377 = N1153 & N1190;
  assign N1378 = N1153 & idx_w_i[7];
  assign N1379 = N1155 & N1190;
  assign N1380 = N1155 & idx_w_i[7];
  assign N1381 = N1157 & N1190;
  assign N1382 = N1157 & idx_w_i[7];
  assign N1383 = N3781 & N1190;
  assign N1384 = N3783 & N1190;
  assign N1385 = N3785 & N1190;
  assign N1386 = N3787 & N1190;
  assign N1387 = N3789 & N1190;
  assign N1388 = N3791 & N1190;
  assign N1389 = N3793 & N1190;
  assign N1390 = N3795 & N1190;
  assign N1391 = N3797 & N1190;
  assign N1392 = N3799 & N1190;
  assign N1393 = N3801 & N1190;
  assign N1394 = N3803 & N1190;
  assign N1395 = N3805 & N1190;
  assign N1396 = N3807 & N1190;
  assign N1397 = N3809 & N1190;
  assign N1398 = N3811 & N1190;
  assign N1399 = N2876 & N1190;
  assign N1400 = N2878 & N1190;
  assign N1401 = N2880 & N1190;
  assign N1402 = N2882 & N1190;
  assign N1403 = N2884 & N1190;
  assign N1404 = N2886 & N1190;
  assign N1405 = N2888 & N1190;
  assign N1406 = N2890 & N1190;
  assign N1407 = N11329 & N1190;
  assign N1408 = N11331 & N1190;
  assign N1409 = N11333 & N1190;
  assign N1410 = N11335 & N1190;
  assign N1411 = N11337 & N1190;
  assign N1412 = N11339 & N1190;
  assign N1413 = N11341 & N1190;
  assign N1414 = N11343 & N1190;
  assign N1415 = ~idx_w_i[8];
  assign N1416 = N1191 & N1415;
  assign N1417 = N1191 & idx_w_i[8];
  assign N1418 = N1193 & N1415;
  assign N1419 = N1193 & idx_w_i[8];
  assign N1420 = N1195 & N1415;
  assign N1421 = N1195 & idx_w_i[8];
  assign N1422 = N1197 & N1415;
  assign N1423 = N1197 & idx_w_i[8];
  assign N1424 = N1199 & N1415;
  assign N1425 = N1199 & idx_w_i[8];
  assign N1426 = N1201 & N1415;
  assign N1427 = N1201 & idx_w_i[8];
  assign N1428 = N1203 & N1415;
  assign N1429 = N1203 & idx_w_i[8];
  assign N1430 = N1205 & N1415;
  assign N1431 = N1205 & idx_w_i[8];
  assign N1432 = N1207 & N1415;
  assign N1433 = N1207 & idx_w_i[8];
  assign N1434 = N1209 & N1415;
  assign N1435 = N1209 & idx_w_i[8];
  assign N1436 = N1211 & N1415;
  assign N1437 = N1211 & idx_w_i[8];
  assign N1438 = N1213 & N1415;
  assign N1439 = N1213 & idx_w_i[8];
  assign N1440 = N1215 & N1415;
  assign N1441 = N1215 & idx_w_i[8];
  assign N1442 = N1217 & N1415;
  assign N1443 = N1217 & idx_w_i[8];
  assign N1444 = N1219 & N1415;
  assign N1445 = N1219 & idx_w_i[8];
  assign N1446 = N1221 & N1415;
  assign N1447 = N1221 & idx_w_i[8];
  assign N1448 = N1223 & N1415;
  assign N1449 = N1223 & idx_w_i[8];
  assign N1450 = N1225 & N1415;
  assign N1451 = N1225 & idx_w_i[8];
  assign N1452 = N1227 & N1415;
  assign N1453 = N1227 & idx_w_i[8];
  assign N1454 = N1229 & N1415;
  assign N1455 = N1229 & idx_w_i[8];
  assign N1456 = N1231 & N1415;
  assign N1457 = N1231 & idx_w_i[8];
  assign N1458 = N1233 & N1415;
  assign N1459 = N1233 & idx_w_i[8];
  assign N1460 = N1235 & N1415;
  assign N1461 = N1235 & idx_w_i[8];
  assign N1462 = N1237 & N1415;
  assign N1463 = N1237 & idx_w_i[8];
  assign N1464 = N1239 & N1415;
  assign N1465 = N1239 & idx_w_i[8];
  assign N1466 = N1241 & N1415;
  assign N1467 = N1241 & idx_w_i[8];
  assign N1468 = N1243 & N1415;
  assign N1469 = N1243 & idx_w_i[8];
  assign N1470 = N1245 & N1415;
  assign N1471 = N1245 & idx_w_i[8];
  assign N1472 = N1247 & N1415;
  assign N1473 = N1247 & idx_w_i[8];
  assign N1474 = N1249 & N1415;
  assign N1475 = N1249 & idx_w_i[8];
  assign N1476 = N1251 & N1415;
  assign N1477 = N1251 & idx_w_i[8];
  assign N1478 = N1253 & N1415;
  assign N1479 = N1253 & idx_w_i[8];
  assign N1480 = N1255 & N1415;
  assign N1481 = N1255 & idx_w_i[8];
  assign N1482 = N1257 & N1415;
  assign N1483 = N1257 & idx_w_i[8];
  assign N1484 = N1259 & N1415;
  assign N1485 = N1259 & idx_w_i[8];
  assign N1486 = N1261 & N1415;
  assign N1487 = N1261 & idx_w_i[8];
  assign N1488 = N1263 & N1415;
  assign N1489 = N1263 & idx_w_i[8];
  assign N1490 = N1265 & N1415;
  assign N1491 = N1265 & idx_w_i[8];
  assign N1492 = N1267 & N1415;
  assign N1493 = N1267 & idx_w_i[8];
  assign N1494 = N1269 & N1415;
  assign N1495 = N1269 & idx_w_i[8];
  assign N1496 = N1271 & N1415;
  assign N1497 = N1271 & idx_w_i[8];
  assign N1498 = N1273 & N1415;
  assign N1499 = N1273 & idx_w_i[8];
  assign N1500 = N1275 & N1415;
  assign N1501 = N1275 & idx_w_i[8];
  assign N1502 = N1277 & N1415;
  assign N1503 = N1277 & idx_w_i[8];
  assign N1504 = N1279 & N1415;
  assign N1505 = N1279 & idx_w_i[8];
  assign N1506 = N1281 & N1415;
  assign N1507 = N1281 & idx_w_i[8];
  assign N1508 = N1283 & N1415;
  assign N1509 = N1283 & idx_w_i[8];
  assign N1510 = N1285 & N1415;
  assign N1511 = N1285 & idx_w_i[8];
  assign N1512 = N1287 & N1415;
  assign N1513 = N1287 & idx_w_i[8];
  assign N1514 = N1289 & N1415;
  assign N1515 = N1289 & idx_w_i[8];
  assign N1516 = N1291 & N1415;
  assign N1517 = N1291 & idx_w_i[8];
  assign N1518 = N1293 & N1415;
  assign N1519 = N1293 & idx_w_i[8];
  assign N1520 = N1295 & N1415;
  assign N1521 = N1295 & idx_w_i[8];
  assign N1522 = N1297 & N1415;
  assign N1523 = N1297 & idx_w_i[8];
  assign N1524 = N1299 & N1415;
  assign N1525 = N1299 & idx_w_i[8];
  assign N1526 = N1301 & N1415;
  assign N1527 = N1301 & idx_w_i[8];
  assign N1528 = N1303 & N1415;
  assign N1529 = N1303 & idx_w_i[8];
  assign N1530 = N1305 & N1415;
  assign N1531 = N1305 & idx_w_i[8];
  assign N1532 = N1307 & N1415;
  assign N1533 = N1307 & idx_w_i[8];
  assign N1534 = N1309 & N1415;
  assign N1535 = N1309 & idx_w_i[8];
  assign N1536 = N1311 & N1415;
  assign N1537 = N1311 & idx_w_i[8];
  assign N1538 = N1313 & N1415;
  assign N1539 = N1313 & idx_w_i[8];
  assign N1540 = N1315 & N1415;
  assign N1541 = N1315 & idx_w_i[8];
  assign N1542 = N1317 & N1415;
  assign N1543 = N1317 & idx_w_i[8];
  assign N1544 = N1319 & N1415;
  assign N1545 = N1319 & idx_w_i[8];
  assign N1546 = N1321 & N1415;
  assign N1547 = N1321 & idx_w_i[8];
  assign N1548 = N1323 & N1415;
  assign N1549 = N1323 & idx_w_i[8];
  assign N1550 = N1325 & N1415;
  assign N1551 = N1325 & idx_w_i[8];
  assign N1552 = N1327 & N1415;
  assign N1553 = N1327 & idx_w_i[8];
  assign N1554 = N1329 & N1415;
  assign N1555 = N1329 & idx_w_i[8];
  assign N1556 = N1331 & N1415;
  assign N1557 = N1331 & idx_w_i[8];
  assign N1558 = N1333 & N1415;
  assign N1559 = N1333 & idx_w_i[8];
  assign N1560 = N1335 & N1415;
  assign N1561 = N1335 & idx_w_i[8];
  assign N1562 = N1337 & N1415;
  assign N1563 = N1337 & idx_w_i[8];
  assign N1564 = N1339 & N1415;
  assign N1565 = N1339 & idx_w_i[8];
  assign N1566 = N1341 & N1415;
  assign N1567 = N1341 & idx_w_i[8];
  assign N1568 = N1343 & N1415;
  assign N1569 = N1343 & idx_w_i[8];
  assign N1570 = N1345 & N1415;
  assign N1571 = N1345 & idx_w_i[8];
  assign N1572 = N1347 & N1415;
  assign N1573 = N1347 & idx_w_i[8];
  assign N1574 = N1349 & N1415;
  assign N1575 = N1349 & idx_w_i[8];
  assign N1576 = N1351 & N1415;
  assign N1577 = N1351 & idx_w_i[8];
  assign N1578 = N1353 & N1415;
  assign N1579 = N1353 & idx_w_i[8];
  assign N1580 = N1355 & N1415;
  assign N1581 = N1355 & idx_w_i[8];
  assign N1582 = N1357 & N1415;
  assign N1583 = N1357 & idx_w_i[8];
  assign N1584 = N1359 & N1415;
  assign N1585 = N1359 & idx_w_i[8];
  assign N1586 = N1361 & N1415;
  assign N1587 = N1361 & idx_w_i[8];
  assign N1588 = N1363 & N1415;
  assign N1589 = N1363 & idx_w_i[8];
  assign N1590 = N1365 & N1415;
  assign N1591 = N1365 & idx_w_i[8];
  assign N1592 = N1367 & N1415;
  assign N1593 = N1367 & idx_w_i[8];
  assign N1594 = N1369 & N1415;
  assign N1595 = N1369 & idx_w_i[8];
  assign N1596 = N1371 & N1415;
  assign N1597 = N1371 & idx_w_i[8];
  assign N1598 = N1373 & N1415;
  assign N1599 = N1373 & idx_w_i[8];
  assign N1600 = N1375 & N1415;
  assign N1601 = N1375 & idx_w_i[8];
  assign N1602 = N1377 & N1415;
  assign N1603 = N1377 & idx_w_i[8];
  assign N1604 = N1379 & N1415;
  assign N1605 = N1379 & idx_w_i[8];
  assign N1606 = N1381 & N1415;
  assign N1607 = N1381 & idx_w_i[8];
  assign N1608 = N1383 & N1415;
  assign N1609 = N1383 & idx_w_i[8];
  assign N1610 = N1384 & N1415;
  assign N1611 = N1384 & idx_w_i[8];
  assign N1612 = N1385 & N1415;
  assign N1613 = N1385 & idx_w_i[8];
  assign N1614 = N1386 & N1415;
  assign N1615 = N1386 & idx_w_i[8];
  assign N1616 = N1387 & N1415;
  assign N1617 = N1387 & idx_w_i[8];
  assign N1618 = N1388 & N1415;
  assign N1619 = N1388 & idx_w_i[8];
  assign N1620 = N1389 & N1415;
  assign N1621 = N1389 & idx_w_i[8];
  assign N1622 = N1390 & N1415;
  assign N1623 = N1390 & idx_w_i[8];
  assign N1624 = N1391 & N1415;
  assign N1625 = N1391 & idx_w_i[8];
  assign N1626 = N1392 & N1415;
  assign N1627 = N1392 & idx_w_i[8];
  assign N1628 = N1393 & N1415;
  assign N1629 = N1393 & idx_w_i[8];
  assign N1630 = N1394 & N1415;
  assign N1631 = N1394 & idx_w_i[8];
  assign N1632 = N1395 & N1415;
  assign N1633 = N1395 & idx_w_i[8];
  assign N1634 = N1396 & N1415;
  assign N1635 = N1396 & idx_w_i[8];
  assign N1636 = N1397 & N1415;
  assign N1637 = N1397 & idx_w_i[8];
  assign N1638 = N1398 & N1415;
  assign N1639 = N1398 & idx_w_i[8];
  assign N1640 = N1399 & N1415;
  assign N1641 = N1399 & idx_w_i[8];
  assign N1642 = N1400 & N1415;
  assign N1643 = N1400 & idx_w_i[8];
  assign N1644 = N1401 & N1415;
  assign N1645 = N1401 & idx_w_i[8];
  assign N1646 = N1402 & N1415;
  assign N1647 = N1402 & idx_w_i[8];
  assign N1648 = N1403 & N1415;
  assign N1649 = N1403 & idx_w_i[8];
  assign N1650 = N1404 & N1415;
  assign N1651 = N1404 & idx_w_i[8];
  assign N1652 = N1405 & N1415;
  assign N1653 = N1405 & idx_w_i[8];
  assign N1654 = N1406 & N1415;
  assign N1655 = N1406 & idx_w_i[8];
  assign N1656 = N1407 & N1415;
  assign N1657 = N1407 & idx_w_i[8];
  assign N1658 = N1408 & N1415;
  assign N1659 = N1408 & idx_w_i[8];
  assign N1660 = N1409 & N1415;
  assign N1661 = N1409 & idx_w_i[8];
  assign N1662 = N1410 & N1415;
  assign N1663 = N1410 & idx_w_i[8];
  assign N1664 = N1411 & N1415;
  assign N1665 = N1411 & idx_w_i[8];
  assign N1666 = N1412 & N1415;
  assign N1667 = N1412 & idx_w_i[8];
  assign N1668 = N1413 & N1415;
  assign N1669 = N1413 & idx_w_i[8];
  assign N1670 = N1414 & N1415;
  assign N1671 = N1414 & idx_w_i[8];
  assign N1672 = N1192 & N1415;
  assign N1673 = N1192 & idx_w_i[8];
  assign N1674 = N1194 & N1415;
  assign N1675 = N1194 & idx_w_i[8];
  assign N1676 = N1196 & N1415;
  assign N1677 = N1196 & idx_w_i[8];
  assign N1678 = N1198 & N1415;
  assign N1679 = N1198 & idx_w_i[8];
  assign N1680 = N1200 & N1415;
  assign N1681 = N1200 & idx_w_i[8];
  assign N1682 = N1202 & N1415;
  assign N1683 = N1202 & idx_w_i[8];
  assign N1684 = N1204 & N1415;
  assign N1685 = N1204 & idx_w_i[8];
  assign N1686 = N1206 & N1415;
  assign N1687 = N1206 & idx_w_i[8];
  assign N1688 = N1208 & N1415;
  assign N1689 = N1208 & idx_w_i[8];
  assign N1690 = N1210 & N1415;
  assign N1691 = N1210 & idx_w_i[8];
  assign N1692 = N1212 & N1415;
  assign N1693 = N1212 & idx_w_i[8];
  assign N1694 = N1214 & N1415;
  assign N1695 = N1214 & idx_w_i[8];
  assign N1696 = N1216 & N1415;
  assign N1697 = N1216 & idx_w_i[8];
  assign N1698 = N1218 & N1415;
  assign N1699 = N1218 & idx_w_i[8];
  assign N1700 = N1220 & N1415;
  assign N1701 = N1220 & idx_w_i[8];
  assign N1702 = N1222 & N1415;
  assign N1703 = N1222 & idx_w_i[8];
  assign N1704 = N1224 & N1415;
  assign N1705 = N1224 & idx_w_i[8];
  assign N1706 = N1226 & N1415;
  assign N1707 = N1226 & idx_w_i[8];
  assign N1708 = N1228 & N1415;
  assign N1709 = N1228 & idx_w_i[8];
  assign N1710 = N1230 & N1415;
  assign N1711 = N1230 & idx_w_i[8];
  assign N1712 = N1232 & N1415;
  assign N1713 = N1232 & idx_w_i[8];
  assign N1714 = N1234 & N1415;
  assign N1715 = N1234 & idx_w_i[8];
  assign N1716 = N1236 & N1415;
  assign N1717 = N1236 & idx_w_i[8];
  assign N1718 = N1238 & N1415;
  assign N1719 = N1238 & idx_w_i[8];
  assign N1720 = N1240 & N1415;
  assign N1721 = N1240 & idx_w_i[8];
  assign N1722 = N1242 & N1415;
  assign N1723 = N1242 & idx_w_i[8];
  assign N1724 = N1244 & N1415;
  assign N1725 = N1244 & idx_w_i[8];
  assign N1726 = N1246 & N1415;
  assign N1727 = N1246 & idx_w_i[8];
  assign N1728 = N1248 & N1415;
  assign N1729 = N1248 & idx_w_i[8];
  assign N1730 = N1250 & N1415;
  assign N1731 = N1250 & idx_w_i[8];
  assign N1732 = N1252 & N1415;
  assign N1733 = N1252 & idx_w_i[8];
  assign N1734 = N1254 & N1415;
  assign N1735 = N1254 & idx_w_i[8];
  assign N1736 = N1256 & N1415;
  assign N1737 = N1256 & idx_w_i[8];
  assign N1738 = N1258 & N1415;
  assign N1739 = N1258 & idx_w_i[8];
  assign N1740 = N1260 & N1415;
  assign N1741 = N1260 & idx_w_i[8];
  assign N1742 = N1262 & N1415;
  assign N1743 = N1262 & idx_w_i[8];
  assign N1744 = N1264 & N1415;
  assign N1745 = N1264 & idx_w_i[8];
  assign N1746 = N1266 & N1415;
  assign N1747 = N1266 & idx_w_i[8];
  assign N1748 = N1268 & N1415;
  assign N1749 = N1268 & idx_w_i[8];
  assign N1750 = N1270 & N1415;
  assign N1751 = N1270 & idx_w_i[8];
  assign N1752 = N1272 & N1415;
  assign N1753 = N1272 & idx_w_i[8];
  assign N1754 = N1274 & N1415;
  assign N1755 = N1274 & idx_w_i[8];
  assign N1756 = N1276 & N1415;
  assign N1757 = N1276 & idx_w_i[8];
  assign N1758 = N1278 & N1415;
  assign N1759 = N1278 & idx_w_i[8];
  assign N1760 = N1280 & N1415;
  assign N1761 = N1280 & idx_w_i[8];
  assign N1762 = N1282 & N1415;
  assign N1763 = N1282 & idx_w_i[8];
  assign N1764 = N1284 & N1415;
  assign N1765 = N1284 & idx_w_i[8];
  assign N1766 = N1286 & N1415;
  assign N1767 = N1286 & idx_w_i[8];
  assign N1768 = N1288 & N1415;
  assign N1769 = N1288 & idx_w_i[8];
  assign N1770 = N1290 & N1415;
  assign N1771 = N1290 & idx_w_i[8];
  assign N1772 = N1292 & N1415;
  assign N1773 = N1292 & idx_w_i[8];
  assign N1774 = N1294 & N1415;
  assign N1775 = N1294 & idx_w_i[8];
  assign N1776 = N1296 & N1415;
  assign N1777 = N1296 & idx_w_i[8];
  assign N1778 = N1298 & N1415;
  assign N1779 = N1298 & idx_w_i[8];
  assign N1780 = N1300 & N1415;
  assign N1781 = N1300 & idx_w_i[8];
  assign N1782 = N1302 & N1415;
  assign N1783 = N1302 & idx_w_i[8];
  assign N1784 = N1304 & N1415;
  assign N1785 = N1304 & idx_w_i[8];
  assign N1786 = N1306 & N1415;
  assign N1787 = N1306 & idx_w_i[8];
  assign N1788 = N1308 & N1415;
  assign N1789 = N1308 & idx_w_i[8];
  assign N1790 = N1310 & N1415;
  assign N1791 = N1310 & idx_w_i[8];
  assign N1792 = N1312 & N1415;
  assign N1793 = N1312 & idx_w_i[8];
  assign N1794 = N1314 & N1415;
  assign N1795 = N1314 & idx_w_i[8];
  assign N1796 = N1316 & N1415;
  assign N1797 = N1316 & idx_w_i[8];
  assign N1798 = N1318 & N1415;
  assign N1799 = N1318 & idx_w_i[8];
  assign N1800 = N1320 & N1415;
  assign N1801 = N1320 & idx_w_i[8];
  assign N1802 = N1322 & N1415;
  assign N1803 = N1322 & idx_w_i[8];
  assign N1804 = N1324 & N1415;
  assign N1805 = N1324 & idx_w_i[8];
  assign N1806 = N1326 & N1415;
  assign N1807 = N1326 & idx_w_i[8];
  assign N1808 = N1328 & N1415;
  assign N1809 = N1328 & idx_w_i[8];
  assign N1810 = N1330 & N1415;
  assign N1811 = N1330 & idx_w_i[8];
  assign N1812 = N1332 & N1415;
  assign N1813 = N1332 & idx_w_i[8];
  assign N1814 = N1334 & N1415;
  assign N1815 = N1334 & idx_w_i[8];
  assign N1816 = N1336 & N1415;
  assign N1817 = N1336 & idx_w_i[8];
  assign N1818 = N1338 & N1415;
  assign N1819 = N1338 & idx_w_i[8];
  assign N1820 = N1340 & N1415;
  assign N1821 = N1340 & idx_w_i[8];
  assign N1822 = N1342 & N1415;
  assign N1823 = N1342 & idx_w_i[8];
  assign N1824 = N1344 & N1415;
  assign N1825 = N1344 & idx_w_i[8];
  assign N1826 = N1346 & N1415;
  assign N1827 = N1346 & idx_w_i[8];
  assign N1828 = N1348 & N1415;
  assign N1829 = N1348 & idx_w_i[8];
  assign N1830 = N1350 & N1415;
  assign N1831 = N1350 & idx_w_i[8];
  assign N1832 = N1352 & N1415;
  assign N1833 = N1352 & idx_w_i[8];
  assign N1834 = N1354 & N1415;
  assign N1835 = N1354 & idx_w_i[8];
  assign N1836 = N1356 & N1415;
  assign N1837 = N1356 & idx_w_i[8];
  assign N1838 = N1358 & N1415;
  assign N1839 = N1358 & idx_w_i[8];
  assign N1840 = N1360 & N1415;
  assign N1841 = N1360 & idx_w_i[8];
  assign N1842 = N1362 & N1415;
  assign N1843 = N1362 & idx_w_i[8];
  assign N1844 = N1364 & N1415;
  assign N1845 = N1364 & idx_w_i[8];
  assign N1846 = N1366 & N1415;
  assign N1847 = N1366 & idx_w_i[8];
  assign N1848 = N1368 & N1415;
  assign N1849 = N1368 & idx_w_i[8];
  assign N1850 = N1370 & N1415;
  assign N1851 = N1370 & idx_w_i[8];
  assign N1852 = N1372 & N1415;
  assign N1853 = N1372 & idx_w_i[8];
  assign N1854 = N1374 & N1415;
  assign N1855 = N1374 & idx_w_i[8];
  assign N1856 = N1376 & N1415;
  assign N1857 = N1376 & idx_w_i[8];
  assign N1858 = N1378 & N1415;
  assign N1859 = N1378 & idx_w_i[8];
  assign N1860 = N1380 & N1415;
  assign N1861 = N1380 & idx_w_i[8];
  assign N1862 = N1382 & N1415;
  assign N1863 = N1382 & idx_w_i[8];
  assign N1864 = N4021 & N1415;
  assign N1865 = N4023 & N1415;
  assign N1866 = N4025 & N1415;
  assign N1867 = N4027 & N1415;
  assign N1868 = N4029 & N1415;
  assign N1869 = N4031 & N1415;
  assign N1870 = N4033 & N1415;
  assign N1871 = N4035 & N1415;
  assign N1872 = N4037 & N1415;
  assign N1873 = N4039 & N1415;
  assign N1874 = N4041 & N1415;
  assign N1875 = N4043 & N1415;
  assign N1876 = N4045 & N1415;
  assign N1877 = N4047 & N1415;
  assign N1878 = N4049 & N1415;
  assign N1879 = N4051 & N1415;
  assign N1880 = N3124 & N1415;
  assign N1881 = N3126 & N1415;
  assign N1882 = N3128 & N1415;
  assign N1883 = N3130 & N1415;
  assign N1884 = N3132 & N1415;
  assign N1885 = N3134 & N1415;
  assign N1886 = N3136 & N1415;
  assign N1887 = N3138 & N1415;
  assign N1888 = N11585 & N1415;
  assign N1889 = N11587 & N1415;
  assign N1890 = N11589 & N1415;
  assign N1891 = N11591 & N1415;
  assign N1892 = N11593 & N1415;
  assign N1893 = N11595 & N1415;
  assign N1894 = N11597 & N1415;
  assign N1895 = N11599 & N1415;
  assign N1897 = N3652 & N1060;
  assign N1898 = N3653 & N1060;
  assign N1899 = N3654 & N1060;
  assign N1900 = N3655 & N1060;
  assign N1901 = N3656 & N1060;
  assign N1902 = N3657 & N1060;
  assign N1903 = N3658 & N1060;
  assign N1904 = N3659 & N1060;
  assign N1905 = N2700 & N1060;
  assign N1906 = N2702 & N1060;
  assign N1907 = N2704 & N1060;
  assign N1908 = N2706 & N1060;
  assign N1909 = N2708 & N1060;
  assign N1910 = N2710 & N1060;
  assign N1911 = N2712 & N1060;
  assign N1912 = N2714 & N1060;
  assign N1913 = N1897 & N1093;
  assign N1914 = N1897 & idx_w_i[6];
  assign N1915 = N1898 & N1093;
  assign N1916 = N1898 & idx_w_i[6];
  assign N1917 = N1899 & N1093;
  assign N1918 = N1899 & idx_w_i[6];
  assign N1919 = N1900 & N1093;
  assign N1920 = N1900 & idx_w_i[6];
  assign N1921 = N1901 & N1093;
  assign N1922 = N1901 & idx_w_i[6];
  assign N1923 = N1902 & N1093;
  assign N1924 = N1902 & idx_w_i[6];
  assign N1925 = N1903 & N1093;
  assign N1926 = N1903 & idx_w_i[6];
  assign N1927 = N1904 & N1093;
  assign N1928 = N1904 & idx_w_i[6];
  assign N1929 = N5102 & N1093;
  assign N1930 = N5103 & N1093;
  assign N1931 = N5104 & N1093;
  assign N1932 = N5105 & N1093;
  assign N1933 = N5106 & N1093;
  assign N1934 = N5107 & N1093;
  assign N1935 = N5108 & N1093;
  assign N1936 = N5109 & N1093;
  assign N1937 = N1905 & N1093;
  assign N1938 = N1905 & idx_w_i[6];
  assign N1939 = N1906 & N1093;
  assign N1940 = N1906 & idx_w_i[6];
  assign N1941 = N1907 & N1093;
  assign N1942 = N1907 & idx_w_i[6];
  assign N1943 = N1908 & N1093;
  assign N1944 = N1908 & idx_w_i[6];
  assign N1945 = N1909 & N1093;
  assign N1946 = N1909 & idx_w_i[6];
  assign N1947 = N1910 & N1093;
  assign N1948 = N1910 & idx_w_i[6];
  assign N1949 = N1911 & N1093;
  assign N1950 = N1911 & idx_w_i[6];
  assign N1951 = N1912 & N1093;
  assign N1952 = N1912 & idx_w_i[6];
  assign N1953 = N5118 & N1093;
  assign N1954 = N5119 & N1093;
  assign N1955 = N5120 & N1093;
  assign N1956 = N5121 & N1093;
  assign N1957 = N5122 & N1093;
  assign N1958 = N5123 & N1093;
  assign N1959 = N5124 & N1093;
  assign N1960 = N5125 & N1093;
  assign N1961 = N3669 & N1093;
  assign N1962 = N3671 & N1093;
  assign N1963 = N3673 & N1093;
  assign N1964 = N3675 & N1093;
  assign N1965 = N3677 & N1093;
  assign N1966 = N3679 & N1093;
  assign N1967 = N3681 & N1093;
  assign N1968 = N3683 & N1093;
  assign N1969 = N3685 & N1093;
  assign N1970 = N3687 & N1093;
  assign N1971 = N3689 & N1093;
  assign N1972 = N3691 & N1093;
  assign N1973 = N3693 & N1093;
  assign N1974 = N3695 & N1093;
  assign N1975 = N3697 & N1093;
  assign N1976 = N3699 & N1093;
  assign N1977 = N2756 & N1093;
  assign N1978 = N2758 & N1093;
  assign N1979 = N2760 & N1093;
  assign N1980 = N2762 & N1093;
  assign N1981 = N2764 & N1093;
  assign N1982 = N2766 & N1093;
  assign N1983 = N2768 & N1093;
  assign N1984 = N2770 & N1093;
  assign N1985 = N11201 & N1093;
  assign N1986 = N11203 & N1093;
  assign N1987 = N11205 & N1093;
  assign N1988 = N11207 & N1093;
  assign N1989 = N11209 & N1093;
  assign N1990 = N11211 & N1093;
  assign N1991 = N11213 & N1093;
  assign N1992 = N11215 & N1093;
  assign N1993 = N1913 & N1190;
  assign N1994 = N1913 & idx_w_i[7];
  assign N1995 = N1915 & N1190;
  assign N1996 = N1915 & idx_w_i[7];
  assign N1997 = N1917 & N1190;
  assign N1998 = N1917 & idx_w_i[7];
  assign N1999 = N1919 & N1190;
  assign N2000 = N1919 & idx_w_i[7];
  assign N2001 = N1921 & N1190;
  assign N2002 = N1921 & idx_w_i[7];
  assign N2003 = N1923 & N1190;
  assign N2004 = N1923 & idx_w_i[7];
  assign N2005 = N1925 & N1190;
  assign N2006 = N1925 & idx_w_i[7];
  assign N2007 = N1927 & N1190;
  assign N2008 = N1927 & idx_w_i[7];
  assign N2009 = N1929 & N1190;
  assign N2010 = N1929 & idx_w_i[7];
  assign N2011 = N1930 & N1190;
  assign N2012 = N1930 & idx_w_i[7];
  assign N2013 = N1931 & N1190;
  assign N2014 = N1931 & idx_w_i[7];
  assign N2015 = N1932 & N1190;
  assign N2016 = N1932 & idx_w_i[7];
  assign N2017 = N1933 & N1190;
  assign N2018 = N1933 & idx_w_i[7];
  assign N2019 = N1934 & N1190;
  assign N2020 = N1934 & idx_w_i[7];
  assign N2021 = N1935 & N1190;
  assign N2022 = N1935 & idx_w_i[7];
  assign N2023 = N1936 & N1190;
  assign N2024 = N1936 & idx_w_i[7];
  assign N2025 = N1937 & N1190;
  assign N2026 = N1937 & idx_w_i[7];
  assign N2027 = N1939 & N1190;
  assign N2028 = N1939 & idx_w_i[7];
  assign N2029 = N1941 & N1190;
  assign N2030 = N1941 & idx_w_i[7];
  assign N2031 = N1943 & N1190;
  assign N2032 = N1943 & idx_w_i[7];
  assign N2033 = N1945 & N1190;
  assign N2034 = N1945 & idx_w_i[7];
  assign N2035 = N1947 & N1190;
  assign N2036 = N1947 & idx_w_i[7];
  assign N2037 = N1949 & N1190;
  assign N2038 = N1949 & idx_w_i[7];
  assign N2039 = N1951 & N1190;
  assign N2040 = N1951 & idx_w_i[7];
  assign N2041 = N1953 & N1190;
  assign N2042 = N1953 & idx_w_i[7];
  assign N2043 = N1954 & N1190;
  assign N2044 = N1954 & idx_w_i[7];
  assign N2045 = N1955 & N1190;
  assign N2046 = N1955 & idx_w_i[7];
  assign N2047 = N1956 & N1190;
  assign N2048 = N1956 & idx_w_i[7];
  assign N2049 = N1957 & N1190;
  assign N2050 = N1957 & idx_w_i[7];
  assign N2051 = N1958 & N1190;
  assign N2052 = N1958 & idx_w_i[7];
  assign N2053 = N1959 & N1190;
  assign N2054 = N1959 & idx_w_i[7];
  assign N2055 = N1960 & N1190;
  assign N2056 = N1960 & idx_w_i[7];
  assign N2057 = N1961 & N1190;
  assign N2058 = N1961 & idx_w_i[7];
  assign N2059 = N1962 & N1190;
  assign N2060 = N1962 & idx_w_i[7];
  assign N2061 = N1963 & N1190;
  assign N2062 = N1963 & idx_w_i[7];
  assign N2063 = N1964 & N1190;
  assign N2064 = N1964 & idx_w_i[7];
  assign N2065 = N1965 & N1190;
  assign N2066 = N1965 & idx_w_i[7];
  assign N2067 = N1966 & N1190;
  assign N2068 = N1966 & idx_w_i[7];
  assign N2069 = N1967 & N1190;
  assign N2070 = N1967 & idx_w_i[7];
  assign N2071 = N1968 & N1190;
  assign N2072 = N1968 & idx_w_i[7];
  assign N2073 = N1969 & N1190;
  assign N2074 = N1969 & idx_w_i[7];
  assign N2075 = N1970 & N1190;
  assign N2076 = N1970 & idx_w_i[7];
  assign N2077 = N1971 & N1190;
  assign N2078 = N1971 & idx_w_i[7];
  assign N2079 = N1972 & N1190;
  assign N2080 = N1972 & idx_w_i[7];
  assign N2081 = N1973 & N1190;
  assign N2082 = N1973 & idx_w_i[7];
  assign N2083 = N1974 & N1190;
  assign N2084 = N1974 & idx_w_i[7];
  assign N2085 = N1975 & N1190;
  assign N2086 = N1975 & idx_w_i[7];
  assign N2087 = N1976 & N1190;
  assign N2088 = N1976 & idx_w_i[7];
  assign N2089 = N1977 & N1190;
  assign N2090 = N1977 & idx_w_i[7];
  assign N2091 = N1978 & N1190;
  assign N2092 = N1978 & idx_w_i[7];
  assign N2093 = N1979 & N1190;
  assign N2094 = N1979 & idx_w_i[7];
  assign N2095 = N1980 & N1190;
  assign N2096 = N1980 & idx_w_i[7];
  assign N2097 = N1981 & N1190;
  assign N2098 = N1981 & idx_w_i[7];
  assign N2099 = N1982 & N1190;
  assign N2100 = N1982 & idx_w_i[7];
  assign N2101 = N1983 & N1190;
  assign N2102 = N1983 & idx_w_i[7];
  assign N2103 = N1984 & N1190;
  assign N2104 = N1984 & idx_w_i[7];
  assign N2105 = N1985 & N1190;
  assign N2106 = N1985 & idx_w_i[7];
  assign N2107 = N1986 & N1190;
  assign N2108 = N1986 & idx_w_i[7];
  assign N2109 = N1987 & N1190;
  assign N2110 = N1987 & idx_w_i[7];
  assign N2111 = N1988 & N1190;
  assign N2112 = N1988 & idx_w_i[7];
  assign N2113 = N1989 & N1190;
  assign N2114 = N1989 & idx_w_i[7];
  assign N2115 = N1990 & N1190;
  assign N2116 = N1990 & idx_w_i[7];
  assign N2117 = N1991 & N1190;
  assign N2118 = N1991 & idx_w_i[7];
  assign N2119 = N1992 & N1190;
  assign N2120 = N1992 & idx_w_i[7];
  assign N2121 = N1914 & N1190;
  assign N2122 = N1914 & idx_w_i[7];
  assign N2123 = N1916 & N1190;
  assign N2124 = N1916 & idx_w_i[7];
  assign N2125 = N1918 & N1190;
  assign N2126 = N1918 & idx_w_i[7];
  assign N2127 = N1920 & N1190;
  assign N2128 = N1920 & idx_w_i[7];
  assign N2129 = N1922 & N1190;
  assign N2130 = N1922 & idx_w_i[7];
  assign N2131 = N1924 & N1190;
  assign N2132 = N1924 & idx_w_i[7];
  assign N2133 = N1926 & N1190;
  assign N2134 = N1926 & idx_w_i[7];
  assign N2135 = N1928 & N1190;
  assign N2136 = N1928 & idx_w_i[7];
  assign N2137 = N5143 & N1190;
  assign N2138 = N5145 & N1190;
  assign N2139 = N5147 & N1190;
  assign N2140 = N5149 & N1190;
  assign N2141 = N5151 & N1190;
  assign N2142 = N5153 & N1190;
  assign N2143 = N5155 & N1190;
  assign N2144 = N5157 & N1190;
  assign N2145 = N1938 & N1190;
  assign N2146 = N1938 & idx_w_i[7];
  assign N2147 = N1940 & N1190;
  assign N2148 = N1940 & idx_w_i[7];
  assign N2149 = N1942 & N1190;
  assign N2150 = N1942 & idx_w_i[7];
  assign N2151 = N1944 & N1190;
  assign N2152 = N1944 & idx_w_i[7];
  assign N2153 = N1946 & N1190;
  assign N2154 = N1946 & idx_w_i[7];
  assign N2155 = N1948 & N1190;
  assign N2156 = N1948 & idx_w_i[7];
  assign N2157 = N1950 & N1190;
  assign N2158 = N1950 & idx_w_i[7];
  assign N2159 = N1952 & N1190;
  assign N2160 = N1952 & idx_w_i[7];
  assign N2161 = N5175 & N1190;
  assign N2162 = N5177 & N1190;
  assign N2163 = N5179 & N1190;
  assign N2164 = N5181 & N1190;
  assign N2165 = N5183 & N1190;
  assign N2166 = N5185 & N1190;
  assign N2167 = N5187 & N1190;
  assign N2168 = N5189 & N1190;
  assign N2169 = N3781 & N1190;
  assign N2170 = N3783 & N1190;
  assign N2171 = N3785 & N1190;
  assign N2172 = N3787 & N1190;
  assign N2173 = N3789 & N1190;
  assign N2174 = N3791 & N1190;
  assign N2175 = N3793 & N1190;
  assign N2176 = N3795 & N1190;
  assign N2177 = N3797 & N1190;
  assign N2178 = N3799 & N1190;
  assign N2179 = N3801 & N1190;
  assign N2180 = N3803 & N1190;
  assign N2181 = N3805 & N1190;
  assign N2182 = N3807 & N1190;
  assign N2183 = N3809 & N1190;
  assign N2184 = N3811 & N1190;
  assign N2185 = N2876 & N1190;
  assign N2186 = N2878 & N1190;
  assign N2187 = N2880 & N1190;
  assign N2188 = N2882 & N1190;
  assign N2189 = N2884 & N1190;
  assign N2190 = N2886 & N1190;
  assign N2191 = N2888 & N1190;
  assign N2192 = N2890 & N1190;
  assign N2193 = N11329 & N1190;
  assign N2194 = N11331 & N1190;
  assign N2195 = N11333 & N1190;
  assign N2196 = N11335 & N1190;
  assign N2197 = N11337 & N1190;
  assign N2198 = N11339 & N1190;
  assign N2199 = N11341 & N1190;
  assign N2200 = N11343 & N1190;
  assign N2201 = N1993 & N1415;
  assign N2202 = N1993 & idx_w_i[8];
  assign N2203 = N1995 & N1415;
  assign N2204 = N1995 & idx_w_i[8];
  assign N2205 = N1997 & N1415;
  assign N2206 = N1997 & idx_w_i[8];
  assign N2207 = N1999 & N1415;
  assign N2208 = N1999 & idx_w_i[8];
  assign N2209 = N2001 & N1415;
  assign N2210 = N2001 & idx_w_i[8];
  assign N2211 = N2003 & N1415;
  assign N2212 = N2003 & idx_w_i[8];
  assign N2213 = N2005 & N1415;
  assign N2214 = N2005 & idx_w_i[8];
  assign N2215 = N2007 & N1415;
  assign N2216 = N2007 & idx_w_i[8];
  assign N2217 = N2009 & N1415;
  assign N2218 = N2009 & idx_w_i[8];
  assign N2219 = N2011 & N1415;
  assign N2220 = N2011 & idx_w_i[8];
  assign N2221 = N2013 & N1415;
  assign N2222 = N2013 & idx_w_i[8];
  assign N2223 = N2015 & N1415;
  assign N2224 = N2015 & idx_w_i[8];
  assign N2225 = N2017 & N1415;
  assign N2226 = N2017 & idx_w_i[8];
  assign N2227 = N2019 & N1415;
  assign N2228 = N2019 & idx_w_i[8];
  assign N2229 = N2021 & N1415;
  assign N2230 = N2021 & idx_w_i[8];
  assign N2231 = N2023 & N1415;
  assign N2232 = N2023 & idx_w_i[8];
  assign N2233 = N2025 & N1415;
  assign N2234 = N2025 & idx_w_i[8];
  assign N2235 = N2027 & N1415;
  assign N2236 = N2027 & idx_w_i[8];
  assign N2237 = N2029 & N1415;
  assign N2238 = N2029 & idx_w_i[8];
  assign N2239 = N2031 & N1415;
  assign N2240 = N2031 & idx_w_i[8];
  assign N2241 = N2033 & N1415;
  assign N2242 = N2033 & idx_w_i[8];
  assign N2243 = N2035 & N1415;
  assign N2244 = N2035 & idx_w_i[8];
  assign N2245 = N2037 & N1415;
  assign N2246 = N2037 & idx_w_i[8];
  assign N2247 = N2039 & N1415;
  assign N2248 = N2039 & idx_w_i[8];
  assign N2249 = N2041 & N1415;
  assign N2250 = N2041 & idx_w_i[8];
  assign N2251 = N2043 & N1415;
  assign N2252 = N2043 & idx_w_i[8];
  assign N2253 = N2045 & N1415;
  assign N2254 = N2045 & idx_w_i[8];
  assign N2255 = N2047 & N1415;
  assign N2256 = N2047 & idx_w_i[8];
  assign N2257 = N2049 & N1415;
  assign N2258 = N2049 & idx_w_i[8];
  assign N2259 = N2051 & N1415;
  assign N2260 = N2051 & idx_w_i[8];
  assign N2261 = N2053 & N1415;
  assign N2262 = N2053 & idx_w_i[8];
  assign N2263 = N2055 & N1415;
  assign N2264 = N2055 & idx_w_i[8];
  assign N2265 = N2057 & N1415;
  assign N2266 = N2057 & idx_w_i[8];
  assign N2267 = N2059 & N1415;
  assign N2268 = N2059 & idx_w_i[8];
  assign N2269 = N2061 & N1415;
  assign N2270 = N2061 & idx_w_i[8];
  assign N2271 = N2063 & N1415;
  assign N2272 = N2063 & idx_w_i[8];
  assign N2273 = N2065 & N1415;
  assign N2274 = N2065 & idx_w_i[8];
  assign N2275 = N2067 & N1415;
  assign N2276 = N2067 & idx_w_i[8];
  assign N2277 = N2069 & N1415;
  assign N2278 = N2069 & idx_w_i[8];
  assign N2279 = N2071 & N1415;
  assign N2280 = N2071 & idx_w_i[8];
  assign N2281 = N2073 & N1415;
  assign N2282 = N2073 & idx_w_i[8];
  assign N2283 = N2075 & N1415;
  assign N2284 = N2075 & idx_w_i[8];
  assign N2285 = N2077 & N1415;
  assign N2286 = N2077 & idx_w_i[8];
  assign N2287 = N2079 & N1415;
  assign N2288 = N2079 & idx_w_i[8];
  assign N2289 = N2081 & N1415;
  assign N2290 = N2081 & idx_w_i[8];
  assign N2291 = N2083 & N1415;
  assign N2292 = N2083 & idx_w_i[8];
  assign N2293 = N2085 & N1415;
  assign N2294 = N2085 & idx_w_i[8];
  assign N2295 = N2087 & N1415;
  assign N2296 = N2087 & idx_w_i[8];
  assign N2297 = N2089 & N1415;
  assign N2298 = N2089 & idx_w_i[8];
  assign N2299 = N2091 & N1415;
  assign N2300 = N2091 & idx_w_i[8];
  assign N2301 = N2093 & N1415;
  assign N2302 = N2093 & idx_w_i[8];
  assign N2303 = N2095 & N1415;
  assign N2304 = N2095 & idx_w_i[8];
  assign N2305 = N2097 & N1415;
  assign N2306 = N2097 & idx_w_i[8];
  assign N2307 = N2099 & N1415;
  assign N2308 = N2099 & idx_w_i[8];
  assign N2309 = N2101 & N1415;
  assign N2310 = N2101 & idx_w_i[8];
  assign N2311 = N2103 & N1415;
  assign N2312 = N2103 & idx_w_i[8];
  assign N2313 = N2105 & N1415;
  assign N2314 = N2105 & idx_w_i[8];
  assign N2315 = N2107 & N1415;
  assign N2316 = N2107 & idx_w_i[8];
  assign N2317 = N2109 & N1415;
  assign N2318 = N2109 & idx_w_i[8];
  assign N2319 = N2111 & N1415;
  assign N2320 = N2111 & idx_w_i[8];
  assign N2321 = N2113 & N1415;
  assign N2322 = N2113 & idx_w_i[8];
  assign N2323 = N2115 & N1415;
  assign N2324 = N2115 & idx_w_i[8];
  assign N2325 = N2117 & N1415;
  assign N2326 = N2117 & idx_w_i[8];
  assign N2327 = N2119 & N1415;
  assign N2328 = N2119 & idx_w_i[8];
  assign N2329 = N2121 & N1415;
  assign N2330 = N2121 & idx_w_i[8];
  assign N2331 = N2123 & N1415;
  assign N2332 = N2123 & idx_w_i[8];
  assign N2333 = N2125 & N1415;
  assign N2334 = N2125 & idx_w_i[8];
  assign N2335 = N2127 & N1415;
  assign N2336 = N2127 & idx_w_i[8];
  assign N2337 = N2129 & N1415;
  assign N2338 = N2129 & idx_w_i[8];
  assign N2339 = N2131 & N1415;
  assign N2340 = N2131 & idx_w_i[8];
  assign N2341 = N2133 & N1415;
  assign N2342 = N2133 & idx_w_i[8];
  assign N2343 = N2135 & N1415;
  assign N2344 = N2135 & idx_w_i[8];
  assign N2345 = N2137 & N1415;
  assign N2346 = N2137 & idx_w_i[8];
  assign N2347 = N2138 & N1415;
  assign N2348 = N2138 & idx_w_i[8];
  assign N2349 = N2139 & N1415;
  assign N2350 = N2139 & idx_w_i[8];
  assign N2351 = N2140 & N1415;
  assign N2352 = N2140 & idx_w_i[8];
  assign N2353 = N2141 & N1415;
  assign N2354 = N2141 & idx_w_i[8];
  assign N2355 = N2142 & N1415;
  assign N2356 = N2142 & idx_w_i[8];
  assign N2357 = N2143 & N1415;
  assign N2358 = N2143 & idx_w_i[8];
  assign N2359 = N2144 & N1415;
  assign N2360 = N2144 & idx_w_i[8];
  assign N2361 = N2145 & N1415;
  assign N2362 = N2145 & idx_w_i[8];
  assign N2363 = N2147 & N1415;
  assign N2364 = N2147 & idx_w_i[8];
  assign N2365 = N2149 & N1415;
  assign N2366 = N2149 & idx_w_i[8];
  assign N2367 = N2151 & N1415;
  assign N2368 = N2151 & idx_w_i[8];
  assign N2369 = N2153 & N1415;
  assign N2370 = N2153 & idx_w_i[8];
  assign N2371 = N2155 & N1415;
  assign N2372 = N2155 & idx_w_i[8];
  assign N2373 = N2157 & N1415;
  assign N2374 = N2157 & idx_w_i[8];
  assign N2375 = N2159 & N1415;
  assign N2376 = N2159 & idx_w_i[8];
  assign N2377 = N2161 & N1415;
  assign N2378 = N2161 & idx_w_i[8];
  assign N2379 = N2162 & N1415;
  assign N2380 = N2162 & idx_w_i[8];
  assign N2381 = N2163 & N1415;
  assign N2382 = N2163 & idx_w_i[8];
  assign N2383 = N2164 & N1415;
  assign N2384 = N2164 & idx_w_i[8];
  assign N2385 = N2165 & N1415;
  assign N2386 = N2165 & idx_w_i[8];
  assign N2387 = N2166 & N1415;
  assign N2388 = N2166 & idx_w_i[8];
  assign N2389 = N2167 & N1415;
  assign N2390 = N2167 & idx_w_i[8];
  assign N2391 = N2168 & N1415;
  assign N2392 = N2168 & idx_w_i[8];
  assign N2393 = N2169 & N1415;
  assign N2394 = N2169 & idx_w_i[8];
  assign N2395 = N2170 & N1415;
  assign N2396 = N2170 & idx_w_i[8];
  assign N2397 = N2171 & N1415;
  assign N2398 = N2171 & idx_w_i[8];
  assign N2399 = N2172 & N1415;
  assign N2400 = N2172 & idx_w_i[8];
  assign N2401 = N2173 & N1415;
  assign N2402 = N2173 & idx_w_i[8];
  assign N2403 = N2174 & N1415;
  assign N2404 = N2174 & idx_w_i[8];
  assign N2405 = N2175 & N1415;
  assign N2406 = N2175 & idx_w_i[8];
  assign N2407 = N2176 & N1415;
  assign N2408 = N2176 & idx_w_i[8];
  assign N2409 = N2177 & N1415;
  assign N2410 = N2177 & idx_w_i[8];
  assign N2411 = N2178 & N1415;
  assign N2412 = N2178 & idx_w_i[8];
  assign N2413 = N2179 & N1415;
  assign N2414 = N2179 & idx_w_i[8];
  assign N2415 = N2180 & N1415;
  assign N2416 = N2180 & idx_w_i[8];
  assign N2417 = N2181 & N1415;
  assign N2418 = N2181 & idx_w_i[8];
  assign N2419 = N2182 & N1415;
  assign N2420 = N2182 & idx_w_i[8];
  assign N2421 = N2183 & N1415;
  assign N2422 = N2183 & idx_w_i[8];
  assign N2423 = N2184 & N1415;
  assign N2424 = N2184 & idx_w_i[8];
  assign N2425 = N2185 & N1415;
  assign N2426 = N2185 & idx_w_i[8];
  assign N2427 = N2186 & N1415;
  assign N2428 = N2186 & idx_w_i[8];
  assign N2429 = N2187 & N1415;
  assign N2430 = N2187 & idx_w_i[8];
  assign N2431 = N2188 & N1415;
  assign N2432 = N2188 & idx_w_i[8];
  assign N2433 = N2189 & N1415;
  assign N2434 = N2189 & idx_w_i[8];
  assign N2435 = N2190 & N1415;
  assign N2436 = N2190 & idx_w_i[8];
  assign N2437 = N2191 & N1415;
  assign N2438 = N2191 & idx_w_i[8];
  assign N2439 = N2192 & N1415;
  assign N2440 = N2192 & idx_w_i[8];
  assign N2441 = N2193 & N1415;
  assign N2442 = N2193 & idx_w_i[8];
  assign N2443 = N2194 & N1415;
  assign N2444 = N2194 & idx_w_i[8];
  assign N2445 = N2195 & N1415;
  assign N2446 = N2195 & idx_w_i[8];
  assign N2447 = N2196 & N1415;
  assign N2448 = N2196 & idx_w_i[8];
  assign N2449 = N2197 & N1415;
  assign N2450 = N2197 & idx_w_i[8];
  assign N2451 = N2198 & N1415;
  assign N2452 = N2198 & idx_w_i[8];
  assign N2453 = N2199 & N1415;
  assign N2454 = N2199 & idx_w_i[8];
  assign N2455 = N2200 & N1415;
  assign N2456 = N2200 & idx_w_i[8];
  assign N2457 = N1994 & N1415;
  assign N2458 = N1994 & idx_w_i[8];
  assign N2459 = N1996 & N1415;
  assign N2460 = N1996 & idx_w_i[8];
  assign N2461 = N1998 & N1415;
  assign N2462 = N1998 & idx_w_i[8];
  assign N2463 = N2000 & N1415;
  assign N2464 = N2000 & idx_w_i[8];
  assign N2465 = N2002 & N1415;
  assign N2466 = N2002 & idx_w_i[8];
  assign N2467 = N2004 & N1415;
  assign N2468 = N2004 & idx_w_i[8];
  assign N2469 = N2006 & N1415;
  assign N2470 = N2006 & idx_w_i[8];
  assign N2471 = N2008 & N1415;
  assign N2472 = N2008 & idx_w_i[8];
  assign N2473 = N2010 & N1415;
  assign N2474 = N2010 & idx_w_i[8];
  assign N2475 = N2012 & N1415;
  assign N2476 = N2012 & idx_w_i[8];
  assign N2477 = N2014 & N1415;
  assign N2478 = N2014 & idx_w_i[8];
  assign N2479 = N2016 & N1415;
  assign N2480 = N2016 & idx_w_i[8];
  assign N2481 = N2018 & N1415;
  assign N2482 = N2018 & idx_w_i[8];
  assign N2483 = N2020 & N1415;
  assign N2484 = N2020 & idx_w_i[8];
  assign N2485 = N2022 & N1415;
  assign N2486 = N2022 & idx_w_i[8];
  assign N2487 = N2024 & N1415;
  assign N2488 = N2024 & idx_w_i[8];
  assign N2489 = N2026 & N1415;
  assign N2490 = N2026 & idx_w_i[8];
  assign N2491 = N2028 & N1415;
  assign N2492 = N2028 & idx_w_i[8];
  assign N2493 = N2030 & N1415;
  assign N2494 = N2030 & idx_w_i[8];
  assign N2495 = N2032 & N1415;
  assign N2496 = N2032 & idx_w_i[8];
  assign N2497 = N2034 & N1415;
  assign N2498 = N2034 & idx_w_i[8];
  assign N2499 = N2036 & N1415;
  assign N2500 = N2036 & idx_w_i[8];
  assign N2501 = N2038 & N1415;
  assign N2502 = N2038 & idx_w_i[8];
  assign N2503 = N2040 & N1415;
  assign N2504 = N2040 & idx_w_i[8];
  assign N2505 = N2042 & N1415;
  assign N2506 = N2042 & idx_w_i[8];
  assign N2507 = N2044 & N1415;
  assign N2508 = N2044 & idx_w_i[8];
  assign N2509 = N2046 & N1415;
  assign N2510 = N2046 & idx_w_i[8];
  assign N2511 = N2048 & N1415;
  assign N2512 = N2048 & idx_w_i[8];
  assign N2513 = N2050 & N1415;
  assign N2514 = N2050 & idx_w_i[8];
  assign N2515 = N2052 & N1415;
  assign N2516 = N2052 & idx_w_i[8];
  assign N2517 = N2054 & N1415;
  assign N2518 = N2054 & idx_w_i[8];
  assign N2519 = N2056 & N1415;
  assign N2520 = N2056 & idx_w_i[8];
  assign N2521 = N2058 & N1415;
  assign N2522 = N2058 & idx_w_i[8];
  assign N2523 = N2060 & N1415;
  assign N2524 = N2060 & idx_w_i[8];
  assign N2525 = N2062 & N1415;
  assign N2526 = N2062 & idx_w_i[8];
  assign N2527 = N2064 & N1415;
  assign N2528 = N2064 & idx_w_i[8];
  assign N2529 = N2066 & N1415;
  assign N2530 = N2066 & idx_w_i[8];
  assign N2531 = N2068 & N1415;
  assign N2532 = N2068 & idx_w_i[8];
  assign N2533 = N2070 & N1415;
  assign N2534 = N2070 & idx_w_i[8];
  assign N2535 = N2072 & N1415;
  assign N2536 = N2072 & idx_w_i[8];
  assign N2537 = N2074 & N1415;
  assign N2538 = N2074 & idx_w_i[8];
  assign N2539 = N2076 & N1415;
  assign N2540 = N2076 & idx_w_i[8];
  assign N2541 = N2078 & N1415;
  assign N2542 = N2078 & idx_w_i[8];
  assign N2543 = N2080 & N1415;
  assign N2544 = N2080 & idx_w_i[8];
  assign N2545 = N2082 & N1415;
  assign N2546 = N2082 & idx_w_i[8];
  assign N2547 = N2084 & N1415;
  assign N2548 = N2084 & idx_w_i[8];
  assign N2549 = N2086 & N1415;
  assign N2550 = N2086 & idx_w_i[8];
  assign N2551 = N2088 & N1415;
  assign N2552 = N2088 & idx_w_i[8];
  assign N2553 = N2090 & N1415;
  assign N2554 = N2090 & idx_w_i[8];
  assign N2555 = N2092 & N1415;
  assign N2556 = N2092 & idx_w_i[8];
  assign N2557 = N2094 & N1415;
  assign N2558 = N2094 & idx_w_i[8];
  assign N2559 = N2096 & N1415;
  assign N2560 = N2096 & idx_w_i[8];
  assign N2561 = N2098 & N1415;
  assign N2562 = N2098 & idx_w_i[8];
  assign N2563 = N2100 & N1415;
  assign N2564 = N2100 & idx_w_i[8];
  assign N2565 = N2102 & N1415;
  assign N2566 = N2102 & idx_w_i[8];
  assign N2567 = N2104 & N1415;
  assign N2568 = N2104 & idx_w_i[8];
  assign N2569 = N2106 & N1415;
  assign N2570 = N2106 & idx_w_i[8];
  assign N2571 = N2108 & N1415;
  assign N2572 = N2108 & idx_w_i[8];
  assign N2573 = N2110 & N1415;
  assign N2574 = N2110 & idx_w_i[8];
  assign N2575 = N2112 & N1415;
  assign N2576 = N2112 & idx_w_i[8];
  assign N2577 = N2114 & N1415;
  assign N2578 = N2114 & idx_w_i[8];
  assign N2579 = N2116 & N1415;
  assign N2580 = N2116 & idx_w_i[8];
  assign N2581 = N2118 & N1415;
  assign N2582 = N2118 & idx_w_i[8];
  assign N2583 = N2120 & N1415;
  assign N2584 = N2120 & idx_w_i[8];
  assign N2585 = N2122 & N1415;
  assign N2586 = N2122 & idx_w_i[8];
  assign N2587 = N2124 & N1415;
  assign N2588 = N2124 & idx_w_i[8];
  assign N2589 = N2126 & N1415;
  assign N2590 = N2126 & idx_w_i[8];
  assign N2591 = N2128 & N1415;
  assign N2592 = N2128 & idx_w_i[8];
  assign N2593 = N2130 & N1415;
  assign N2594 = N2130 & idx_w_i[8];
  assign N2595 = N2132 & N1415;
  assign N2596 = N2132 & idx_w_i[8];
  assign N2597 = N2134 & N1415;
  assign N2598 = N2134 & idx_w_i[8];
  assign N2599 = N2136 & N1415;
  assign N2600 = N2136 & idx_w_i[8];
  assign N2601 = N5375 & N1415;
  assign N2602 = N5377 & N1415;
  assign N2603 = N5379 & N1415;
  assign N2604 = N5381 & N1415;
  assign N2605 = N5383 & N1415;
  assign N2606 = N5385 & N1415;
  assign N2607 = N5387 & N1415;
  assign N2608 = N5389 & N1415;
  assign N2609 = N2146 & N1415;
  assign N2610 = N2146 & idx_w_i[8];
  assign N2611 = N2148 & N1415;
  assign N2612 = N2148 & idx_w_i[8];
  assign N2613 = N2150 & N1415;
  assign N2614 = N2150 & idx_w_i[8];
  assign N2615 = N2152 & N1415;
  assign N2616 = N2152 & idx_w_i[8];
  assign N2617 = N2154 & N1415;
  assign N2618 = N2154 & idx_w_i[8];
  assign N2619 = N2156 & N1415;
  assign N2620 = N2156 & idx_w_i[8];
  assign N2621 = N2158 & N1415;
  assign N2622 = N2158 & idx_w_i[8];
  assign N2623 = N2160 & N1415;
  assign N2624 = N2160 & idx_w_i[8];
  assign N2625 = N5407 & N1415;
  assign N2626 = N5409 & N1415;
  assign N2627 = N5411 & N1415;
  assign N2628 = N5413 & N1415;
  assign N2629 = N5415 & N1415;
  assign N2630 = N5417 & N1415;
  assign N2631 = N5419 & N1415;
  assign N2632 = N5421 & N1415;
  assign N2633 = N4021 & N1415;
  assign N2634 = N4023 & N1415;
  assign N2635 = N4025 & N1415;
  assign N2636 = N4027 & N1415;
  assign N2637 = N4029 & N1415;
  assign N2638 = N4031 & N1415;
  assign N2639 = N4033 & N1415;
  assign N2640 = N4035 & N1415;
  assign N2641 = N4037 & N1415;
  assign N2642 = N4039 & N1415;
  assign N2643 = N4041 & N1415;
  assign N2644 = N4043 & N1415;
  assign N2645 = N4045 & N1415;
  assign N2646 = N4047 & N1415;
  assign N2647 = N4049 & N1415;
  assign N2648 = N4051 & N1415;
  assign N2649 = N3124 & N1415;
  assign N2650 = N3126 & N1415;
  assign N2651 = N3128 & N1415;
  assign N2652 = N3130 & N1415;
  assign N2653 = N3132 & N1415;
  assign N2654 = N3134 & N1415;
  assign N2655 = N3136 & N1415;
  assign N2656 = N3138 & N1415;
  assign N2657 = N11585 & N1415;
  assign N2658 = N11587 & N1415;
  assign N2659 = N11589 & N1415;
  assign N2660 = N11591 & N1415;
  assign N2661 = N11593 & N1415;
  assign N2662 = N11595 & N1415;
  assign N2663 = N11597 & N1415;
  assign N2664 = N11599 & N1415;
  assign N2666 = ~correct_i;
  assign N2667 = ~N1896;
  assign N2668 = ~N2665;
  assign N2673 = ~N2672;
  assign N2676 = ~N2675;
  assign N2678 = ~N2677;
  assign N2681 = ~N2680;
  assign N2683 = ~N2682;
  assign N2686 = ~N2685;
  assign N2689 = ~idx_w_i[3];
  assign N2690 = N11096 & N2689;
  assign N2691 = N11098 & N2689;
  assign N2692 = N11100 & N2689;
  assign N2693 = N11102 & N2689;
  assign N2694 = N11097 & N2689;
  assign N2695 = N11099 & N2689;
  assign N2696 = N11101 & N2689;
  assign N2697 = N11103 & N2689;
  assign N2698 = ~idx_w_i[4];
  assign N2699 = N2690 & N2698;
  assign N2700 = N2690 & idx_w_i[4];
  assign N2701 = N2691 & N2698;
  assign N2702 = N2691 & idx_w_i[4];
  assign N2703 = N2692 & N2698;
  assign N2704 = N2692 & idx_w_i[4];
  assign N2705 = N2693 & N2698;
  assign N2706 = N2693 & idx_w_i[4];
  assign N2707 = N2694 & N2698;
  assign N2708 = N2694 & idx_w_i[4];
  assign N2709 = N2695 & N2698;
  assign N2710 = N2695 & idx_w_i[4];
  assign N2711 = N2696 & N2698;
  assign N2712 = N2696 & idx_w_i[4];
  assign N2713 = N2697 & N2698;
  assign N2714 = N2697 & idx_w_i[4];
  assign N2715 = N11105 & N2698;
  assign N2716 = N11107 & N2698;
  assign N2717 = N11109 & N2698;
  assign N2718 = N11111 & N2698;
  assign N2719 = N11113 & N2698;
  assign N2720 = N11115 & N2698;
  assign N2721 = N11117 & N2698;
  assign N2722 = N11119 & N2698;
  assign N2723 = N2699 & N1060;
  assign N2724 = N2699 & idx_w_i[5];
  assign N2725 = N2701 & N1060;
  assign N2726 = N2701 & idx_w_i[5];
  assign N2727 = N2703 & N1060;
  assign N2728 = N2703 & idx_w_i[5];
  assign N2729 = N2705 & N1060;
  assign N2730 = N2705 & idx_w_i[5];
  assign N2731 = N2707 & N1060;
  assign N2732 = N2707 & idx_w_i[5];
  assign N2733 = N2709 & N1060;
  assign N2734 = N2709 & idx_w_i[5];
  assign N2735 = N2711 & N1060;
  assign N2736 = N2711 & idx_w_i[5];
  assign N2737 = N2713 & N1060;
  assign N2738 = N2713 & idx_w_i[5];
  assign N2739 = N2715 & N1060;
  assign N2740 = N2715 & idx_w_i[5];
  assign N2741 = N2716 & N1060;
  assign N2742 = N2716 & idx_w_i[5];
  assign N2743 = N2717 & N1060;
  assign N2744 = N2717 & idx_w_i[5];
  assign N2745 = N2718 & N1060;
  assign N2746 = N2718 & idx_w_i[5];
  assign N2747 = N2719 & N1060;
  assign N2748 = N2719 & idx_w_i[5];
  assign N2749 = N2720 & N1060;
  assign N2750 = N2720 & idx_w_i[5];
  assign N2751 = N2721 & N1060;
  assign N2752 = N2721 & idx_w_i[5];
  assign N2753 = N2722 & N1060;
  assign N2754 = N2722 & idx_w_i[5];
  assign N2755 = N2700 & N1060;
  assign N2756 = N2700 & idx_w_i[5];
  assign N2757 = N2702 & N1060;
  assign N2758 = N2702 & idx_w_i[5];
  assign N2759 = N2704 & N1060;
  assign N2760 = N2704 & idx_w_i[5];
  assign N2761 = N2706 & N1060;
  assign N2762 = N2706 & idx_w_i[5];
  assign N2763 = N2708 & N1060;
  assign N2764 = N2708 & idx_w_i[5];
  assign N2765 = N2710 & N1060;
  assign N2766 = N2710 & idx_w_i[5];
  assign N2767 = N2712 & N1060;
  assign N2768 = N2712 & idx_w_i[5];
  assign N2769 = N2714 & N1060;
  assign N2770 = N2714 & idx_w_i[5];
  assign N2771 = N11137 & N1060;
  assign N2772 = N11139 & N1060;
  assign N2773 = N11141 & N1060;
  assign N2774 = N11143 & N1060;
  assign N2775 = N11145 & N1060;
  assign N2776 = N11147 & N1060;
  assign N2777 = N11149 & N1060;
  assign N2778 = N11151 & N1060;
  assign N2779 = N2723 & N1093;
  assign N2780 = N2723 & idx_w_i[6];
  assign N2781 = N2725 & N1093;
  assign N2782 = N2725 & idx_w_i[6];
  assign N2783 = N2727 & N1093;
  assign N2784 = N2727 & idx_w_i[6];
  assign N2785 = N2729 & N1093;
  assign N2786 = N2729 & idx_w_i[6];
  assign N2787 = N2731 & N1093;
  assign N2788 = N2731 & idx_w_i[6];
  assign N2789 = N2733 & N1093;
  assign N2790 = N2733 & idx_w_i[6];
  assign N2791 = N2735 & N1093;
  assign N2792 = N2735 & idx_w_i[6];
  assign N2793 = N2737 & N1093;
  assign N2794 = N2737 & idx_w_i[6];
  assign N2795 = N2739 & N1093;
  assign N2796 = N2739 & idx_w_i[6];
  assign N2797 = N2741 & N1093;
  assign N2798 = N2741 & idx_w_i[6];
  assign N2799 = N2743 & N1093;
  assign N2800 = N2743 & idx_w_i[6];
  assign N2801 = N2745 & N1093;
  assign N2802 = N2745 & idx_w_i[6];
  assign N2803 = N2747 & N1093;
  assign N2804 = N2747 & idx_w_i[6];
  assign N2805 = N2749 & N1093;
  assign N2806 = N2749 & idx_w_i[6];
  assign N2807 = N2751 & N1093;
  assign N2808 = N2751 & idx_w_i[6];
  assign N2809 = N2753 & N1093;
  assign N2810 = N2753 & idx_w_i[6];
  assign N2811 = N2755 & N1093;
  assign N2812 = N2755 & idx_w_i[6];
  assign N2813 = N2757 & N1093;
  assign N2814 = N2757 & idx_w_i[6];
  assign N2815 = N2759 & N1093;
  assign N2816 = N2759 & idx_w_i[6];
  assign N2817 = N2761 & N1093;
  assign N2818 = N2761 & idx_w_i[6];
  assign N2819 = N2763 & N1093;
  assign N2820 = N2763 & idx_w_i[6];
  assign N2821 = N2765 & N1093;
  assign N2822 = N2765 & idx_w_i[6];
  assign N2823 = N2767 & N1093;
  assign N2824 = N2767 & idx_w_i[6];
  assign N2825 = N2769 & N1093;
  assign N2826 = N2769 & idx_w_i[6];
  assign N2827 = N2771 & N1093;
  assign N2828 = N2771 & idx_w_i[6];
  assign N2829 = N2772 & N1093;
  assign N2830 = N2772 & idx_w_i[6];
  assign N2831 = N2773 & N1093;
  assign N2832 = N2773 & idx_w_i[6];
  assign N2833 = N2774 & N1093;
  assign N2834 = N2774 & idx_w_i[6];
  assign N2835 = N2775 & N1093;
  assign N2836 = N2775 & idx_w_i[6];
  assign N2837 = N2776 & N1093;
  assign N2838 = N2776 & idx_w_i[6];
  assign N2839 = N2777 & N1093;
  assign N2840 = N2777 & idx_w_i[6];
  assign N2841 = N2778 & N1093;
  assign N2842 = N2778 & idx_w_i[6];
  assign N2843 = N2724 & N1093;
  assign N2844 = N2724 & idx_w_i[6];
  assign N2845 = N2726 & N1093;
  assign N2846 = N2726 & idx_w_i[6];
  assign N2847 = N2728 & N1093;
  assign N2848 = N2728 & idx_w_i[6];
  assign N2849 = N2730 & N1093;
  assign N2850 = N2730 & idx_w_i[6];
  assign N2851 = N2732 & N1093;
  assign N2852 = N2732 & idx_w_i[6];
  assign N2853 = N2734 & N1093;
  assign N2854 = N2734 & idx_w_i[6];
  assign N2855 = N2736 & N1093;
  assign N2856 = N2736 & idx_w_i[6];
  assign N2857 = N2738 & N1093;
  assign N2858 = N2738 & idx_w_i[6];
  assign N2859 = N2740 & N1093;
  assign N2860 = N2740 & idx_w_i[6];
  assign N2861 = N2742 & N1093;
  assign N2862 = N2742 & idx_w_i[6];
  assign N2863 = N2744 & N1093;
  assign N2864 = N2744 & idx_w_i[6];
  assign N2865 = N2746 & N1093;
  assign N2866 = N2746 & idx_w_i[6];
  assign N2867 = N2748 & N1093;
  assign N2868 = N2748 & idx_w_i[6];
  assign N2869 = N2750 & N1093;
  assign N2870 = N2750 & idx_w_i[6];
  assign N2871 = N2752 & N1093;
  assign N2872 = N2752 & idx_w_i[6];
  assign N2873 = N2754 & N1093;
  assign N2874 = N2754 & idx_w_i[6];
  assign N2875 = N2756 & N1093;
  assign N2876 = N2756 & idx_w_i[6];
  assign N2877 = N2758 & N1093;
  assign N2878 = N2758 & idx_w_i[6];
  assign N2879 = N2760 & N1093;
  assign N2880 = N2760 & idx_w_i[6];
  assign N2881 = N2762 & N1093;
  assign N2882 = N2762 & idx_w_i[6];
  assign N2883 = N2764 & N1093;
  assign N2884 = N2764 & idx_w_i[6];
  assign N2885 = N2766 & N1093;
  assign N2886 = N2766 & idx_w_i[6];
  assign N2887 = N2768 & N1093;
  assign N2888 = N2768 & idx_w_i[6];
  assign N2889 = N2770 & N1093;
  assign N2890 = N2770 & idx_w_i[6];
  assign N2891 = N11201 & N1093;
  assign N2892 = N11203 & N1093;
  assign N2893 = N11205 & N1093;
  assign N2894 = N11207 & N1093;
  assign N2895 = N11209 & N1093;
  assign N2896 = N11211 & N1093;
  assign N2897 = N11213 & N1093;
  assign N2898 = N11215 & N1093;
  assign N2899 = N2779 & N1190;
  assign N2900 = N2779 & idx_w_i[7];
  assign N2901 = N2781 & N1190;
  assign N2902 = N2781 & idx_w_i[7];
  assign N2903 = N2783 & N1190;
  assign N2904 = N2783 & idx_w_i[7];
  assign N2905 = N2785 & N1190;
  assign N2906 = N2785 & idx_w_i[7];
  assign N2907 = N2787 & N1190;
  assign N2908 = N2787 & idx_w_i[7];
  assign N2909 = N2789 & N1190;
  assign N2910 = N2789 & idx_w_i[7];
  assign N2911 = N2791 & N1190;
  assign N2912 = N2791 & idx_w_i[7];
  assign N2913 = N2793 & N1190;
  assign N2914 = N2793 & idx_w_i[7];
  assign N2915 = N2795 & N1190;
  assign N2916 = N2795 & idx_w_i[7];
  assign N2917 = N2797 & N1190;
  assign N2918 = N2797 & idx_w_i[7];
  assign N2919 = N2799 & N1190;
  assign N2920 = N2799 & idx_w_i[7];
  assign N2921 = N2801 & N1190;
  assign N2922 = N2801 & idx_w_i[7];
  assign N2923 = N2803 & N1190;
  assign N2924 = N2803 & idx_w_i[7];
  assign N2925 = N2805 & N1190;
  assign N2926 = N2805 & idx_w_i[7];
  assign N2927 = N2807 & N1190;
  assign N2928 = N2807 & idx_w_i[7];
  assign N2929 = N2809 & N1190;
  assign N2930 = N2809 & idx_w_i[7];
  assign N2931 = N2811 & N1190;
  assign N2932 = N2811 & idx_w_i[7];
  assign N2933 = N2813 & N1190;
  assign N2934 = N2813 & idx_w_i[7];
  assign N2935 = N2815 & N1190;
  assign N2936 = N2815 & idx_w_i[7];
  assign N2937 = N2817 & N1190;
  assign N2938 = N2817 & idx_w_i[7];
  assign N2939 = N2819 & N1190;
  assign N2940 = N2819 & idx_w_i[7];
  assign N2941 = N2821 & N1190;
  assign N2942 = N2821 & idx_w_i[7];
  assign N2943 = N2823 & N1190;
  assign N2944 = N2823 & idx_w_i[7];
  assign N2945 = N2825 & N1190;
  assign N2946 = N2825 & idx_w_i[7];
  assign N2947 = N2827 & N1190;
  assign N2948 = N2827 & idx_w_i[7];
  assign N2949 = N2829 & N1190;
  assign N2950 = N2829 & idx_w_i[7];
  assign N2951 = N2831 & N1190;
  assign N2952 = N2831 & idx_w_i[7];
  assign N2953 = N2833 & N1190;
  assign N2954 = N2833 & idx_w_i[7];
  assign N2955 = N2835 & N1190;
  assign N2956 = N2835 & idx_w_i[7];
  assign N2957 = N2837 & N1190;
  assign N2958 = N2837 & idx_w_i[7];
  assign N2959 = N2839 & N1190;
  assign N2960 = N2839 & idx_w_i[7];
  assign N2961 = N2841 & N1190;
  assign N2962 = N2841 & idx_w_i[7];
  assign N2963 = N2843 & N1190;
  assign N2964 = N2843 & idx_w_i[7];
  assign N2965 = N2845 & N1190;
  assign N2966 = N2845 & idx_w_i[7];
  assign N2967 = N2847 & N1190;
  assign N2968 = N2847 & idx_w_i[7];
  assign N2969 = N2849 & N1190;
  assign N2970 = N2849 & idx_w_i[7];
  assign N2971 = N2851 & N1190;
  assign N2972 = N2851 & idx_w_i[7];
  assign N2973 = N2853 & N1190;
  assign N2974 = N2853 & idx_w_i[7];
  assign N2975 = N2855 & N1190;
  assign N2976 = N2855 & idx_w_i[7];
  assign N2977 = N2857 & N1190;
  assign N2978 = N2857 & idx_w_i[7];
  assign N2979 = N2859 & N1190;
  assign N2980 = N2859 & idx_w_i[7];
  assign N2981 = N2861 & N1190;
  assign N2982 = N2861 & idx_w_i[7];
  assign N2983 = N2863 & N1190;
  assign N2984 = N2863 & idx_w_i[7];
  assign N2985 = N2865 & N1190;
  assign N2986 = N2865 & idx_w_i[7];
  assign N2987 = N2867 & N1190;
  assign N2988 = N2867 & idx_w_i[7];
  assign N2989 = N2869 & N1190;
  assign N2990 = N2869 & idx_w_i[7];
  assign N2991 = N2871 & N1190;
  assign N2992 = N2871 & idx_w_i[7];
  assign N2993 = N2873 & N1190;
  assign N2994 = N2873 & idx_w_i[7];
  assign N2995 = N2875 & N1190;
  assign N2996 = N2875 & idx_w_i[7];
  assign N2997 = N2877 & N1190;
  assign N2998 = N2877 & idx_w_i[7];
  assign N2999 = N2879 & N1190;
  assign N3000 = N2879 & idx_w_i[7];
  assign N3001 = N2881 & N1190;
  assign N3002 = N2881 & idx_w_i[7];
  assign N3003 = N2883 & N1190;
  assign N3004 = N2883 & idx_w_i[7];
  assign N3005 = N2885 & N1190;
  assign N3006 = N2885 & idx_w_i[7];
  assign N3007 = N2887 & N1190;
  assign N3008 = N2887 & idx_w_i[7];
  assign N3009 = N2889 & N1190;
  assign N3010 = N2889 & idx_w_i[7];
  assign N3011 = N2891 & N1190;
  assign N3012 = N2891 & idx_w_i[7];
  assign N3013 = N2892 & N1190;
  assign N3014 = N2892 & idx_w_i[7];
  assign N3015 = N2893 & N1190;
  assign N3016 = N2893 & idx_w_i[7];
  assign N3017 = N2894 & N1190;
  assign N3018 = N2894 & idx_w_i[7];
  assign N3019 = N2895 & N1190;
  assign N3020 = N2895 & idx_w_i[7];
  assign N3021 = N2896 & N1190;
  assign N3022 = N2896 & idx_w_i[7];
  assign N3023 = N2897 & N1190;
  assign N3024 = N2897 & idx_w_i[7];
  assign N3025 = N2898 & N1190;
  assign N3026 = N2898 & idx_w_i[7];
  assign N3027 = N2780 & N1190;
  assign N3028 = N2780 & idx_w_i[7];
  assign N3029 = N2782 & N1190;
  assign N3030 = N2782 & idx_w_i[7];
  assign N3031 = N2784 & N1190;
  assign N3032 = N2784 & idx_w_i[7];
  assign N3033 = N2786 & N1190;
  assign N3034 = N2786 & idx_w_i[7];
  assign N3035 = N2788 & N1190;
  assign N3036 = N2788 & idx_w_i[7];
  assign N3037 = N2790 & N1190;
  assign N3038 = N2790 & idx_w_i[7];
  assign N3039 = N2792 & N1190;
  assign N3040 = N2792 & idx_w_i[7];
  assign N3041 = N2794 & N1190;
  assign N3042 = N2794 & idx_w_i[7];
  assign N3043 = N2796 & N1190;
  assign N3044 = N2796 & idx_w_i[7];
  assign N3045 = N2798 & N1190;
  assign N3046 = N2798 & idx_w_i[7];
  assign N3047 = N2800 & N1190;
  assign N3048 = N2800 & idx_w_i[7];
  assign N3049 = N2802 & N1190;
  assign N3050 = N2802 & idx_w_i[7];
  assign N3051 = N2804 & N1190;
  assign N3052 = N2804 & idx_w_i[7];
  assign N3053 = N2806 & N1190;
  assign N3054 = N2806 & idx_w_i[7];
  assign N3055 = N2808 & N1190;
  assign N3056 = N2808 & idx_w_i[7];
  assign N3057 = N2810 & N1190;
  assign N3058 = N2810 & idx_w_i[7];
  assign N3059 = N2812 & N1190;
  assign N3060 = N2812 & idx_w_i[7];
  assign N3061 = N2814 & N1190;
  assign N3062 = N2814 & idx_w_i[7];
  assign N3063 = N2816 & N1190;
  assign N3064 = N2816 & idx_w_i[7];
  assign N3065 = N2818 & N1190;
  assign N3066 = N2818 & idx_w_i[7];
  assign N3067 = N2820 & N1190;
  assign N3068 = N2820 & idx_w_i[7];
  assign N3069 = N2822 & N1190;
  assign N3070 = N2822 & idx_w_i[7];
  assign N3071 = N2824 & N1190;
  assign N3072 = N2824 & idx_w_i[7];
  assign N3073 = N2826 & N1190;
  assign N3074 = N2826 & idx_w_i[7];
  assign N3075 = N2828 & N1190;
  assign N3076 = N2828 & idx_w_i[7];
  assign N3077 = N2830 & N1190;
  assign N3078 = N2830 & idx_w_i[7];
  assign N3079 = N2832 & N1190;
  assign N3080 = N2832 & idx_w_i[7];
  assign N3081 = N2834 & N1190;
  assign N3082 = N2834 & idx_w_i[7];
  assign N3083 = N2836 & N1190;
  assign N3084 = N2836 & idx_w_i[7];
  assign N3085 = N2838 & N1190;
  assign N3086 = N2838 & idx_w_i[7];
  assign N3087 = N2840 & N1190;
  assign N3088 = N2840 & idx_w_i[7];
  assign N3089 = N2842 & N1190;
  assign N3090 = N2842 & idx_w_i[7];
  assign N3091 = N2844 & N1190;
  assign N3092 = N2844 & idx_w_i[7];
  assign N3093 = N2846 & N1190;
  assign N3094 = N2846 & idx_w_i[7];
  assign N3095 = N2848 & N1190;
  assign N3096 = N2848 & idx_w_i[7];
  assign N3097 = N2850 & N1190;
  assign N3098 = N2850 & idx_w_i[7];
  assign N3099 = N2852 & N1190;
  assign N3100 = N2852 & idx_w_i[7];
  assign N3101 = N2854 & N1190;
  assign N3102 = N2854 & idx_w_i[7];
  assign N3103 = N2856 & N1190;
  assign N3104 = N2856 & idx_w_i[7];
  assign N3105 = N2858 & N1190;
  assign N3106 = N2858 & idx_w_i[7];
  assign N3107 = N2860 & N1190;
  assign N3108 = N2860 & idx_w_i[7];
  assign N3109 = N2862 & N1190;
  assign N3110 = N2862 & idx_w_i[7];
  assign N3111 = N2864 & N1190;
  assign N3112 = N2864 & idx_w_i[7];
  assign N3113 = N2866 & N1190;
  assign N3114 = N2866 & idx_w_i[7];
  assign N3115 = N2868 & N1190;
  assign N3116 = N2868 & idx_w_i[7];
  assign N3117 = N2870 & N1190;
  assign N3118 = N2870 & idx_w_i[7];
  assign N3119 = N2872 & N1190;
  assign N3120 = N2872 & idx_w_i[7];
  assign N3121 = N2874 & N1190;
  assign N3122 = N2874 & idx_w_i[7];
  assign N3123 = N2876 & N1190;
  assign N3124 = N2876 & idx_w_i[7];
  assign N3125 = N2878 & N1190;
  assign N3126 = N2878 & idx_w_i[7];
  assign N3127 = N2880 & N1190;
  assign N3128 = N2880 & idx_w_i[7];
  assign N3129 = N2882 & N1190;
  assign N3130 = N2882 & idx_w_i[7];
  assign N3131 = N2884 & N1190;
  assign N3132 = N2884 & idx_w_i[7];
  assign N3133 = N2886 & N1190;
  assign N3134 = N2886 & idx_w_i[7];
  assign N3135 = N2888 & N1190;
  assign N3136 = N2888 & idx_w_i[7];
  assign N3137 = N2890 & N1190;
  assign N3138 = N2890 & idx_w_i[7];
  assign N3139 = N11329 & N1190;
  assign N3140 = N11331 & N1190;
  assign N3141 = N11333 & N1190;
  assign N3142 = N11335 & N1190;
  assign N3143 = N11337 & N1190;
  assign N3144 = N11339 & N1190;
  assign N3145 = N11341 & N1190;
  assign N3146 = N11343 & N1190;
  assign N3147 = N2899 & N1415;
  assign N3148 = N2899 & idx_w_i[8];
  assign N3149 = N2901 & N1415;
  assign N3150 = N2901 & idx_w_i[8];
  assign N3151 = N2903 & N1415;
  assign N3152 = N2903 & idx_w_i[8];
  assign N3153 = N2905 & N1415;
  assign N3154 = N2905 & idx_w_i[8];
  assign N3155 = N2907 & N1415;
  assign N3156 = N2907 & idx_w_i[8];
  assign N3157 = N2909 & N1415;
  assign N3158 = N2909 & idx_w_i[8];
  assign N3159 = N2911 & N1415;
  assign N3160 = N2911 & idx_w_i[8];
  assign N3161 = N2913 & N1415;
  assign N3162 = N2913 & idx_w_i[8];
  assign N3163 = N2915 & N1415;
  assign N3164 = N2915 & idx_w_i[8];
  assign N3165 = N2917 & N1415;
  assign N3166 = N2917 & idx_w_i[8];
  assign N3167 = N2919 & N1415;
  assign N3168 = N2919 & idx_w_i[8];
  assign N3169 = N2921 & N1415;
  assign N3170 = N2921 & idx_w_i[8];
  assign N3171 = N2923 & N1415;
  assign N3172 = N2923 & idx_w_i[8];
  assign N3173 = N2925 & N1415;
  assign N3174 = N2925 & idx_w_i[8];
  assign N3175 = N2927 & N1415;
  assign N3176 = N2927 & idx_w_i[8];
  assign N3177 = N2929 & N1415;
  assign N3178 = N2929 & idx_w_i[8];
  assign N3179 = N2931 & N1415;
  assign N3180 = N2931 & idx_w_i[8];
  assign N3181 = N2933 & N1415;
  assign N3182 = N2933 & idx_w_i[8];
  assign N3183 = N2935 & N1415;
  assign N3184 = N2935 & idx_w_i[8];
  assign N3185 = N2937 & N1415;
  assign N3186 = N2937 & idx_w_i[8];
  assign N3187 = N2939 & N1415;
  assign N3188 = N2939 & idx_w_i[8];
  assign N3189 = N2941 & N1415;
  assign N3190 = N2941 & idx_w_i[8];
  assign N3191 = N2943 & N1415;
  assign N3192 = N2943 & idx_w_i[8];
  assign N3193 = N2945 & N1415;
  assign N3194 = N2945 & idx_w_i[8];
  assign N3195 = N2947 & N1415;
  assign N3196 = N2947 & idx_w_i[8];
  assign N3197 = N2949 & N1415;
  assign N3198 = N2949 & idx_w_i[8];
  assign N3199 = N2951 & N1415;
  assign N3200 = N2951 & idx_w_i[8];
  assign N3201 = N2953 & N1415;
  assign N3202 = N2953 & idx_w_i[8];
  assign N3203 = N2955 & N1415;
  assign N3204 = N2955 & idx_w_i[8];
  assign N3205 = N2957 & N1415;
  assign N3206 = N2957 & idx_w_i[8];
  assign N3207 = N2959 & N1415;
  assign N3208 = N2959 & idx_w_i[8];
  assign N3209 = N2961 & N1415;
  assign N3210 = N2961 & idx_w_i[8];
  assign N3211 = N2963 & N1415;
  assign N3212 = N2963 & idx_w_i[8];
  assign N3213 = N2965 & N1415;
  assign N3214 = N2965 & idx_w_i[8];
  assign N3215 = N2967 & N1415;
  assign N3216 = N2967 & idx_w_i[8];
  assign N3217 = N2969 & N1415;
  assign N3218 = N2969 & idx_w_i[8];
  assign N3219 = N2971 & N1415;
  assign N3220 = N2971 & idx_w_i[8];
  assign N3221 = N2973 & N1415;
  assign N3222 = N2973 & idx_w_i[8];
  assign N3223 = N2975 & N1415;
  assign N3224 = N2975 & idx_w_i[8];
  assign N3225 = N2977 & N1415;
  assign N3226 = N2977 & idx_w_i[8];
  assign N3227 = N2979 & N1415;
  assign N3228 = N2979 & idx_w_i[8];
  assign N3229 = N2981 & N1415;
  assign N3230 = N2981 & idx_w_i[8];
  assign N3231 = N2983 & N1415;
  assign N3232 = N2983 & idx_w_i[8];
  assign N3233 = N2985 & N1415;
  assign N3234 = N2985 & idx_w_i[8];
  assign N3235 = N2987 & N1415;
  assign N3236 = N2987 & idx_w_i[8];
  assign N3237 = N2989 & N1415;
  assign N3238 = N2989 & idx_w_i[8];
  assign N3239 = N2991 & N1415;
  assign N3240 = N2991 & idx_w_i[8];
  assign N3241 = N2993 & N1415;
  assign N3242 = N2993 & idx_w_i[8];
  assign N3243 = N2995 & N1415;
  assign N3244 = N2995 & idx_w_i[8];
  assign N3245 = N2997 & N1415;
  assign N3246 = N2997 & idx_w_i[8];
  assign N3247 = N2999 & N1415;
  assign N3248 = N2999 & idx_w_i[8];
  assign N3249 = N3001 & N1415;
  assign N3250 = N3001 & idx_w_i[8];
  assign N3251 = N3003 & N1415;
  assign N3252 = N3003 & idx_w_i[8];
  assign N3253 = N3005 & N1415;
  assign N3254 = N3005 & idx_w_i[8];
  assign N3255 = N3007 & N1415;
  assign N3256 = N3007 & idx_w_i[8];
  assign N3257 = N3009 & N1415;
  assign N3258 = N3009 & idx_w_i[8];
  assign N3259 = N3011 & N1415;
  assign N3260 = N3011 & idx_w_i[8];
  assign N3261 = N3013 & N1415;
  assign N3262 = N3013 & idx_w_i[8];
  assign N3263 = N3015 & N1415;
  assign N3264 = N3015 & idx_w_i[8];
  assign N3265 = N3017 & N1415;
  assign N3266 = N3017 & idx_w_i[8];
  assign N3267 = N3019 & N1415;
  assign N3268 = N3019 & idx_w_i[8];
  assign N3269 = N3021 & N1415;
  assign N3270 = N3021 & idx_w_i[8];
  assign N3271 = N3023 & N1415;
  assign N3272 = N3023 & idx_w_i[8];
  assign N3273 = N3025 & N1415;
  assign N3274 = N3025 & idx_w_i[8];
  assign N3275 = N3027 & N1415;
  assign N3276 = N3027 & idx_w_i[8];
  assign N3277 = N3029 & N1415;
  assign N3278 = N3029 & idx_w_i[8];
  assign N3279 = N3031 & N1415;
  assign N3280 = N3031 & idx_w_i[8];
  assign N3281 = N3033 & N1415;
  assign N3282 = N3033 & idx_w_i[8];
  assign N3283 = N3035 & N1415;
  assign N3284 = N3035 & idx_w_i[8];
  assign N3285 = N3037 & N1415;
  assign N3286 = N3037 & idx_w_i[8];
  assign N3287 = N3039 & N1415;
  assign N3288 = N3039 & idx_w_i[8];
  assign N3289 = N3041 & N1415;
  assign N3290 = N3041 & idx_w_i[8];
  assign N3291 = N3043 & N1415;
  assign N3292 = N3043 & idx_w_i[8];
  assign N3293 = N3045 & N1415;
  assign N3294 = N3045 & idx_w_i[8];
  assign N3295 = N3047 & N1415;
  assign N3296 = N3047 & idx_w_i[8];
  assign N3297 = N3049 & N1415;
  assign N3298 = N3049 & idx_w_i[8];
  assign N3299 = N3051 & N1415;
  assign N3300 = N3051 & idx_w_i[8];
  assign N3301 = N3053 & N1415;
  assign N3302 = N3053 & idx_w_i[8];
  assign N3303 = N3055 & N1415;
  assign N3304 = N3055 & idx_w_i[8];
  assign N3305 = N3057 & N1415;
  assign N3306 = N3057 & idx_w_i[8];
  assign N3307 = N3059 & N1415;
  assign N3308 = N3059 & idx_w_i[8];
  assign N3309 = N3061 & N1415;
  assign N3310 = N3061 & idx_w_i[8];
  assign N3311 = N3063 & N1415;
  assign N3312 = N3063 & idx_w_i[8];
  assign N3313 = N3065 & N1415;
  assign N3314 = N3065 & idx_w_i[8];
  assign N3315 = N3067 & N1415;
  assign N3316 = N3067 & idx_w_i[8];
  assign N3317 = N3069 & N1415;
  assign N3318 = N3069 & idx_w_i[8];
  assign N3319 = N3071 & N1415;
  assign N3320 = N3071 & idx_w_i[8];
  assign N3321 = N3073 & N1415;
  assign N3322 = N3073 & idx_w_i[8];
  assign N3323 = N3075 & N1415;
  assign N3324 = N3075 & idx_w_i[8];
  assign N3325 = N3077 & N1415;
  assign N3326 = N3077 & idx_w_i[8];
  assign N3327 = N3079 & N1415;
  assign N3328 = N3079 & idx_w_i[8];
  assign N3329 = N3081 & N1415;
  assign N3330 = N3081 & idx_w_i[8];
  assign N3331 = N3083 & N1415;
  assign N3332 = N3083 & idx_w_i[8];
  assign N3333 = N3085 & N1415;
  assign N3334 = N3085 & idx_w_i[8];
  assign N3335 = N3087 & N1415;
  assign N3336 = N3087 & idx_w_i[8];
  assign N3337 = N3089 & N1415;
  assign N3338 = N3089 & idx_w_i[8];
  assign N3339 = N3091 & N1415;
  assign N3340 = N3091 & idx_w_i[8];
  assign N3341 = N3093 & N1415;
  assign N3342 = N3093 & idx_w_i[8];
  assign N3343 = N3095 & N1415;
  assign N3344 = N3095 & idx_w_i[8];
  assign N3345 = N3097 & N1415;
  assign N3346 = N3097 & idx_w_i[8];
  assign N3347 = N3099 & N1415;
  assign N3348 = N3099 & idx_w_i[8];
  assign N3349 = N3101 & N1415;
  assign N3350 = N3101 & idx_w_i[8];
  assign N3351 = N3103 & N1415;
  assign N3352 = N3103 & idx_w_i[8];
  assign N3353 = N3105 & N1415;
  assign N3354 = N3105 & idx_w_i[8];
  assign N3355 = N3107 & N1415;
  assign N3356 = N3107 & idx_w_i[8];
  assign N3357 = N3109 & N1415;
  assign N3358 = N3109 & idx_w_i[8];
  assign N3359 = N3111 & N1415;
  assign N3360 = N3111 & idx_w_i[8];
  assign N3361 = N3113 & N1415;
  assign N3362 = N3113 & idx_w_i[8];
  assign N3363 = N3115 & N1415;
  assign N3364 = N3115 & idx_w_i[8];
  assign N3365 = N3117 & N1415;
  assign N3366 = N3117 & idx_w_i[8];
  assign N3367 = N3119 & N1415;
  assign N3368 = N3119 & idx_w_i[8];
  assign N3369 = N3121 & N1415;
  assign N3370 = N3121 & idx_w_i[8];
  assign N3371 = N3123 & N1415;
  assign N3372 = N3123 & idx_w_i[8];
  assign N3373 = N3125 & N1415;
  assign N3374 = N3125 & idx_w_i[8];
  assign N3375 = N3127 & N1415;
  assign N3376 = N3127 & idx_w_i[8];
  assign N3377 = N3129 & N1415;
  assign N3378 = N3129 & idx_w_i[8];
  assign N3379 = N3131 & N1415;
  assign N3380 = N3131 & idx_w_i[8];
  assign N3381 = N3133 & N1415;
  assign N3382 = N3133 & idx_w_i[8];
  assign N3383 = N3135 & N1415;
  assign N3384 = N3135 & idx_w_i[8];
  assign N3385 = N3137 & N1415;
  assign N3386 = N3137 & idx_w_i[8];
  assign N3387 = N3139 & N1415;
  assign N3388 = N3139 & idx_w_i[8];
  assign N3389 = N3140 & N1415;
  assign N3390 = N3140 & idx_w_i[8];
  assign N3391 = N3141 & N1415;
  assign N3392 = N3141 & idx_w_i[8];
  assign N3393 = N3142 & N1415;
  assign N3394 = N3142 & idx_w_i[8];
  assign N3395 = N3143 & N1415;
  assign N3396 = N3143 & idx_w_i[8];
  assign N3397 = N3144 & N1415;
  assign N3398 = N3144 & idx_w_i[8];
  assign N3399 = N3145 & N1415;
  assign N3400 = N3145 & idx_w_i[8];
  assign N3401 = N3146 & N1415;
  assign N3402 = N3146 & idx_w_i[8];
  assign N3403 = N2900 & N1415;
  assign N3404 = N2900 & idx_w_i[8];
  assign N3405 = N2902 & N1415;
  assign N3406 = N2902 & idx_w_i[8];
  assign N3407 = N2904 & N1415;
  assign N3408 = N2904 & idx_w_i[8];
  assign N3409 = N2906 & N1415;
  assign N3410 = N2906 & idx_w_i[8];
  assign N3411 = N2908 & N1415;
  assign N3412 = N2908 & idx_w_i[8];
  assign N3413 = N2910 & N1415;
  assign N3414 = N2910 & idx_w_i[8];
  assign N3415 = N2912 & N1415;
  assign N3416 = N2912 & idx_w_i[8];
  assign N3417 = N2914 & N1415;
  assign N3418 = N2914 & idx_w_i[8];
  assign N3419 = N2916 & N1415;
  assign N3420 = N2916 & idx_w_i[8];
  assign N3421 = N2918 & N1415;
  assign N3422 = N2918 & idx_w_i[8];
  assign N3423 = N2920 & N1415;
  assign N3424 = N2920 & idx_w_i[8];
  assign N3425 = N2922 & N1415;
  assign N3426 = N2922 & idx_w_i[8];
  assign N3427 = N2924 & N1415;
  assign N3428 = N2924 & idx_w_i[8];
  assign N3429 = N2926 & N1415;
  assign N3430 = N2926 & idx_w_i[8];
  assign N3431 = N2928 & N1415;
  assign N3432 = N2928 & idx_w_i[8];
  assign N3433 = N2930 & N1415;
  assign N3434 = N2930 & idx_w_i[8];
  assign N3435 = N2932 & N1415;
  assign N3436 = N2932 & idx_w_i[8];
  assign N3437 = N2934 & N1415;
  assign N3438 = N2934 & idx_w_i[8];
  assign N3439 = N2936 & N1415;
  assign N3440 = N2936 & idx_w_i[8];
  assign N3441 = N2938 & N1415;
  assign N3442 = N2938 & idx_w_i[8];
  assign N3443 = N2940 & N1415;
  assign N3444 = N2940 & idx_w_i[8];
  assign N3445 = N2942 & N1415;
  assign N3446 = N2942 & idx_w_i[8];
  assign N3447 = N2944 & N1415;
  assign N3448 = N2944 & idx_w_i[8];
  assign N3449 = N2946 & N1415;
  assign N3450 = N2946 & idx_w_i[8];
  assign N3451 = N2948 & N1415;
  assign N3452 = N2948 & idx_w_i[8];
  assign N3453 = N2950 & N1415;
  assign N3454 = N2950 & idx_w_i[8];
  assign N3455 = N2952 & N1415;
  assign N3456 = N2952 & idx_w_i[8];
  assign N3457 = N2954 & N1415;
  assign N3458 = N2954 & idx_w_i[8];
  assign N3459 = N2956 & N1415;
  assign N3460 = N2956 & idx_w_i[8];
  assign N3461 = N2958 & N1415;
  assign N3462 = N2958 & idx_w_i[8];
  assign N3463 = N2960 & N1415;
  assign N3464 = N2960 & idx_w_i[8];
  assign N3465 = N2962 & N1415;
  assign N3466 = N2962 & idx_w_i[8];
  assign N3467 = N2964 & N1415;
  assign N3468 = N2964 & idx_w_i[8];
  assign N3469 = N2966 & N1415;
  assign N3470 = N2966 & idx_w_i[8];
  assign N3471 = N2968 & N1415;
  assign N3472 = N2968 & idx_w_i[8];
  assign N3473 = N2970 & N1415;
  assign N3474 = N2970 & idx_w_i[8];
  assign N3475 = N2972 & N1415;
  assign N3476 = N2972 & idx_w_i[8];
  assign N3477 = N2974 & N1415;
  assign N3478 = N2974 & idx_w_i[8];
  assign N3479 = N2976 & N1415;
  assign N3480 = N2976 & idx_w_i[8];
  assign N3481 = N2978 & N1415;
  assign N3482 = N2978 & idx_w_i[8];
  assign N3483 = N2980 & N1415;
  assign N3484 = N2980 & idx_w_i[8];
  assign N3485 = N2982 & N1415;
  assign N3486 = N2982 & idx_w_i[8];
  assign N3487 = N2984 & N1415;
  assign N3488 = N2984 & idx_w_i[8];
  assign N3489 = N2986 & N1415;
  assign N3490 = N2986 & idx_w_i[8];
  assign N3491 = N2988 & N1415;
  assign N3492 = N2988 & idx_w_i[8];
  assign N3493 = N2990 & N1415;
  assign N3494 = N2990 & idx_w_i[8];
  assign N3495 = N2992 & N1415;
  assign N3496 = N2992 & idx_w_i[8];
  assign N3497 = N2994 & N1415;
  assign N3498 = N2994 & idx_w_i[8];
  assign N3499 = N2996 & N1415;
  assign N3500 = N2996 & idx_w_i[8];
  assign N3501 = N2998 & N1415;
  assign N3502 = N2998 & idx_w_i[8];
  assign N3503 = N3000 & N1415;
  assign N3504 = N3000 & idx_w_i[8];
  assign N3505 = N3002 & N1415;
  assign N3506 = N3002 & idx_w_i[8];
  assign N3507 = N3004 & N1415;
  assign N3508 = N3004 & idx_w_i[8];
  assign N3509 = N3006 & N1415;
  assign N3510 = N3006 & idx_w_i[8];
  assign N3511 = N3008 & N1415;
  assign N3512 = N3008 & idx_w_i[8];
  assign N3513 = N3010 & N1415;
  assign N3514 = N3010 & idx_w_i[8];
  assign N3515 = N3012 & N1415;
  assign N3516 = N3012 & idx_w_i[8];
  assign N3517 = N3014 & N1415;
  assign N3518 = N3014 & idx_w_i[8];
  assign N3519 = N3016 & N1415;
  assign N3520 = N3016 & idx_w_i[8];
  assign N3521 = N3018 & N1415;
  assign N3522 = N3018 & idx_w_i[8];
  assign N3523 = N3020 & N1415;
  assign N3524 = N3020 & idx_w_i[8];
  assign N3525 = N3022 & N1415;
  assign N3526 = N3022 & idx_w_i[8];
  assign N3527 = N3024 & N1415;
  assign N3528 = N3024 & idx_w_i[8];
  assign N3529 = N3026 & N1415;
  assign N3530 = N3026 & idx_w_i[8];
  assign N3531 = N3028 & N1415;
  assign N3532 = N3028 & idx_w_i[8];
  assign N3533 = N3030 & N1415;
  assign N3534 = N3030 & idx_w_i[8];
  assign N3535 = N3032 & N1415;
  assign N3536 = N3032 & idx_w_i[8];
  assign N3537 = N3034 & N1415;
  assign N3538 = N3034 & idx_w_i[8];
  assign N3539 = N3036 & N1415;
  assign N3540 = N3036 & idx_w_i[8];
  assign N3541 = N3038 & N1415;
  assign N3542 = N3038 & idx_w_i[8];
  assign N3543 = N3040 & N1415;
  assign N3544 = N3040 & idx_w_i[8];
  assign N3545 = N3042 & N1415;
  assign N3546 = N3042 & idx_w_i[8];
  assign N3547 = N3044 & N1415;
  assign N3548 = N3044 & idx_w_i[8];
  assign N3549 = N3046 & N1415;
  assign N3550 = N3046 & idx_w_i[8];
  assign N3551 = N3048 & N1415;
  assign N3552 = N3048 & idx_w_i[8];
  assign N3553 = N3050 & N1415;
  assign N3554 = N3050 & idx_w_i[8];
  assign N3555 = N3052 & N1415;
  assign N3556 = N3052 & idx_w_i[8];
  assign N3557 = N3054 & N1415;
  assign N3558 = N3054 & idx_w_i[8];
  assign N3559 = N3056 & N1415;
  assign N3560 = N3056 & idx_w_i[8];
  assign N3561 = N3058 & N1415;
  assign N3562 = N3058 & idx_w_i[8];
  assign N3563 = N3060 & N1415;
  assign N3564 = N3060 & idx_w_i[8];
  assign N3565 = N3062 & N1415;
  assign N3566 = N3062 & idx_w_i[8];
  assign N3567 = N3064 & N1415;
  assign N3568 = N3064 & idx_w_i[8];
  assign N3569 = N3066 & N1415;
  assign N3570 = N3066 & idx_w_i[8];
  assign N3571 = N3068 & N1415;
  assign N3572 = N3068 & idx_w_i[8];
  assign N3573 = N3070 & N1415;
  assign N3574 = N3070 & idx_w_i[8];
  assign N3575 = N3072 & N1415;
  assign N3576 = N3072 & idx_w_i[8];
  assign N3577 = N3074 & N1415;
  assign N3578 = N3074 & idx_w_i[8];
  assign N3579 = N3076 & N1415;
  assign N3580 = N3076 & idx_w_i[8];
  assign N3581 = N3078 & N1415;
  assign N3582 = N3078 & idx_w_i[8];
  assign N3583 = N3080 & N1415;
  assign N3584 = N3080 & idx_w_i[8];
  assign N3585 = N3082 & N1415;
  assign N3586 = N3082 & idx_w_i[8];
  assign N3587 = N3084 & N1415;
  assign N3588 = N3084 & idx_w_i[8];
  assign N3589 = N3086 & N1415;
  assign N3590 = N3086 & idx_w_i[8];
  assign N3591 = N3088 & N1415;
  assign N3592 = N3088 & idx_w_i[8];
  assign N3593 = N3090 & N1415;
  assign N3594 = N3090 & idx_w_i[8];
  assign N3595 = N3092 & N1415;
  assign N3596 = N3092 & idx_w_i[8];
  assign N3597 = N3094 & N1415;
  assign N3598 = N3094 & idx_w_i[8];
  assign N3599 = N3096 & N1415;
  assign N3600 = N3096 & idx_w_i[8];
  assign N3601 = N3098 & N1415;
  assign N3602 = N3098 & idx_w_i[8];
  assign N3603 = N3100 & N1415;
  assign N3604 = N3100 & idx_w_i[8];
  assign N3605 = N3102 & N1415;
  assign N3606 = N3102 & idx_w_i[8];
  assign N3607 = N3104 & N1415;
  assign N3608 = N3104 & idx_w_i[8];
  assign N3609 = N3106 & N1415;
  assign N3610 = N3106 & idx_w_i[8];
  assign N3611 = N3108 & N1415;
  assign N3612 = N3108 & idx_w_i[8];
  assign N3613 = N3110 & N1415;
  assign N3614 = N3110 & idx_w_i[8];
  assign N3615 = N3112 & N1415;
  assign N3616 = N3112 & idx_w_i[8];
  assign N3617 = N3114 & N1415;
  assign N3618 = N3114 & idx_w_i[8];
  assign N3619 = N3116 & N1415;
  assign N3620 = N3116 & idx_w_i[8];
  assign N3621 = N3118 & N1415;
  assign N3622 = N3118 & idx_w_i[8];
  assign N3623 = N3120 & N1415;
  assign N3624 = N3120 & idx_w_i[8];
  assign N3625 = N3122 & N1415;
  assign N3626 = N3122 & idx_w_i[8];
  assign N3627 = N3124 & N1415;
  assign N3628 = N3124 & idx_w_i[8];
  assign N3629 = N3126 & N1415;
  assign N3630 = N3126 & idx_w_i[8];
  assign N3631 = N3128 & N1415;
  assign N3632 = N3128 & idx_w_i[8];
  assign N3633 = N3130 & N1415;
  assign N3634 = N3130 & idx_w_i[8];
  assign N3635 = N3132 & N1415;
  assign N3636 = N3132 & idx_w_i[8];
  assign N3637 = N3134 & N1415;
  assign N3638 = N3134 & idx_w_i[8];
  assign N3639 = N3136 & N1415;
  assign N3640 = N3136 & idx_w_i[8];
  assign N3641 = N3138 & N1415;
  assign N3642 = N3138 & idx_w_i[8];
  assign N3643 = N11585 & N1415;
  assign N3644 = N11587 & N1415;
  assign N3645 = N11589 & N1415;
  assign N3646 = N11591 & N1415;
  assign N3647 = N11593 & N1415;
  assign N3648 = N11595 & N1415;
  assign N3649 = N11597 & N1415;
  assign N3650 = N11599 & N1415;
  assign N3652 = N2690 & N2698;
  assign N3653 = N2691 & N2698;
  assign N3654 = N2692 & N2698;
  assign N3655 = N2693 & N2698;
  assign N3656 = N2694 & N2698;
  assign N3657 = N2695 & N2698;
  assign N3658 = N2696 & N2698;
  assign N3659 = N2697 & N2698;
  assign N3660 = N11105 & N2698;
  assign N3661 = N11107 & N2698;
  assign N3662 = N11109 & N2698;
  assign N3663 = N11111 & N2698;
  assign N3664 = N11113 & N2698;
  assign N3665 = N11115 & N2698;
  assign N3666 = N11117 & N2698;
  assign N3667 = N11119 & N2698;
  assign N3668 = N3652 & N1060;
  assign N3669 = N3652 & idx_w_i[5];
  assign N3670 = N3653 & N1060;
  assign N3671 = N3653 & idx_w_i[5];
  assign N3672 = N3654 & N1060;
  assign N3673 = N3654 & idx_w_i[5];
  assign N3674 = N3655 & N1060;
  assign N3675 = N3655 & idx_w_i[5];
  assign N3676 = N3656 & N1060;
  assign N3677 = N3656 & idx_w_i[5];
  assign N3678 = N3657 & N1060;
  assign N3679 = N3657 & idx_w_i[5];
  assign N3680 = N3658 & N1060;
  assign N3681 = N3658 & idx_w_i[5];
  assign N3682 = N3659 & N1060;
  assign N3683 = N3659 & idx_w_i[5];
  assign N3684 = N3660 & N1060;
  assign N3685 = N3660 & idx_w_i[5];
  assign N3686 = N3661 & N1060;
  assign N3687 = N3661 & idx_w_i[5];
  assign N3688 = N3662 & N1060;
  assign N3689 = N3662 & idx_w_i[5];
  assign N3690 = N3663 & N1060;
  assign N3691 = N3663 & idx_w_i[5];
  assign N3692 = N3664 & N1060;
  assign N3693 = N3664 & idx_w_i[5];
  assign N3694 = N3665 & N1060;
  assign N3695 = N3665 & idx_w_i[5];
  assign N3696 = N3666 & N1060;
  assign N3697 = N3666 & idx_w_i[5];
  assign N3698 = N3667 & N1060;
  assign N3699 = N3667 & idx_w_i[5];
  assign N3700 = N2700 & N1060;
  assign N3701 = N2702 & N1060;
  assign N3702 = N2704 & N1060;
  assign N3703 = N2706 & N1060;
  assign N3704 = N2708 & N1060;
  assign N3705 = N2710 & N1060;
  assign N3706 = N2712 & N1060;
  assign N3707 = N2714 & N1060;
  assign N3708 = N11137 & N1060;
  assign N3709 = N11139 & N1060;
  assign N3710 = N11141 & N1060;
  assign N3711 = N11143 & N1060;
  assign N3712 = N11145 & N1060;
  assign N3713 = N11147 & N1060;
  assign N3714 = N11149 & N1060;
  assign N3715 = N11151 & N1060;
  assign N3716 = N3668 & N1093;
  assign N3717 = N3668 & idx_w_i[6];
  assign N3718 = N3670 & N1093;
  assign N3719 = N3670 & idx_w_i[6];
  assign N3720 = N3672 & N1093;
  assign N3721 = N3672 & idx_w_i[6];
  assign N3722 = N3674 & N1093;
  assign N3723 = N3674 & idx_w_i[6];
  assign N3724 = N3676 & N1093;
  assign N3725 = N3676 & idx_w_i[6];
  assign N3726 = N3678 & N1093;
  assign N3727 = N3678 & idx_w_i[6];
  assign N3728 = N3680 & N1093;
  assign N3729 = N3680 & idx_w_i[6];
  assign N3730 = N3682 & N1093;
  assign N3731 = N3682 & idx_w_i[6];
  assign N3732 = N3684 & N1093;
  assign N3733 = N3684 & idx_w_i[6];
  assign N3734 = N3686 & N1093;
  assign N3735 = N3686 & idx_w_i[6];
  assign N3736 = N3688 & N1093;
  assign N3737 = N3688 & idx_w_i[6];
  assign N3738 = N3690 & N1093;
  assign N3739 = N3690 & idx_w_i[6];
  assign N3740 = N3692 & N1093;
  assign N3741 = N3692 & idx_w_i[6];
  assign N3742 = N3694 & N1093;
  assign N3743 = N3694 & idx_w_i[6];
  assign N3744 = N3696 & N1093;
  assign N3745 = N3696 & idx_w_i[6];
  assign N3746 = N3698 & N1093;
  assign N3747 = N3698 & idx_w_i[6];
  assign N3748 = N3700 & N1093;
  assign N3749 = N3700 & idx_w_i[6];
  assign N3750 = N3701 & N1093;
  assign N3751 = N3701 & idx_w_i[6];
  assign N3752 = N3702 & N1093;
  assign N3753 = N3702 & idx_w_i[6];
  assign N3754 = N3703 & N1093;
  assign N3755 = N3703 & idx_w_i[6];
  assign N3756 = N3704 & N1093;
  assign N3757 = N3704 & idx_w_i[6];
  assign N3758 = N3705 & N1093;
  assign N3759 = N3705 & idx_w_i[6];
  assign N3760 = N3706 & N1093;
  assign N3761 = N3706 & idx_w_i[6];
  assign N3762 = N3707 & N1093;
  assign N3763 = N3707 & idx_w_i[6];
  assign N3764 = N3708 & N1093;
  assign N3765 = N3708 & idx_w_i[6];
  assign N3766 = N3709 & N1093;
  assign N3767 = N3709 & idx_w_i[6];
  assign N3768 = N3710 & N1093;
  assign N3769 = N3710 & idx_w_i[6];
  assign N3770 = N3711 & N1093;
  assign N3771 = N3711 & idx_w_i[6];
  assign N3772 = N3712 & N1093;
  assign N3773 = N3712 & idx_w_i[6];
  assign N3774 = N3713 & N1093;
  assign N3775 = N3713 & idx_w_i[6];
  assign N3776 = N3714 & N1093;
  assign N3777 = N3714 & idx_w_i[6];
  assign N3778 = N3715 & N1093;
  assign N3779 = N3715 & idx_w_i[6];
  assign N3780 = N3669 & N1093;
  assign N3781 = N3669 & idx_w_i[6];
  assign N3782 = N3671 & N1093;
  assign N3783 = N3671 & idx_w_i[6];
  assign N3784 = N3673 & N1093;
  assign N3785 = N3673 & idx_w_i[6];
  assign N3786 = N3675 & N1093;
  assign N3787 = N3675 & idx_w_i[6];
  assign N3788 = N3677 & N1093;
  assign N3789 = N3677 & idx_w_i[6];
  assign N3790 = N3679 & N1093;
  assign N3791 = N3679 & idx_w_i[6];
  assign N3792 = N3681 & N1093;
  assign N3793 = N3681 & idx_w_i[6];
  assign N3794 = N3683 & N1093;
  assign N3795 = N3683 & idx_w_i[6];
  assign N3796 = N3685 & N1093;
  assign N3797 = N3685 & idx_w_i[6];
  assign N3798 = N3687 & N1093;
  assign N3799 = N3687 & idx_w_i[6];
  assign N3800 = N3689 & N1093;
  assign N3801 = N3689 & idx_w_i[6];
  assign N3802 = N3691 & N1093;
  assign N3803 = N3691 & idx_w_i[6];
  assign N3804 = N3693 & N1093;
  assign N3805 = N3693 & idx_w_i[6];
  assign N3806 = N3695 & N1093;
  assign N3807 = N3695 & idx_w_i[6];
  assign N3808 = N3697 & N1093;
  assign N3809 = N3697 & idx_w_i[6];
  assign N3810 = N3699 & N1093;
  assign N3811 = N3699 & idx_w_i[6];
  assign N3812 = N2756 & N1093;
  assign N3813 = N2758 & N1093;
  assign N3814 = N2760 & N1093;
  assign N3815 = N2762 & N1093;
  assign N3816 = N2764 & N1093;
  assign N3817 = N2766 & N1093;
  assign N3818 = N2768 & N1093;
  assign N3819 = N2770 & N1093;
  assign N3820 = N11201 & N1093;
  assign N3821 = N11203 & N1093;
  assign N3822 = N11205 & N1093;
  assign N3823 = N11207 & N1093;
  assign N3824 = N11209 & N1093;
  assign N3825 = N11211 & N1093;
  assign N3826 = N11213 & N1093;
  assign N3827 = N11215 & N1093;
  assign N3828 = N3716 & N1190;
  assign N3829 = N3716 & idx_w_i[7];
  assign N3830 = N3718 & N1190;
  assign N3831 = N3718 & idx_w_i[7];
  assign N3832 = N3720 & N1190;
  assign N3833 = N3720 & idx_w_i[7];
  assign N3834 = N3722 & N1190;
  assign N3835 = N3722 & idx_w_i[7];
  assign N3836 = N3724 & N1190;
  assign N3837 = N3724 & idx_w_i[7];
  assign N3838 = N3726 & N1190;
  assign N3839 = N3726 & idx_w_i[7];
  assign N3840 = N3728 & N1190;
  assign N3841 = N3728 & idx_w_i[7];
  assign N3842 = N3730 & N1190;
  assign N3843 = N3730 & idx_w_i[7];
  assign N3844 = N3732 & N1190;
  assign N3845 = N3732 & idx_w_i[7];
  assign N3846 = N3734 & N1190;
  assign N3847 = N3734 & idx_w_i[7];
  assign N3848 = N3736 & N1190;
  assign N3849 = N3736 & idx_w_i[7];
  assign N3850 = N3738 & N1190;
  assign N3851 = N3738 & idx_w_i[7];
  assign N3852 = N3740 & N1190;
  assign N3853 = N3740 & idx_w_i[7];
  assign N3854 = N3742 & N1190;
  assign N3855 = N3742 & idx_w_i[7];
  assign N3856 = N3744 & N1190;
  assign N3857 = N3744 & idx_w_i[7];
  assign N3858 = N3746 & N1190;
  assign N3859 = N3746 & idx_w_i[7];
  assign N3860 = N3748 & N1190;
  assign N3861 = N3748 & idx_w_i[7];
  assign N3862 = N3750 & N1190;
  assign N3863 = N3750 & idx_w_i[7];
  assign N3864 = N3752 & N1190;
  assign N3865 = N3752 & idx_w_i[7];
  assign N3866 = N3754 & N1190;
  assign N3867 = N3754 & idx_w_i[7];
  assign N3868 = N3756 & N1190;
  assign N3869 = N3756 & idx_w_i[7];
  assign N3870 = N3758 & N1190;
  assign N3871 = N3758 & idx_w_i[7];
  assign N3872 = N3760 & N1190;
  assign N3873 = N3760 & idx_w_i[7];
  assign N3874 = N3762 & N1190;
  assign N3875 = N3762 & idx_w_i[7];
  assign N3876 = N3764 & N1190;
  assign N3877 = N3764 & idx_w_i[7];
  assign N3878 = N3766 & N1190;
  assign N3879 = N3766 & idx_w_i[7];
  assign N3880 = N3768 & N1190;
  assign N3881 = N3768 & idx_w_i[7];
  assign N3882 = N3770 & N1190;
  assign N3883 = N3770 & idx_w_i[7];
  assign N3884 = N3772 & N1190;
  assign N3885 = N3772 & idx_w_i[7];
  assign N3886 = N3774 & N1190;
  assign N3887 = N3774 & idx_w_i[7];
  assign N3888 = N3776 & N1190;
  assign N3889 = N3776 & idx_w_i[7];
  assign N3890 = N3778 & N1190;
  assign N3891 = N3778 & idx_w_i[7];
  assign N3892 = N3780 & N1190;
  assign N3893 = N3780 & idx_w_i[7];
  assign N3894 = N3782 & N1190;
  assign N3895 = N3782 & idx_w_i[7];
  assign N3896 = N3784 & N1190;
  assign N3897 = N3784 & idx_w_i[7];
  assign N3898 = N3786 & N1190;
  assign N3899 = N3786 & idx_w_i[7];
  assign N3900 = N3788 & N1190;
  assign N3901 = N3788 & idx_w_i[7];
  assign N3902 = N3790 & N1190;
  assign N3903 = N3790 & idx_w_i[7];
  assign N3904 = N3792 & N1190;
  assign N3905 = N3792 & idx_w_i[7];
  assign N3906 = N3794 & N1190;
  assign N3907 = N3794 & idx_w_i[7];
  assign N3908 = N3796 & N1190;
  assign N3909 = N3796 & idx_w_i[7];
  assign N3910 = N3798 & N1190;
  assign N3911 = N3798 & idx_w_i[7];
  assign N3912 = N3800 & N1190;
  assign N3913 = N3800 & idx_w_i[7];
  assign N3914 = N3802 & N1190;
  assign N3915 = N3802 & idx_w_i[7];
  assign N3916 = N3804 & N1190;
  assign N3917 = N3804 & idx_w_i[7];
  assign N3918 = N3806 & N1190;
  assign N3919 = N3806 & idx_w_i[7];
  assign N3920 = N3808 & N1190;
  assign N3921 = N3808 & idx_w_i[7];
  assign N3922 = N3810 & N1190;
  assign N3923 = N3810 & idx_w_i[7];
  assign N3924 = N3812 & N1190;
  assign N3925 = N3812 & idx_w_i[7];
  assign N3926 = N3813 & N1190;
  assign N3927 = N3813 & idx_w_i[7];
  assign N3928 = N3814 & N1190;
  assign N3929 = N3814 & idx_w_i[7];
  assign N3930 = N3815 & N1190;
  assign N3931 = N3815 & idx_w_i[7];
  assign N3932 = N3816 & N1190;
  assign N3933 = N3816 & idx_w_i[7];
  assign N3934 = N3817 & N1190;
  assign N3935 = N3817 & idx_w_i[7];
  assign N3936 = N3818 & N1190;
  assign N3937 = N3818 & idx_w_i[7];
  assign N3938 = N3819 & N1190;
  assign N3939 = N3819 & idx_w_i[7];
  assign N3940 = N3820 & N1190;
  assign N3941 = N3820 & idx_w_i[7];
  assign N3942 = N3821 & N1190;
  assign N3943 = N3821 & idx_w_i[7];
  assign N3944 = N3822 & N1190;
  assign N3945 = N3822 & idx_w_i[7];
  assign N3946 = N3823 & N1190;
  assign N3947 = N3823 & idx_w_i[7];
  assign N3948 = N3824 & N1190;
  assign N3949 = N3824 & idx_w_i[7];
  assign N3950 = N3825 & N1190;
  assign N3951 = N3825 & idx_w_i[7];
  assign N3952 = N3826 & N1190;
  assign N3953 = N3826 & idx_w_i[7];
  assign N3954 = N3827 & N1190;
  assign N3955 = N3827 & idx_w_i[7];
  assign N3956 = N3717 & N1190;
  assign N3957 = N3717 & idx_w_i[7];
  assign N3958 = N3719 & N1190;
  assign N3959 = N3719 & idx_w_i[7];
  assign N3960 = N3721 & N1190;
  assign N3961 = N3721 & idx_w_i[7];
  assign N3962 = N3723 & N1190;
  assign N3963 = N3723 & idx_w_i[7];
  assign N3964 = N3725 & N1190;
  assign N3965 = N3725 & idx_w_i[7];
  assign N3966 = N3727 & N1190;
  assign N3967 = N3727 & idx_w_i[7];
  assign N3968 = N3729 & N1190;
  assign N3969 = N3729 & idx_w_i[7];
  assign N3970 = N3731 & N1190;
  assign N3971 = N3731 & idx_w_i[7];
  assign N3972 = N3733 & N1190;
  assign N3973 = N3733 & idx_w_i[7];
  assign N3974 = N3735 & N1190;
  assign N3975 = N3735 & idx_w_i[7];
  assign N3976 = N3737 & N1190;
  assign N3977 = N3737 & idx_w_i[7];
  assign N3978 = N3739 & N1190;
  assign N3979 = N3739 & idx_w_i[7];
  assign N3980 = N3741 & N1190;
  assign N3981 = N3741 & idx_w_i[7];
  assign N3982 = N3743 & N1190;
  assign N3983 = N3743 & idx_w_i[7];
  assign N3984 = N3745 & N1190;
  assign N3985 = N3745 & idx_w_i[7];
  assign N3986 = N3747 & N1190;
  assign N3987 = N3747 & idx_w_i[7];
  assign N3988 = N3749 & N1190;
  assign N3989 = N3749 & idx_w_i[7];
  assign N3990 = N3751 & N1190;
  assign N3991 = N3751 & idx_w_i[7];
  assign N3992 = N3753 & N1190;
  assign N3993 = N3753 & idx_w_i[7];
  assign N3994 = N3755 & N1190;
  assign N3995 = N3755 & idx_w_i[7];
  assign N3996 = N3757 & N1190;
  assign N3997 = N3757 & idx_w_i[7];
  assign N3998 = N3759 & N1190;
  assign N3999 = N3759 & idx_w_i[7];
  assign N4000 = N3761 & N1190;
  assign N4001 = N3761 & idx_w_i[7];
  assign N4002 = N3763 & N1190;
  assign N4003 = N3763 & idx_w_i[7];
  assign N4004 = N3765 & N1190;
  assign N4005 = N3765 & idx_w_i[7];
  assign N4006 = N3767 & N1190;
  assign N4007 = N3767 & idx_w_i[7];
  assign N4008 = N3769 & N1190;
  assign N4009 = N3769 & idx_w_i[7];
  assign N4010 = N3771 & N1190;
  assign N4011 = N3771 & idx_w_i[7];
  assign N4012 = N3773 & N1190;
  assign N4013 = N3773 & idx_w_i[7];
  assign N4014 = N3775 & N1190;
  assign N4015 = N3775 & idx_w_i[7];
  assign N4016 = N3777 & N1190;
  assign N4017 = N3777 & idx_w_i[7];
  assign N4018 = N3779 & N1190;
  assign N4019 = N3779 & idx_w_i[7];
  assign N4020 = N3781 & N1190;
  assign N4021 = N3781 & idx_w_i[7];
  assign N4022 = N3783 & N1190;
  assign N4023 = N3783 & idx_w_i[7];
  assign N4024 = N3785 & N1190;
  assign N4025 = N3785 & idx_w_i[7];
  assign N4026 = N3787 & N1190;
  assign N4027 = N3787 & idx_w_i[7];
  assign N4028 = N3789 & N1190;
  assign N4029 = N3789 & idx_w_i[7];
  assign N4030 = N3791 & N1190;
  assign N4031 = N3791 & idx_w_i[7];
  assign N4032 = N3793 & N1190;
  assign N4033 = N3793 & idx_w_i[7];
  assign N4034 = N3795 & N1190;
  assign N4035 = N3795 & idx_w_i[7];
  assign N4036 = N3797 & N1190;
  assign N4037 = N3797 & idx_w_i[7];
  assign N4038 = N3799 & N1190;
  assign N4039 = N3799 & idx_w_i[7];
  assign N4040 = N3801 & N1190;
  assign N4041 = N3801 & idx_w_i[7];
  assign N4042 = N3803 & N1190;
  assign N4043 = N3803 & idx_w_i[7];
  assign N4044 = N3805 & N1190;
  assign N4045 = N3805 & idx_w_i[7];
  assign N4046 = N3807 & N1190;
  assign N4047 = N3807 & idx_w_i[7];
  assign N4048 = N3809 & N1190;
  assign N4049 = N3809 & idx_w_i[7];
  assign N4050 = N3811 & N1190;
  assign N4051 = N3811 & idx_w_i[7];
  assign N4052 = N2876 & N1190;
  assign N4053 = N2878 & N1190;
  assign N4054 = N2880 & N1190;
  assign N4055 = N2882 & N1190;
  assign N4056 = N2884 & N1190;
  assign N4057 = N2886 & N1190;
  assign N4058 = N2888 & N1190;
  assign N4059 = N2890 & N1190;
  assign N4060 = N11329 & N1190;
  assign N4061 = N11331 & N1190;
  assign N4062 = N11333 & N1190;
  assign N4063 = N11335 & N1190;
  assign N4064 = N11337 & N1190;
  assign N4065 = N11339 & N1190;
  assign N4066 = N11341 & N1190;
  assign N4067 = N11343 & N1190;
  assign N4068 = N3828 & N1415;
  assign N4069 = N3828 & idx_w_i[8];
  assign N4070 = N3830 & N1415;
  assign N4071 = N3830 & idx_w_i[8];
  assign N4072 = N3832 & N1415;
  assign N4073 = N3832 & idx_w_i[8];
  assign N4074 = N3834 & N1415;
  assign N4075 = N3834 & idx_w_i[8];
  assign N4076 = N3836 & N1415;
  assign N4077 = N3836 & idx_w_i[8];
  assign N4078 = N3838 & N1415;
  assign N4079 = N3838 & idx_w_i[8];
  assign N4080 = N3840 & N1415;
  assign N4081 = N3840 & idx_w_i[8];
  assign N4082 = N3842 & N1415;
  assign N4083 = N3842 & idx_w_i[8];
  assign N4084 = N3844 & N1415;
  assign N4085 = N3844 & idx_w_i[8];
  assign N4086 = N3846 & N1415;
  assign N4087 = N3846 & idx_w_i[8];
  assign N4088 = N3848 & N1415;
  assign N4089 = N3848 & idx_w_i[8];
  assign N4090 = N3850 & N1415;
  assign N4091 = N3850 & idx_w_i[8];
  assign N4092 = N3852 & N1415;
  assign N4093 = N3852 & idx_w_i[8];
  assign N4094 = N3854 & N1415;
  assign N4095 = N3854 & idx_w_i[8];
  assign N4096 = N3856 & N1415;
  assign N4097 = N3856 & idx_w_i[8];
  assign N4098 = N3858 & N1415;
  assign N4099 = N3858 & idx_w_i[8];
  assign N4100 = N3860 & N1415;
  assign N4101 = N3860 & idx_w_i[8];
  assign N4102 = N3862 & N1415;
  assign N4103 = N3862 & idx_w_i[8];
  assign N4104 = N3864 & N1415;
  assign N4105 = N3864 & idx_w_i[8];
  assign N4106 = N3866 & N1415;
  assign N4107 = N3866 & idx_w_i[8];
  assign N4108 = N3868 & N1415;
  assign N4109 = N3868 & idx_w_i[8];
  assign N4110 = N3870 & N1415;
  assign N4111 = N3870 & idx_w_i[8];
  assign N4112 = N3872 & N1415;
  assign N4113 = N3872 & idx_w_i[8];
  assign N4114 = N3874 & N1415;
  assign N4115 = N3874 & idx_w_i[8];
  assign N4116 = N3876 & N1415;
  assign N4117 = N3876 & idx_w_i[8];
  assign N4118 = N3878 & N1415;
  assign N4119 = N3878 & idx_w_i[8];
  assign N4120 = N3880 & N1415;
  assign N4121 = N3880 & idx_w_i[8];
  assign N4122 = N3882 & N1415;
  assign N4123 = N3882 & idx_w_i[8];
  assign N4124 = N3884 & N1415;
  assign N4125 = N3884 & idx_w_i[8];
  assign N4126 = N3886 & N1415;
  assign N4127 = N3886 & idx_w_i[8];
  assign N4128 = N3888 & N1415;
  assign N4129 = N3888 & idx_w_i[8];
  assign N4130 = N3890 & N1415;
  assign N4131 = N3890 & idx_w_i[8];
  assign N4132 = N3892 & N1415;
  assign N4133 = N3892 & idx_w_i[8];
  assign N4134 = N3894 & N1415;
  assign N4135 = N3894 & idx_w_i[8];
  assign N4136 = N3896 & N1415;
  assign N4137 = N3896 & idx_w_i[8];
  assign N4138 = N3898 & N1415;
  assign N4139 = N3898 & idx_w_i[8];
  assign N4140 = N3900 & N1415;
  assign N4141 = N3900 & idx_w_i[8];
  assign N4142 = N3902 & N1415;
  assign N4143 = N3902 & idx_w_i[8];
  assign N4144 = N3904 & N1415;
  assign N4145 = N3904 & idx_w_i[8];
  assign N4146 = N3906 & N1415;
  assign N4147 = N3906 & idx_w_i[8];
  assign N4148 = N3908 & N1415;
  assign N4149 = N3908 & idx_w_i[8];
  assign N4150 = N3910 & N1415;
  assign N4151 = N3910 & idx_w_i[8];
  assign N4152 = N3912 & N1415;
  assign N4153 = N3912 & idx_w_i[8];
  assign N4154 = N3914 & N1415;
  assign N4155 = N3914 & idx_w_i[8];
  assign N4156 = N3916 & N1415;
  assign N4157 = N3916 & idx_w_i[8];
  assign N4158 = N3918 & N1415;
  assign N4159 = N3918 & idx_w_i[8];
  assign N4160 = N3920 & N1415;
  assign N4161 = N3920 & idx_w_i[8];
  assign N4162 = N3922 & N1415;
  assign N4163 = N3922 & idx_w_i[8];
  assign N4164 = N3924 & N1415;
  assign N4165 = N3924 & idx_w_i[8];
  assign N4166 = N3926 & N1415;
  assign N4167 = N3926 & idx_w_i[8];
  assign N4168 = N3928 & N1415;
  assign N4169 = N3928 & idx_w_i[8];
  assign N4170 = N3930 & N1415;
  assign N4171 = N3930 & idx_w_i[8];
  assign N4172 = N3932 & N1415;
  assign N4173 = N3932 & idx_w_i[8];
  assign N4174 = N3934 & N1415;
  assign N4175 = N3934 & idx_w_i[8];
  assign N4176 = N3936 & N1415;
  assign N4177 = N3936 & idx_w_i[8];
  assign N4178 = N3938 & N1415;
  assign N4179 = N3938 & idx_w_i[8];
  assign N4180 = N3940 & N1415;
  assign N4181 = N3940 & idx_w_i[8];
  assign N4182 = N3942 & N1415;
  assign N4183 = N3942 & idx_w_i[8];
  assign N4184 = N3944 & N1415;
  assign N4185 = N3944 & idx_w_i[8];
  assign N4186 = N3946 & N1415;
  assign N4187 = N3946 & idx_w_i[8];
  assign N4188 = N3948 & N1415;
  assign N4189 = N3948 & idx_w_i[8];
  assign N4190 = N3950 & N1415;
  assign N4191 = N3950 & idx_w_i[8];
  assign N4192 = N3952 & N1415;
  assign N4193 = N3952 & idx_w_i[8];
  assign N4194 = N3954 & N1415;
  assign N4195 = N3954 & idx_w_i[8];
  assign N4196 = N3956 & N1415;
  assign N4197 = N3956 & idx_w_i[8];
  assign N4198 = N3958 & N1415;
  assign N4199 = N3958 & idx_w_i[8];
  assign N4200 = N3960 & N1415;
  assign N4201 = N3960 & idx_w_i[8];
  assign N4202 = N3962 & N1415;
  assign N4203 = N3962 & idx_w_i[8];
  assign N4204 = N3964 & N1415;
  assign N4205 = N3964 & idx_w_i[8];
  assign N4206 = N3966 & N1415;
  assign N4207 = N3966 & idx_w_i[8];
  assign N4208 = N3968 & N1415;
  assign N4209 = N3968 & idx_w_i[8];
  assign N4210 = N3970 & N1415;
  assign N4211 = N3970 & idx_w_i[8];
  assign N4212 = N3972 & N1415;
  assign N4213 = N3972 & idx_w_i[8];
  assign N4214 = N3974 & N1415;
  assign N4215 = N3974 & idx_w_i[8];
  assign N4216 = N3976 & N1415;
  assign N4217 = N3976 & idx_w_i[8];
  assign N4218 = N3978 & N1415;
  assign N4219 = N3978 & idx_w_i[8];
  assign N4220 = N3980 & N1415;
  assign N4221 = N3980 & idx_w_i[8];
  assign N4222 = N3982 & N1415;
  assign N4223 = N3982 & idx_w_i[8];
  assign N4224 = N3984 & N1415;
  assign N4225 = N3984 & idx_w_i[8];
  assign N4226 = N3986 & N1415;
  assign N4227 = N3986 & idx_w_i[8];
  assign N4228 = N3988 & N1415;
  assign N4229 = N3988 & idx_w_i[8];
  assign N4230 = N3990 & N1415;
  assign N4231 = N3990 & idx_w_i[8];
  assign N4232 = N3992 & N1415;
  assign N4233 = N3992 & idx_w_i[8];
  assign N4234 = N3994 & N1415;
  assign N4235 = N3994 & idx_w_i[8];
  assign N4236 = N3996 & N1415;
  assign N4237 = N3996 & idx_w_i[8];
  assign N4238 = N3998 & N1415;
  assign N4239 = N3998 & idx_w_i[8];
  assign N4240 = N4000 & N1415;
  assign N4241 = N4000 & idx_w_i[8];
  assign N4242 = N4002 & N1415;
  assign N4243 = N4002 & idx_w_i[8];
  assign N4244 = N4004 & N1415;
  assign N4245 = N4004 & idx_w_i[8];
  assign N4246 = N4006 & N1415;
  assign N4247 = N4006 & idx_w_i[8];
  assign N4248 = N4008 & N1415;
  assign N4249 = N4008 & idx_w_i[8];
  assign N4250 = N4010 & N1415;
  assign N4251 = N4010 & idx_w_i[8];
  assign N4252 = N4012 & N1415;
  assign N4253 = N4012 & idx_w_i[8];
  assign N4254 = N4014 & N1415;
  assign N4255 = N4014 & idx_w_i[8];
  assign N4256 = N4016 & N1415;
  assign N4257 = N4016 & idx_w_i[8];
  assign N4258 = N4018 & N1415;
  assign N4259 = N4018 & idx_w_i[8];
  assign N4260 = N4020 & N1415;
  assign N4261 = N4020 & idx_w_i[8];
  assign N4262 = N4022 & N1415;
  assign N4263 = N4022 & idx_w_i[8];
  assign N4264 = N4024 & N1415;
  assign N4265 = N4024 & idx_w_i[8];
  assign N4266 = N4026 & N1415;
  assign N4267 = N4026 & idx_w_i[8];
  assign N4268 = N4028 & N1415;
  assign N4269 = N4028 & idx_w_i[8];
  assign N4270 = N4030 & N1415;
  assign N4271 = N4030 & idx_w_i[8];
  assign N4272 = N4032 & N1415;
  assign N4273 = N4032 & idx_w_i[8];
  assign N4274 = N4034 & N1415;
  assign N4275 = N4034 & idx_w_i[8];
  assign N4276 = N4036 & N1415;
  assign N4277 = N4036 & idx_w_i[8];
  assign N4278 = N4038 & N1415;
  assign N4279 = N4038 & idx_w_i[8];
  assign N4280 = N4040 & N1415;
  assign N4281 = N4040 & idx_w_i[8];
  assign N4282 = N4042 & N1415;
  assign N4283 = N4042 & idx_w_i[8];
  assign N4284 = N4044 & N1415;
  assign N4285 = N4044 & idx_w_i[8];
  assign N4286 = N4046 & N1415;
  assign N4287 = N4046 & idx_w_i[8];
  assign N4288 = N4048 & N1415;
  assign N4289 = N4048 & idx_w_i[8];
  assign N4290 = N4050 & N1415;
  assign N4291 = N4050 & idx_w_i[8];
  assign N4292 = N4052 & N1415;
  assign N4293 = N4052 & idx_w_i[8];
  assign N4294 = N4053 & N1415;
  assign N4295 = N4053 & idx_w_i[8];
  assign N4296 = N4054 & N1415;
  assign N4297 = N4054 & idx_w_i[8];
  assign N4298 = N4055 & N1415;
  assign N4299 = N4055 & idx_w_i[8];
  assign N4300 = N4056 & N1415;
  assign N4301 = N4056 & idx_w_i[8];
  assign N4302 = N4057 & N1415;
  assign N4303 = N4057 & idx_w_i[8];
  assign N4304 = N4058 & N1415;
  assign N4305 = N4058 & idx_w_i[8];
  assign N4306 = N4059 & N1415;
  assign N4307 = N4059 & idx_w_i[8];
  assign N4308 = N4060 & N1415;
  assign N4309 = N4060 & idx_w_i[8];
  assign N4310 = N4061 & N1415;
  assign N4311 = N4061 & idx_w_i[8];
  assign N4312 = N4062 & N1415;
  assign N4313 = N4062 & idx_w_i[8];
  assign N4314 = N4063 & N1415;
  assign N4315 = N4063 & idx_w_i[8];
  assign N4316 = N4064 & N1415;
  assign N4317 = N4064 & idx_w_i[8];
  assign N4318 = N4065 & N1415;
  assign N4319 = N4065 & idx_w_i[8];
  assign N4320 = N4066 & N1415;
  assign N4321 = N4066 & idx_w_i[8];
  assign N4322 = N4067 & N1415;
  assign N4323 = N4067 & idx_w_i[8];
  assign N4324 = N3829 & N1415;
  assign N4325 = N3829 & idx_w_i[8];
  assign N4326 = N3831 & N1415;
  assign N4327 = N3831 & idx_w_i[8];
  assign N4328 = N3833 & N1415;
  assign N4329 = N3833 & idx_w_i[8];
  assign N4330 = N3835 & N1415;
  assign N4331 = N3835 & idx_w_i[8];
  assign N4332 = N3837 & N1415;
  assign N4333 = N3837 & idx_w_i[8];
  assign N4334 = N3839 & N1415;
  assign N4335 = N3839 & idx_w_i[8];
  assign N4336 = N3841 & N1415;
  assign N4337 = N3841 & idx_w_i[8];
  assign N4338 = N3843 & N1415;
  assign N4339 = N3843 & idx_w_i[8];
  assign N4340 = N3845 & N1415;
  assign N4341 = N3845 & idx_w_i[8];
  assign N4342 = N3847 & N1415;
  assign N4343 = N3847 & idx_w_i[8];
  assign N4344 = N3849 & N1415;
  assign N4345 = N3849 & idx_w_i[8];
  assign N4346 = N3851 & N1415;
  assign N4347 = N3851 & idx_w_i[8];
  assign N4348 = N3853 & N1415;
  assign N4349 = N3853 & idx_w_i[8];
  assign N4350 = N3855 & N1415;
  assign N4351 = N3855 & idx_w_i[8];
  assign N4352 = N3857 & N1415;
  assign N4353 = N3857 & idx_w_i[8];
  assign N4354 = N3859 & N1415;
  assign N4355 = N3859 & idx_w_i[8];
  assign N4356 = N3861 & N1415;
  assign N4357 = N3861 & idx_w_i[8];
  assign N4358 = N3863 & N1415;
  assign N4359 = N3863 & idx_w_i[8];
  assign N4360 = N3865 & N1415;
  assign N4361 = N3865 & idx_w_i[8];
  assign N4362 = N3867 & N1415;
  assign N4363 = N3867 & idx_w_i[8];
  assign N4364 = N3869 & N1415;
  assign N4365 = N3869 & idx_w_i[8];
  assign N4366 = N3871 & N1415;
  assign N4367 = N3871 & idx_w_i[8];
  assign N4368 = N3873 & N1415;
  assign N4369 = N3873 & idx_w_i[8];
  assign N4370 = N3875 & N1415;
  assign N4371 = N3875 & idx_w_i[8];
  assign N4372 = N3877 & N1415;
  assign N4373 = N3877 & idx_w_i[8];
  assign N4374 = N3879 & N1415;
  assign N4375 = N3879 & idx_w_i[8];
  assign N4376 = N3881 & N1415;
  assign N4377 = N3881 & idx_w_i[8];
  assign N4378 = N3883 & N1415;
  assign N4379 = N3883 & idx_w_i[8];
  assign N4380 = N3885 & N1415;
  assign N4381 = N3885 & idx_w_i[8];
  assign N4382 = N3887 & N1415;
  assign N4383 = N3887 & idx_w_i[8];
  assign N4384 = N3889 & N1415;
  assign N4385 = N3889 & idx_w_i[8];
  assign N4386 = N3891 & N1415;
  assign N4387 = N3891 & idx_w_i[8];
  assign N4388 = N3893 & N1415;
  assign N4389 = N3893 & idx_w_i[8];
  assign N4390 = N3895 & N1415;
  assign N4391 = N3895 & idx_w_i[8];
  assign N4392 = N3897 & N1415;
  assign N4393 = N3897 & idx_w_i[8];
  assign N4394 = N3899 & N1415;
  assign N4395 = N3899 & idx_w_i[8];
  assign N4396 = N3901 & N1415;
  assign N4397 = N3901 & idx_w_i[8];
  assign N4398 = N3903 & N1415;
  assign N4399 = N3903 & idx_w_i[8];
  assign N4400 = N3905 & N1415;
  assign N4401 = N3905 & idx_w_i[8];
  assign N4402 = N3907 & N1415;
  assign N4403 = N3907 & idx_w_i[8];
  assign N4404 = N3909 & N1415;
  assign N4405 = N3909 & idx_w_i[8];
  assign N4406 = N3911 & N1415;
  assign N4407 = N3911 & idx_w_i[8];
  assign N4408 = N3913 & N1415;
  assign N4409 = N3913 & idx_w_i[8];
  assign N4410 = N3915 & N1415;
  assign N4411 = N3915 & idx_w_i[8];
  assign N4412 = N3917 & N1415;
  assign N4413 = N3917 & idx_w_i[8];
  assign N4414 = N3919 & N1415;
  assign N4415 = N3919 & idx_w_i[8];
  assign N4416 = N3921 & N1415;
  assign N4417 = N3921 & idx_w_i[8];
  assign N4418 = N3923 & N1415;
  assign N4419 = N3923 & idx_w_i[8];
  assign N4420 = N3925 & N1415;
  assign N4421 = N3925 & idx_w_i[8];
  assign N4422 = N3927 & N1415;
  assign N4423 = N3927 & idx_w_i[8];
  assign N4424 = N3929 & N1415;
  assign N4425 = N3929 & idx_w_i[8];
  assign N4426 = N3931 & N1415;
  assign N4427 = N3931 & idx_w_i[8];
  assign N4428 = N3933 & N1415;
  assign N4429 = N3933 & idx_w_i[8];
  assign N4430 = N3935 & N1415;
  assign N4431 = N3935 & idx_w_i[8];
  assign N4432 = N3937 & N1415;
  assign N4433 = N3937 & idx_w_i[8];
  assign N4434 = N3939 & N1415;
  assign N4435 = N3939 & idx_w_i[8];
  assign N4436 = N3941 & N1415;
  assign N4437 = N3941 & idx_w_i[8];
  assign N4438 = N3943 & N1415;
  assign N4439 = N3943 & idx_w_i[8];
  assign N4440 = N3945 & N1415;
  assign N4441 = N3945 & idx_w_i[8];
  assign N4442 = N3947 & N1415;
  assign N4443 = N3947 & idx_w_i[8];
  assign N4444 = N3949 & N1415;
  assign N4445 = N3949 & idx_w_i[8];
  assign N4446 = N3951 & N1415;
  assign N4447 = N3951 & idx_w_i[8];
  assign N4448 = N3953 & N1415;
  assign N4449 = N3953 & idx_w_i[8];
  assign N4450 = N3955 & N1415;
  assign N4451 = N3955 & idx_w_i[8];
  assign N4452 = N3957 & N1415;
  assign N4453 = N3957 & idx_w_i[8];
  assign N4454 = N3959 & N1415;
  assign N4455 = N3959 & idx_w_i[8];
  assign N4456 = N3961 & N1415;
  assign N4457 = N3961 & idx_w_i[8];
  assign N4458 = N3963 & N1415;
  assign N4459 = N3963 & idx_w_i[8];
  assign N4460 = N3965 & N1415;
  assign N4461 = N3965 & idx_w_i[8];
  assign N4462 = N3967 & N1415;
  assign N4463 = N3967 & idx_w_i[8];
  assign N4464 = N3969 & N1415;
  assign N4465 = N3969 & idx_w_i[8];
  assign N4466 = N3971 & N1415;
  assign N4467 = N3971 & idx_w_i[8];
  assign N4468 = N3973 & N1415;
  assign N4469 = N3973 & idx_w_i[8];
  assign N4470 = N3975 & N1415;
  assign N4471 = N3975 & idx_w_i[8];
  assign N4472 = N3977 & N1415;
  assign N4473 = N3977 & idx_w_i[8];
  assign N4474 = N3979 & N1415;
  assign N4475 = N3979 & idx_w_i[8];
  assign N4476 = N3981 & N1415;
  assign N4477 = N3981 & idx_w_i[8];
  assign N4478 = N3983 & N1415;
  assign N4479 = N3983 & idx_w_i[8];
  assign N4480 = N3985 & N1415;
  assign N4481 = N3985 & idx_w_i[8];
  assign N4482 = N3987 & N1415;
  assign N4483 = N3987 & idx_w_i[8];
  assign N4484 = N3989 & N1415;
  assign N4485 = N3989 & idx_w_i[8];
  assign N4486 = N3991 & N1415;
  assign N4487 = N3991 & idx_w_i[8];
  assign N4488 = N3993 & N1415;
  assign N4489 = N3993 & idx_w_i[8];
  assign N4490 = N3995 & N1415;
  assign N4491 = N3995 & idx_w_i[8];
  assign N4492 = N3997 & N1415;
  assign N4493 = N3997 & idx_w_i[8];
  assign N4494 = N3999 & N1415;
  assign N4495 = N3999 & idx_w_i[8];
  assign N4496 = N4001 & N1415;
  assign N4497 = N4001 & idx_w_i[8];
  assign N4498 = N4003 & N1415;
  assign N4499 = N4003 & idx_w_i[8];
  assign N4500 = N4005 & N1415;
  assign N4501 = N4005 & idx_w_i[8];
  assign N4502 = N4007 & N1415;
  assign N4503 = N4007 & idx_w_i[8];
  assign N4504 = N4009 & N1415;
  assign N4505 = N4009 & idx_w_i[8];
  assign N4506 = N4011 & N1415;
  assign N4507 = N4011 & idx_w_i[8];
  assign N4508 = N4013 & N1415;
  assign N4509 = N4013 & idx_w_i[8];
  assign N4510 = N4015 & N1415;
  assign N4511 = N4015 & idx_w_i[8];
  assign N4512 = N4017 & N1415;
  assign N4513 = N4017 & idx_w_i[8];
  assign N4514 = N4019 & N1415;
  assign N4515 = N4019 & idx_w_i[8];
  assign N4516 = N4021 & N1415;
  assign N4517 = N4021 & idx_w_i[8];
  assign N4518 = N4023 & N1415;
  assign N4519 = N4023 & idx_w_i[8];
  assign N4520 = N4025 & N1415;
  assign N4521 = N4025 & idx_w_i[8];
  assign N4522 = N4027 & N1415;
  assign N4523 = N4027 & idx_w_i[8];
  assign N4524 = N4029 & N1415;
  assign N4525 = N4029 & idx_w_i[8];
  assign N4526 = N4031 & N1415;
  assign N4527 = N4031 & idx_w_i[8];
  assign N4528 = N4033 & N1415;
  assign N4529 = N4033 & idx_w_i[8];
  assign N4530 = N4035 & N1415;
  assign N4531 = N4035 & idx_w_i[8];
  assign N4532 = N4037 & N1415;
  assign N4533 = N4037 & idx_w_i[8];
  assign N4534 = N4039 & N1415;
  assign N4535 = N4039 & idx_w_i[8];
  assign N4536 = N4041 & N1415;
  assign N4537 = N4041 & idx_w_i[8];
  assign N4538 = N4043 & N1415;
  assign N4539 = N4043 & idx_w_i[8];
  assign N4540 = N4045 & N1415;
  assign N4541 = N4045 & idx_w_i[8];
  assign N4542 = N4047 & N1415;
  assign N4543 = N4047 & idx_w_i[8];
  assign N4544 = N4049 & N1415;
  assign N4545 = N4049 & idx_w_i[8];
  assign N4546 = N4051 & N1415;
  assign N4547 = N4051 & idx_w_i[8];
  assign N4548 = N3124 & N1415;
  assign N4549 = N3126 & N1415;
  assign N4550 = N3128 & N1415;
  assign N4551 = N3130 & N1415;
  assign N4552 = N3132 & N1415;
  assign N4553 = N3134 & N1415;
  assign N4554 = N3136 & N1415;
  assign N4555 = N3138 & N1415;
  assign N4556 = N11585 & N1415;
  assign N4557 = N11587 & N1415;
  assign N4558 = N11589 & N1415;
  assign N4559 = N11591 & N1415;
  assign N4560 = N11593 & N1415;
  assign N4561 = N11595 & N1415;
  assign N4562 = N11597 & N1415;
  assign N4563 = N11599 & N1415;
  assign N5077 = N3651 ^ N4564;
  assign N5078 = N11104 & N2698;
  assign N5079 = N11106 & N2698;
  assign N5080 = N11108 & N2698;
  assign N5081 = N11110 & N2698;
  assign N5082 = N11112 & N2698;
  assign N5083 = N11114 & N2698;
  assign N5084 = N11116 & N2698;
  assign N5085 = N11118 & N2698;
  assign N5086 = N5078 & N1060;
  assign N5087 = N5078 & idx_w_i[5];
  assign N5088 = N5079 & N1060;
  assign N5089 = N5079 & idx_w_i[5];
  assign N5090 = N5080 & N1060;
  assign N5091 = N5080 & idx_w_i[5];
  assign N5092 = N5081 & N1060;
  assign N5093 = N5081 & idx_w_i[5];
  assign N5094 = N5082 & N1060;
  assign N5095 = N5082 & idx_w_i[5];
  assign N5096 = N5083 & N1060;
  assign N5097 = N5083 & idx_w_i[5];
  assign N5098 = N5084 & N1060;
  assign N5099 = N5084 & idx_w_i[5];
  assign N5100 = N5085 & N1060;
  assign N5101 = N5085 & idx_w_i[5];
  assign N5102 = N3660 & N1060;
  assign N5103 = N3661 & N1060;
  assign N5104 = N3662 & N1060;
  assign N5105 = N3663 & N1060;
  assign N5106 = N3664 & N1060;
  assign N5107 = N3665 & N1060;
  assign N5108 = N3666 & N1060;
  assign N5109 = N3667 & N1060;
  assign N5110 = N11121 & N1060;
  assign N5111 = N11123 & N1060;
  assign N5112 = N11125 & N1060;
  assign N5113 = N11127 & N1060;
  assign N5114 = N11129 & N1060;
  assign N5115 = N11131 & N1060;
  assign N5116 = N11133 & N1060;
  assign N5117 = N11135 & N1060;
  assign N5118 = N11137 & N1060;
  assign N5119 = N11139 & N1060;
  assign N5120 = N11141 & N1060;
  assign N5121 = N11143 & N1060;
  assign N5122 = N11145 & N1060;
  assign N5123 = N11147 & N1060;
  assign N5124 = N11149 & N1060;
  assign N5125 = N11151 & N1060;
  assign N5126 = N5086 & N1093;
  assign N5127 = N5086 & idx_w_i[6];
  assign N5128 = N5088 & N1093;
  assign N5129 = N5088 & idx_w_i[6];
  assign N5130 = N5090 & N1093;
  assign N5131 = N5090 & idx_w_i[6];
  assign N5132 = N5092 & N1093;
  assign N5133 = N5092 & idx_w_i[6];
  assign N5134 = N5094 & N1093;
  assign N5135 = N5094 & idx_w_i[6];
  assign N5136 = N5096 & N1093;
  assign N5137 = N5096 & idx_w_i[6];
  assign N5138 = N5098 & N1093;
  assign N5139 = N5098 & idx_w_i[6];
  assign N5140 = N5100 & N1093;
  assign N5141 = N5100 & idx_w_i[6];
  assign N5142 = N5102 & N1093;
  assign N5143 = N5102 & idx_w_i[6];
  assign N5144 = N5103 & N1093;
  assign N5145 = N5103 & idx_w_i[6];
  assign N5146 = N5104 & N1093;
  assign N5147 = N5104 & idx_w_i[6];
  assign N5148 = N5105 & N1093;
  assign N5149 = N5105 & idx_w_i[6];
  assign N5150 = N5106 & N1093;
  assign N5151 = N5106 & idx_w_i[6];
  assign N5152 = N5107 & N1093;
  assign N5153 = N5107 & idx_w_i[6];
  assign N5154 = N5108 & N1093;
  assign N5155 = N5108 & idx_w_i[6];
  assign N5156 = N5109 & N1093;
  assign N5157 = N5109 & idx_w_i[6];
  assign N5158 = N5110 & N1093;
  assign N5159 = N5110 & idx_w_i[6];
  assign N5160 = N5111 & N1093;
  assign N5161 = N5111 & idx_w_i[6];
  assign N5162 = N5112 & N1093;
  assign N5163 = N5112 & idx_w_i[6];
  assign N5164 = N5113 & N1093;
  assign N5165 = N5113 & idx_w_i[6];
  assign N5166 = N5114 & N1093;
  assign N5167 = N5114 & idx_w_i[6];
  assign N5168 = N5115 & N1093;
  assign N5169 = N5115 & idx_w_i[6];
  assign N5170 = N5116 & N1093;
  assign N5171 = N5116 & idx_w_i[6];
  assign N5172 = N5117 & N1093;
  assign N5173 = N5117 & idx_w_i[6];
  assign N5174 = N5118 & N1093;
  assign N5175 = N5118 & idx_w_i[6];
  assign N5176 = N5119 & N1093;
  assign N5177 = N5119 & idx_w_i[6];
  assign N5178 = N5120 & N1093;
  assign N5179 = N5120 & idx_w_i[6];
  assign N5180 = N5121 & N1093;
  assign N5181 = N5121 & idx_w_i[6];
  assign N5182 = N5122 & N1093;
  assign N5183 = N5122 & idx_w_i[6];
  assign N5184 = N5123 & N1093;
  assign N5185 = N5123 & idx_w_i[6];
  assign N5186 = N5124 & N1093;
  assign N5187 = N5124 & idx_w_i[6];
  assign N5188 = N5125 & N1093;
  assign N5189 = N5125 & idx_w_i[6];
  assign N5190 = N5087 & N1093;
  assign N5191 = N5087 & idx_w_i[6];
  assign N5192 = N5089 & N1093;
  assign N5193 = N5089 & idx_w_i[6];
  assign N5194 = N5091 & N1093;
  assign N5195 = N5091 & idx_w_i[6];
  assign N5196 = N5093 & N1093;
  assign N5197 = N5093 & idx_w_i[6];
  assign N5198 = N5095 & N1093;
  assign N5199 = N5095 & idx_w_i[6];
  assign N5200 = N5097 & N1093;
  assign N5201 = N5097 & idx_w_i[6];
  assign N5202 = N5099 & N1093;
  assign N5203 = N5099 & idx_w_i[6];
  assign N5204 = N5101 & N1093;
  assign N5205 = N5101 & idx_w_i[6];
  assign N5206 = N3685 & N1093;
  assign N5207 = N3687 & N1093;
  assign N5208 = N3689 & N1093;
  assign N5209 = N3691 & N1093;
  assign N5210 = N3693 & N1093;
  assign N5211 = N3695 & N1093;
  assign N5212 = N3697 & N1093;
  assign N5213 = N3699 & N1093;
  assign N5214 = N11185 & N1093;
  assign N5215 = N11187 & N1093;
  assign N5216 = N11189 & N1093;
  assign N5217 = N11191 & N1093;
  assign N5218 = N11193 & N1093;
  assign N5219 = N11195 & N1093;
  assign N5220 = N11197 & N1093;
  assign N5221 = N11199 & N1093;
  assign N5222 = N11201 & N1093;
  assign N5223 = N11203 & N1093;
  assign N5224 = N11205 & N1093;
  assign N5225 = N11207 & N1093;
  assign N5226 = N11209 & N1093;
  assign N5227 = N11211 & N1093;
  assign N5228 = N11213 & N1093;
  assign N5229 = N11215 & N1093;
  assign N5230 = N5126 & N1190;
  assign N5231 = N5126 & idx_w_i[7];
  assign N5232 = N5128 & N1190;
  assign N5233 = N5128 & idx_w_i[7];
  assign N5234 = N5130 & N1190;
  assign N5235 = N5130 & idx_w_i[7];
  assign N5236 = N5132 & N1190;
  assign N5237 = N5132 & idx_w_i[7];
  assign N5238 = N5134 & N1190;
  assign N5239 = N5134 & idx_w_i[7];
  assign N5240 = N5136 & N1190;
  assign N5241 = N5136 & idx_w_i[7];
  assign N5242 = N5138 & N1190;
  assign N5243 = N5138 & idx_w_i[7];
  assign N5244 = N5140 & N1190;
  assign N5245 = N5140 & idx_w_i[7];
  assign N5246 = N5142 & N1190;
  assign N5247 = N5142 & idx_w_i[7];
  assign N5248 = N5144 & N1190;
  assign N5249 = N5144 & idx_w_i[7];
  assign N5250 = N5146 & N1190;
  assign N5251 = N5146 & idx_w_i[7];
  assign N5252 = N5148 & N1190;
  assign N5253 = N5148 & idx_w_i[7];
  assign N5254 = N5150 & N1190;
  assign N5255 = N5150 & idx_w_i[7];
  assign N5256 = N5152 & N1190;
  assign N5257 = N5152 & idx_w_i[7];
  assign N5258 = N5154 & N1190;
  assign N5259 = N5154 & idx_w_i[7];
  assign N5260 = N5156 & N1190;
  assign N5261 = N5156 & idx_w_i[7];
  assign N5262 = N5158 & N1190;
  assign N5263 = N5158 & idx_w_i[7];
  assign N5264 = N5160 & N1190;
  assign N5265 = N5160 & idx_w_i[7];
  assign N5266 = N5162 & N1190;
  assign N5267 = N5162 & idx_w_i[7];
  assign N5268 = N5164 & N1190;
  assign N5269 = N5164 & idx_w_i[7];
  assign N5270 = N5166 & N1190;
  assign N5271 = N5166 & idx_w_i[7];
  assign N5272 = N5168 & N1190;
  assign N5273 = N5168 & idx_w_i[7];
  assign N5274 = N5170 & N1190;
  assign N5275 = N5170 & idx_w_i[7];
  assign N5276 = N5172 & N1190;
  assign N5277 = N5172 & idx_w_i[7];
  assign N5278 = N5174 & N1190;
  assign N5279 = N5174 & idx_w_i[7];
  assign N5280 = N5176 & N1190;
  assign N5281 = N5176 & idx_w_i[7];
  assign N5282 = N5178 & N1190;
  assign N5283 = N5178 & idx_w_i[7];
  assign N5284 = N5180 & N1190;
  assign N5285 = N5180 & idx_w_i[7];
  assign N5286 = N5182 & N1190;
  assign N5287 = N5182 & idx_w_i[7];
  assign N5288 = N5184 & N1190;
  assign N5289 = N5184 & idx_w_i[7];
  assign N5290 = N5186 & N1190;
  assign N5291 = N5186 & idx_w_i[7];
  assign N5292 = N5188 & N1190;
  assign N5293 = N5188 & idx_w_i[7];
  assign N5294 = N5190 & N1190;
  assign N5295 = N5190 & idx_w_i[7];
  assign N5296 = N5192 & N1190;
  assign N5297 = N5192 & idx_w_i[7];
  assign N5298 = N5194 & N1190;
  assign N5299 = N5194 & idx_w_i[7];
  assign N5300 = N5196 & N1190;
  assign N5301 = N5196 & idx_w_i[7];
  assign N5302 = N5198 & N1190;
  assign N5303 = N5198 & idx_w_i[7];
  assign N5304 = N5200 & N1190;
  assign N5305 = N5200 & idx_w_i[7];
  assign N5306 = N5202 & N1190;
  assign N5307 = N5202 & idx_w_i[7];
  assign N5308 = N5204 & N1190;
  assign N5309 = N5204 & idx_w_i[7];
  assign N5310 = N5206 & N1190;
  assign N5311 = N5206 & idx_w_i[7];
  assign N5312 = N5207 & N1190;
  assign N5313 = N5207 & idx_w_i[7];
  assign N5314 = N5208 & N1190;
  assign N5315 = N5208 & idx_w_i[7];
  assign N5316 = N5209 & N1190;
  assign N5317 = N5209 & idx_w_i[7];
  assign N5318 = N5210 & N1190;
  assign N5319 = N5210 & idx_w_i[7];
  assign N5320 = N5211 & N1190;
  assign N5321 = N5211 & idx_w_i[7];
  assign N5322 = N5212 & N1190;
  assign N5323 = N5212 & idx_w_i[7];
  assign N5324 = N5213 & N1190;
  assign N5325 = N5213 & idx_w_i[7];
  assign N5326 = N5214 & N1190;
  assign N5327 = N5214 & idx_w_i[7];
  assign N5328 = N5215 & N1190;
  assign N5329 = N5215 & idx_w_i[7];
  assign N5330 = N5216 & N1190;
  assign N5331 = N5216 & idx_w_i[7];
  assign N5332 = N5217 & N1190;
  assign N5333 = N5217 & idx_w_i[7];
  assign N5334 = N5218 & N1190;
  assign N5335 = N5218 & idx_w_i[7];
  assign N5336 = N5219 & N1190;
  assign N5337 = N5219 & idx_w_i[7];
  assign N5338 = N5220 & N1190;
  assign N5339 = N5220 & idx_w_i[7];
  assign N5340 = N5221 & N1190;
  assign N5341 = N5221 & idx_w_i[7];
  assign N5342 = N5222 & N1190;
  assign N5343 = N5222 & idx_w_i[7];
  assign N5344 = N5223 & N1190;
  assign N5345 = N5223 & idx_w_i[7];
  assign N5346 = N5224 & N1190;
  assign N5347 = N5224 & idx_w_i[7];
  assign N5348 = N5225 & N1190;
  assign N5349 = N5225 & idx_w_i[7];
  assign N5350 = N5226 & N1190;
  assign N5351 = N5226 & idx_w_i[7];
  assign N5352 = N5227 & N1190;
  assign N5353 = N5227 & idx_w_i[7];
  assign N5354 = N5228 & N1190;
  assign N5355 = N5228 & idx_w_i[7];
  assign N5356 = N5229 & N1190;
  assign N5357 = N5229 & idx_w_i[7];
  assign N5358 = N5127 & N1190;
  assign N5359 = N5127 & idx_w_i[7];
  assign N5360 = N5129 & N1190;
  assign N5361 = N5129 & idx_w_i[7];
  assign N5362 = N5131 & N1190;
  assign N5363 = N5131 & idx_w_i[7];
  assign N5364 = N5133 & N1190;
  assign N5365 = N5133 & idx_w_i[7];
  assign N5366 = N5135 & N1190;
  assign N5367 = N5135 & idx_w_i[7];
  assign N5368 = N5137 & N1190;
  assign N5369 = N5137 & idx_w_i[7];
  assign N5370 = N5139 & N1190;
  assign N5371 = N5139 & idx_w_i[7];
  assign N5372 = N5141 & N1190;
  assign N5373 = N5141 & idx_w_i[7];
  assign N5374 = N5143 & N1190;
  assign N5375 = N5143 & idx_w_i[7];
  assign N5376 = N5145 & N1190;
  assign N5377 = N5145 & idx_w_i[7];
  assign N5378 = N5147 & N1190;
  assign N5379 = N5147 & idx_w_i[7];
  assign N5380 = N5149 & N1190;
  assign N5381 = N5149 & idx_w_i[7];
  assign N5382 = N5151 & N1190;
  assign N5383 = N5151 & idx_w_i[7];
  assign N5384 = N5153 & N1190;
  assign N5385 = N5153 & idx_w_i[7];
  assign N5386 = N5155 & N1190;
  assign N5387 = N5155 & idx_w_i[7];
  assign N5388 = N5157 & N1190;
  assign N5389 = N5157 & idx_w_i[7];
  assign N5390 = N5159 & N1190;
  assign N5391 = N5159 & idx_w_i[7];
  assign N5392 = N5161 & N1190;
  assign N5393 = N5161 & idx_w_i[7];
  assign N5394 = N5163 & N1190;
  assign N5395 = N5163 & idx_w_i[7];
  assign N5396 = N5165 & N1190;
  assign N5397 = N5165 & idx_w_i[7];
  assign N5398 = N5167 & N1190;
  assign N5399 = N5167 & idx_w_i[7];
  assign N5400 = N5169 & N1190;
  assign N5401 = N5169 & idx_w_i[7];
  assign N5402 = N5171 & N1190;
  assign N5403 = N5171 & idx_w_i[7];
  assign N5404 = N5173 & N1190;
  assign N5405 = N5173 & idx_w_i[7];
  assign N5406 = N5175 & N1190;
  assign N5407 = N5175 & idx_w_i[7];
  assign N5408 = N5177 & N1190;
  assign N5409 = N5177 & idx_w_i[7];
  assign N5410 = N5179 & N1190;
  assign N5411 = N5179 & idx_w_i[7];
  assign N5412 = N5181 & N1190;
  assign N5413 = N5181 & idx_w_i[7];
  assign N5414 = N5183 & N1190;
  assign N5415 = N5183 & idx_w_i[7];
  assign N5416 = N5185 & N1190;
  assign N5417 = N5185 & idx_w_i[7];
  assign N5418 = N5187 & N1190;
  assign N5419 = N5187 & idx_w_i[7];
  assign N5420 = N5189 & N1190;
  assign N5421 = N5189 & idx_w_i[7];
  assign N5422 = N5191 & N1190;
  assign N5423 = N5191 & idx_w_i[7];
  assign N5424 = N5193 & N1190;
  assign N5425 = N5193 & idx_w_i[7];
  assign N5426 = N5195 & N1190;
  assign N5427 = N5195 & idx_w_i[7];
  assign N5428 = N5197 & N1190;
  assign N5429 = N5197 & idx_w_i[7];
  assign N5430 = N5199 & N1190;
  assign N5431 = N5199 & idx_w_i[7];
  assign N5432 = N5201 & N1190;
  assign N5433 = N5201 & idx_w_i[7];
  assign N5434 = N5203 & N1190;
  assign N5435 = N5203 & idx_w_i[7];
  assign N5436 = N5205 & N1190;
  assign N5437 = N5205 & idx_w_i[7];
  assign N5438 = N3797 & N1190;
  assign N5439 = N3799 & N1190;
  assign N5440 = N3801 & N1190;
  assign N5441 = N3803 & N1190;
  assign N5442 = N3805 & N1190;
  assign N5443 = N3807 & N1190;
  assign N5444 = N3809 & N1190;
  assign N5445 = N3811 & N1190;
  assign N5446 = N11313 & N1190;
  assign N5447 = N11315 & N1190;
  assign N5448 = N11317 & N1190;
  assign N5449 = N11319 & N1190;
  assign N5450 = N11321 & N1190;
  assign N5451 = N11323 & N1190;
  assign N5452 = N11325 & N1190;
  assign N5453 = N11327 & N1190;
  assign N5454 = N11329 & N1190;
  assign N5455 = N11331 & N1190;
  assign N5456 = N11333 & N1190;
  assign N5457 = N11335 & N1190;
  assign N5458 = N11337 & N1190;
  assign N5459 = N11339 & N1190;
  assign N5460 = N11341 & N1190;
  assign N5461 = N11343 & N1190;
  assign N5462 = N5230 & N1415;
  assign N5463 = N5230 & idx_w_i[8];
  assign N5464 = N5232 & N1415;
  assign N5465 = N5232 & idx_w_i[8];
  assign N5466 = N5234 & N1415;
  assign N5467 = N5234 & idx_w_i[8];
  assign N5468 = N5236 & N1415;
  assign N5469 = N5236 & idx_w_i[8];
  assign N5470 = N5238 & N1415;
  assign N5471 = N5238 & idx_w_i[8];
  assign N5472 = N5240 & N1415;
  assign N5473 = N5240 & idx_w_i[8];
  assign N5474 = N5242 & N1415;
  assign N5475 = N5242 & idx_w_i[8];
  assign N5476 = N5244 & N1415;
  assign N5477 = N5244 & idx_w_i[8];
  assign N5478 = N5246 & N1415;
  assign N5479 = N5246 & idx_w_i[8];
  assign N5480 = N5248 & N1415;
  assign N5481 = N5248 & idx_w_i[8];
  assign N5482 = N5250 & N1415;
  assign N5483 = N5250 & idx_w_i[8];
  assign N5484 = N5252 & N1415;
  assign N5485 = N5252 & idx_w_i[8];
  assign N5486 = N5254 & N1415;
  assign N5487 = N5254 & idx_w_i[8];
  assign N5488 = N5256 & N1415;
  assign N5489 = N5256 & idx_w_i[8];
  assign N5490 = N5258 & N1415;
  assign N5491 = N5258 & idx_w_i[8];
  assign N5492 = N5260 & N1415;
  assign N5493 = N5260 & idx_w_i[8];
  assign N5494 = N5262 & N1415;
  assign N5495 = N5262 & idx_w_i[8];
  assign N5496 = N5264 & N1415;
  assign N5497 = N5264 & idx_w_i[8];
  assign N5498 = N5266 & N1415;
  assign N5499 = N5266 & idx_w_i[8];
  assign N5500 = N5268 & N1415;
  assign N5501 = N5268 & idx_w_i[8];
  assign N5502 = N5270 & N1415;
  assign N5503 = N5270 & idx_w_i[8];
  assign N5504 = N5272 & N1415;
  assign N5505 = N5272 & idx_w_i[8];
  assign N5506 = N5274 & N1415;
  assign N5507 = N5274 & idx_w_i[8];
  assign N5508 = N5276 & N1415;
  assign N5509 = N5276 & idx_w_i[8];
  assign N5510 = N5278 & N1415;
  assign N5511 = N5278 & idx_w_i[8];
  assign N5512 = N5280 & N1415;
  assign N5513 = N5280 & idx_w_i[8];
  assign N5514 = N5282 & N1415;
  assign N5515 = N5282 & idx_w_i[8];
  assign N5516 = N5284 & N1415;
  assign N5517 = N5284 & idx_w_i[8];
  assign N5518 = N5286 & N1415;
  assign N5519 = N5286 & idx_w_i[8];
  assign N5520 = N5288 & N1415;
  assign N5521 = N5288 & idx_w_i[8];
  assign N5522 = N5290 & N1415;
  assign N5523 = N5290 & idx_w_i[8];
  assign N5524 = N5292 & N1415;
  assign N5525 = N5292 & idx_w_i[8];
  assign N5526 = N5294 & N1415;
  assign N5527 = N5294 & idx_w_i[8];
  assign N5528 = N5296 & N1415;
  assign N5529 = N5296 & idx_w_i[8];
  assign N5530 = N5298 & N1415;
  assign N5531 = N5298 & idx_w_i[8];
  assign N5532 = N5300 & N1415;
  assign N5533 = N5300 & idx_w_i[8];
  assign N5534 = N5302 & N1415;
  assign N5535 = N5302 & idx_w_i[8];
  assign N5536 = N5304 & N1415;
  assign N5537 = N5304 & idx_w_i[8];
  assign N5538 = N5306 & N1415;
  assign N5539 = N5306 & idx_w_i[8];
  assign N5540 = N5308 & N1415;
  assign N5541 = N5308 & idx_w_i[8];
  assign N5542 = N5310 & N1415;
  assign N5543 = N5310 & idx_w_i[8];
  assign N5544 = N5312 & N1415;
  assign N5545 = N5312 & idx_w_i[8];
  assign N5546 = N5314 & N1415;
  assign N5547 = N5314 & idx_w_i[8];
  assign N5548 = N5316 & N1415;
  assign N5549 = N5316 & idx_w_i[8];
  assign N5550 = N5318 & N1415;
  assign N5551 = N5318 & idx_w_i[8];
  assign N5552 = N5320 & N1415;
  assign N5553 = N5320 & idx_w_i[8];
  assign N5554 = N5322 & N1415;
  assign N5555 = N5322 & idx_w_i[8];
  assign N5556 = N5324 & N1415;
  assign N5557 = N5324 & idx_w_i[8];
  assign N5558 = N5326 & N1415;
  assign N5559 = N5326 & idx_w_i[8];
  assign N5560 = N5328 & N1415;
  assign N5561 = N5328 & idx_w_i[8];
  assign N5562 = N5330 & N1415;
  assign N5563 = N5330 & idx_w_i[8];
  assign N5564 = N5332 & N1415;
  assign N5565 = N5332 & idx_w_i[8];
  assign N5566 = N5334 & N1415;
  assign N5567 = N5334 & idx_w_i[8];
  assign N5568 = N5336 & N1415;
  assign N5569 = N5336 & idx_w_i[8];
  assign N5570 = N5338 & N1415;
  assign N5571 = N5338 & idx_w_i[8];
  assign N5572 = N5340 & N1415;
  assign N5573 = N5340 & idx_w_i[8];
  assign N5574 = N5342 & N1415;
  assign N5575 = N5342 & idx_w_i[8];
  assign N5576 = N5344 & N1415;
  assign N5577 = N5344 & idx_w_i[8];
  assign N5578 = N5346 & N1415;
  assign N5579 = N5346 & idx_w_i[8];
  assign N5580 = N5348 & N1415;
  assign N5581 = N5348 & idx_w_i[8];
  assign N5582 = N5350 & N1415;
  assign N5583 = N5350 & idx_w_i[8];
  assign N5584 = N5352 & N1415;
  assign N5585 = N5352 & idx_w_i[8];
  assign N5586 = N5354 & N1415;
  assign N5587 = N5354 & idx_w_i[8];
  assign N5588 = N5356 & N1415;
  assign N5589 = N5356 & idx_w_i[8];
  assign N5590 = N5358 & N1415;
  assign N5591 = N5358 & idx_w_i[8];
  assign N5592 = N5360 & N1415;
  assign N5593 = N5360 & idx_w_i[8];
  assign N5594 = N5362 & N1415;
  assign N5595 = N5362 & idx_w_i[8];
  assign N5596 = N5364 & N1415;
  assign N5597 = N5364 & idx_w_i[8];
  assign N5598 = N5366 & N1415;
  assign N5599 = N5366 & idx_w_i[8];
  assign N5600 = N5368 & N1415;
  assign N5601 = N5368 & idx_w_i[8];
  assign N5602 = N5370 & N1415;
  assign N5603 = N5370 & idx_w_i[8];
  assign N5604 = N5372 & N1415;
  assign N5605 = N5372 & idx_w_i[8];
  assign N5606 = N5374 & N1415;
  assign N5607 = N5374 & idx_w_i[8];
  assign N5608 = N5376 & N1415;
  assign N5609 = N5376 & idx_w_i[8];
  assign N5610 = N5378 & N1415;
  assign N5611 = N5378 & idx_w_i[8];
  assign N5612 = N5380 & N1415;
  assign N5613 = N5380 & idx_w_i[8];
  assign N5614 = N5382 & N1415;
  assign N5615 = N5382 & idx_w_i[8];
  assign N5616 = N5384 & N1415;
  assign N5617 = N5384 & idx_w_i[8];
  assign N5618 = N5386 & N1415;
  assign N5619 = N5386 & idx_w_i[8];
  assign N5620 = N5388 & N1415;
  assign N5621 = N5388 & idx_w_i[8];
  assign N5622 = N5390 & N1415;
  assign N5623 = N5390 & idx_w_i[8];
  assign N5624 = N5392 & N1415;
  assign N5625 = N5392 & idx_w_i[8];
  assign N5626 = N5394 & N1415;
  assign N5627 = N5394 & idx_w_i[8];
  assign N5628 = N5396 & N1415;
  assign N5629 = N5396 & idx_w_i[8];
  assign N5630 = N5398 & N1415;
  assign N5631 = N5398 & idx_w_i[8];
  assign N5632 = N5400 & N1415;
  assign N5633 = N5400 & idx_w_i[8];
  assign N5634 = N5402 & N1415;
  assign N5635 = N5402 & idx_w_i[8];
  assign N5636 = N5404 & N1415;
  assign N5637 = N5404 & idx_w_i[8];
  assign N5638 = N5406 & N1415;
  assign N5639 = N5406 & idx_w_i[8];
  assign N5640 = N5408 & N1415;
  assign N5641 = N5408 & idx_w_i[8];
  assign N5642 = N5410 & N1415;
  assign N5643 = N5410 & idx_w_i[8];
  assign N5644 = N5412 & N1415;
  assign N5645 = N5412 & idx_w_i[8];
  assign N5646 = N5414 & N1415;
  assign N5647 = N5414 & idx_w_i[8];
  assign N5648 = N5416 & N1415;
  assign N5649 = N5416 & idx_w_i[8];
  assign N5650 = N5418 & N1415;
  assign N5651 = N5418 & idx_w_i[8];
  assign N5652 = N5420 & N1415;
  assign N5653 = N5420 & idx_w_i[8];
  assign N5654 = N5422 & N1415;
  assign N5655 = N5422 & idx_w_i[8];
  assign N5656 = N5424 & N1415;
  assign N5657 = N5424 & idx_w_i[8];
  assign N5658 = N5426 & N1415;
  assign N5659 = N5426 & idx_w_i[8];
  assign N5660 = N5428 & N1415;
  assign N5661 = N5428 & idx_w_i[8];
  assign N5662 = N5430 & N1415;
  assign N5663 = N5430 & idx_w_i[8];
  assign N5664 = N5432 & N1415;
  assign N5665 = N5432 & idx_w_i[8];
  assign N5666 = N5434 & N1415;
  assign N5667 = N5434 & idx_w_i[8];
  assign N5668 = N5436 & N1415;
  assign N5669 = N5436 & idx_w_i[8];
  assign N5670 = N5438 & N1415;
  assign N5671 = N5438 & idx_w_i[8];
  assign N5672 = N5439 & N1415;
  assign N5673 = N5439 & idx_w_i[8];
  assign N5674 = N5440 & N1415;
  assign N5675 = N5440 & idx_w_i[8];
  assign N5676 = N5441 & N1415;
  assign N5677 = N5441 & idx_w_i[8];
  assign N5678 = N5442 & N1415;
  assign N5679 = N5442 & idx_w_i[8];
  assign N5680 = N5443 & N1415;
  assign N5681 = N5443 & idx_w_i[8];
  assign N5682 = N5444 & N1415;
  assign N5683 = N5444 & idx_w_i[8];
  assign N5684 = N5445 & N1415;
  assign N5685 = N5445 & idx_w_i[8];
  assign N5686 = N5446 & N1415;
  assign N5687 = N5446 & idx_w_i[8];
  assign N5688 = N5447 & N1415;
  assign N5689 = N5447 & idx_w_i[8];
  assign N5690 = N5448 & N1415;
  assign N5691 = N5448 & idx_w_i[8];
  assign N5692 = N5449 & N1415;
  assign N5693 = N5449 & idx_w_i[8];
  assign N5694 = N5450 & N1415;
  assign N5695 = N5450 & idx_w_i[8];
  assign N5696 = N5451 & N1415;
  assign N5697 = N5451 & idx_w_i[8];
  assign N5698 = N5452 & N1415;
  assign N5699 = N5452 & idx_w_i[8];
  assign N5700 = N5453 & N1415;
  assign N5701 = N5453 & idx_w_i[8];
  assign N5702 = N5454 & N1415;
  assign N5703 = N5454 & idx_w_i[8];
  assign N5704 = N5455 & N1415;
  assign N5705 = N5455 & idx_w_i[8];
  assign N5706 = N5456 & N1415;
  assign N5707 = N5456 & idx_w_i[8];
  assign N5708 = N5457 & N1415;
  assign N5709 = N5457 & idx_w_i[8];
  assign N5710 = N5458 & N1415;
  assign N5711 = N5458 & idx_w_i[8];
  assign N5712 = N5459 & N1415;
  assign N5713 = N5459 & idx_w_i[8];
  assign N5714 = N5460 & N1415;
  assign N5715 = N5460 & idx_w_i[8];
  assign N5716 = N5461 & N1415;
  assign N5717 = N5461 & idx_w_i[8];
  assign N5718 = N5231 & N1415;
  assign N5719 = N5231 & idx_w_i[8];
  assign N5720 = N5233 & N1415;
  assign N5721 = N5233 & idx_w_i[8];
  assign N5722 = N5235 & N1415;
  assign N5723 = N5235 & idx_w_i[8];
  assign N5724 = N5237 & N1415;
  assign N5725 = N5237 & idx_w_i[8];
  assign N5726 = N5239 & N1415;
  assign N5727 = N5239 & idx_w_i[8];
  assign N5728 = N5241 & N1415;
  assign N5729 = N5241 & idx_w_i[8];
  assign N5730 = N5243 & N1415;
  assign N5731 = N5243 & idx_w_i[8];
  assign N5732 = N5245 & N1415;
  assign N5733 = N5245 & idx_w_i[8];
  assign N5734 = N5247 & N1415;
  assign N5735 = N5247 & idx_w_i[8];
  assign N5736 = N5249 & N1415;
  assign N5737 = N5249 & idx_w_i[8];
  assign N5738 = N5251 & N1415;
  assign N5739 = N5251 & idx_w_i[8];
  assign N5740 = N5253 & N1415;
  assign N5741 = N5253 & idx_w_i[8];
  assign N5742 = N5255 & N1415;
  assign N5743 = N5255 & idx_w_i[8];
  assign N5744 = N5257 & N1415;
  assign N5745 = N5257 & idx_w_i[8];
  assign N5746 = N5259 & N1415;
  assign N5747 = N5259 & idx_w_i[8];
  assign N5748 = N5261 & N1415;
  assign N5749 = N5261 & idx_w_i[8];
  assign N5750 = N5263 & N1415;
  assign N5751 = N5263 & idx_w_i[8];
  assign N5752 = N5265 & N1415;
  assign N5753 = N5265 & idx_w_i[8];
  assign N5754 = N5267 & N1415;
  assign N5755 = N5267 & idx_w_i[8];
  assign N5756 = N5269 & N1415;
  assign N5757 = N5269 & idx_w_i[8];
  assign N5758 = N5271 & N1415;
  assign N5759 = N5271 & idx_w_i[8];
  assign N5760 = N5273 & N1415;
  assign N5761 = N5273 & idx_w_i[8];
  assign N5762 = N5275 & N1415;
  assign N5763 = N5275 & idx_w_i[8];
  assign N5764 = N5277 & N1415;
  assign N5765 = N5277 & idx_w_i[8];
  assign N5766 = N5279 & N1415;
  assign N5767 = N5279 & idx_w_i[8];
  assign N5768 = N5281 & N1415;
  assign N5769 = N5281 & idx_w_i[8];
  assign N5770 = N5283 & N1415;
  assign N5771 = N5283 & idx_w_i[8];
  assign N5772 = N5285 & N1415;
  assign N5773 = N5285 & idx_w_i[8];
  assign N5774 = N5287 & N1415;
  assign N5775 = N5287 & idx_w_i[8];
  assign N5776 = N5289 & N1415;
  assign N5777 = N5289 & idx_w_i[8];
  assign N5778 = N5291 & N1415;
  assign N5779 = N5291 & idx_w_i[8];
  assign N5780 = N5293 & N1415;
  assign N5781 = N5293 & idx_w_i[8];
  assign N5782 = N5295 & N1415;
  assign N5783 = N5295 & idx_w_i[8];
  assign N5784 = N5297 & N1415;
  assign N5785 = N5297 & idx_w_i[8];
  assign N5786 = N5299 & N1415;
  assign N5787 = N5299 & idx_w_i[8];
  assign N5788 = N5301 & N1415;
  assign N5789 = N5301 & idx_w_i[8];
  assign N5790 = N5303 & N1415;
  assign N5791 = N5303 & idx_w_i[8];
  assign N5792 = N5305 & N1415;
  assign N5793 = N5305 & idx_w_i[8];
  assign N5794 = N5307 & N1415;
  assign N5795 = N5307 & idx_w_i[8];
  assign N5796 = N5309 & N1415;
  assign N5797 = N5309 & idx_w_i[8];
  assign N5798 = N5311 & N1415;
  assign N5799 = N5311 & idx_w_i[8];
  assign N5800 = N5313 & N1415;
  assign N5801 = N5313 & idx_w_i[8];
  assign N5802 = N5315 & N1415;
  assign N5803 = N5315 & idx_w_i[8];
  assign N5804 = N5317 & N1415;
  assign N5805 = N5317 & idx_w_i[8];
  assign N5806 = N5319 & N1415;
  assign N5807 = N5319 & idx_w_i[8];
  assign N5808 = N5321 & N1415;
  assign N5809 = N5321 & idx_w_i[8];
  assign N5810 = N5323 & N1415;
  assign N5811 = N5323 & idx_w_i[8];
  assign N5812 = N5325 & N1415;
  assign N5813 = N5325 & idx_w_i[8];
  assign N5814 = N5327 & N1415;
  assign N5815 = N5327 & idx_w_i[8];
  assign N5816 = N5329 & N1415;
  assign N5817 = N5329 & idx_w_i[8];
  assign N5818 = N5331 & N1415;
  assign N5819 = N5331 & idx_w_i[8];
  assign N5820 = N5333 & N1415;
  assign N5821 = N5333 & idx_w_i[8];
  assign N5822 = N5335 & N1415;
  assign N5823 = N5335 & idx_w_i[8];
  assign N5824 = N5337 & N1415;
  assign N5825 = N5337 & idx_w_i[8];
  assign N5826 = N5339 & N1415;
  assign N5827 = N5339 & idx_w_i[8];
  assign N5828 = N5341 & N1415;
  assign N5829 = N5341 & idx_w_i[8];
  assign N5830 = N5343 & N1415;
  assign N5831 = N5343 & idx_w_i[8];
  assign N5832 = N5345 & N1415;
  assign N5833 = N5345 & idx_w_i[8];
  assign N5834 = N5347 & N1415;
  assign N5835 = N5347 & idx_w_i[8];
  assign N5836 = N5349 & N1415;
  assign N5837 = N5349 & idx_w_i[8];
  assign N5838 = N5351 & N1415;
  assign N5839 = N5351 & idx_w_i[8];
  assign N5840 = N5353 & N1415;
  assign N5841 = N5353 & idx_w_i[8];
  assign N5842 = N5355 & N1415;
  assign N5843 = N5355 & idx_w_i[8];
  assign N5844 = N5357 & N1415;
  assign N5845 = N5357 & idx_w_i[8];
  assign N5846 = N5359 & N1415;
  assign N5847 = N5359 & idx_w_i[8];
  assign N5848 = N5361 & N1415;
  assign N5849 = N5361 & idx_w_i[8];
  assign N5850 = N5363 & N1415;
  assign N5851 = N5363 & idx_w_i[8];
  assign N5852 = N5365 & N1415;
  assign N5853 = N5365 & idx_w_i[8];
  assign N5854 = N5367 & N1415;
  assign N5855 = N5367 & idx_w_i[8];
  assign N5856 = N5369 & N1415;
  assign N5857 = N5369 & idx_w_i[8];
  assign N5858 = N5371 & N1415;
  assign N5859 = N5371 & idx_w_i[8];
  assign N5860 = N5373 & N1415;
  assign N5861 = N5373 & idx_w_i[8];
  assign N5862 = N5375 & N1415;
  assign N5863 = N5375 & idx_w_i[8];
  assign N5864 = N5377 & N1415;
  assign N5865 = N5377 & idx_w_i[8];
  assign N5866 = N5379 & N1415;
  assign N5867 = N5379 & idx_w_i[8];
  assign N5868 = N5381 & N1415;
  assign N5869 = N5381 & idx_w_i[8];
  assign N5870 = N5383 & N1415;
  assign N5871 = N5383 & idx_w_i[8];
  assign N5872 = N5385 & N1415;
  assign N5873 = N5385 & idx_w_i[8];
  assign N5874 = N5387 & N1415;
  assign N5875 = N5387 & idx_w_i[8];
  assign N5876 = N5389 & N1415;
  assign N5877 = N5389 & idx_w_i[8];
  assign N5878 = N5391 & N1415;
  assign N5879 = N5391 & idx_w_i[8];
  assign N5880 = N5393 & N1415;
  assign N5881 = N5393 & idx_w_i[8];
  assign N5882 = N5395 & N1415;
  assign N5883 = N5395 & idx_w_i[8];
  assign N5884 = N5397 & N1415;
  assign N5885 = N5397 & idx_w_i[8];
  assign N5886 = N5399 & N1415;
  assign N5887 = N5399 & idx_w_i[8];
  assign N5888 = N5401 & N1415;
  assign N5889 = N5401 & idx_w_i[8];
  assign N5890 = N5403 & N1415;
  assign N5891 = N5403 & idx_w_i[8];
  assign N5892 = N5405 & N1415;
  assign N5893 = N5405 & idx_w_i[8];
  assign N5894 = N5407 & N1415;
  assign N5895 = N5407 & idx_w_i[8];
  assign N5896 = N5409 & N1415;
  assign N5897 = N5409 & idx_w_i[8];
  assign N5898 = N5411 & N1415;
  assign N5899 = N5411 & idx_w_i[8];
  assign N5900 = N5413 & N1415;
  assign N5901 = N5413 & idx_w_i[8];
  assign N5902 = N5415 & N1415;
  assign N5903 = N5415 & idx_w_i[8];
  assign N5904 = N5417 & N1415;
  assign N5905 = N5417 & idx_w_i[8];
  assign N5906 = N5419 & N1415;
  assign N5907 = N5419 & idx_w_i[8];
  assign N5908 = N5421 & N1415;
  assign N5909 = N5421 & idx_w_i[8];
  assign N5910 = N5423 & N1415;
  assign N5911 = N5423 & idx_w_i[8];
  assign N5912 = N5425 & N1415;
  assign N5913 = N5425 & idx_w_i[8];
  assign N5914 = N5427 & N1415;
  assign N5915 = N5427 & idx_w_i[8];
  assign N5916 = N5429 & N1415;
  assign N5917 = N5429 & idx_w_i[8];
  assign N5918 = N5431 & N1415;
  assign N5919 = N5431 & idx_w_i[8];
  assign N5920 = N5433 & N1415;
  assign N5921 = N5433 & idx_w_i[8];
  assign N5922 = N5435 & N1415;
  assign N5923 = N5435 & idx_w_i[8];
  assign N5924 = N5437 & N1415;
  assign N5925 = N5437 & idx_w_i[8];
  assign N5926 = N4037 & N1415;
  assign N5927 = N4039 & N1415;
  assign N5928 = N4041 & N1415;
  assign N5929 = N4043 & N1415;
  assign N5930 = N4045 & N1415;
  assign N5931 = N4047 & N1415;
  assign N5932 = N4049 & N1415;
  assign N5933 = N4051 & N1415;
  assign N5934 = N11569 & N1415;
  assign N5935 = N11571 & N1415;
  assign N5936 = N11573 & N1415;
  assign N5937 = N11575 & N1415;
  assign N5938 = N11577 & N1415;
  assign N5939 = N11579 & N1415;
  assign N5940 = N11581 & N1415;
  assign N5941 = N11583 & N1415;
  assign N5942 = N11585 & N1415;
  assign N5943 = N11587 & N1415;
  assign N5944 = N11589 & N1415;
  assign N5945 = N11591 & N1415;
  assign N5946 = N11593 & N1415;
  assign N5947 = N11595 & N1415;
  assign N5948 = N11597 & N1415;
  assign N5949 = N11599 & N1415;
  assign N5951 = N11104 & N2698;
  assign N5952 = N11106 & N2698;
  assign N5953 = N11108 & N2698;
  assign N5954 = N11110 & N2698;
  assign N5955 = N11112 & N2698;
  assign N5956 = N11114 & N2698;
  assign N5957 = N11116 & N2698;
  assign N5958 = N11118 & N2698;
  assign N5959 = N5951 & N1060;
  assign N5960 = N5951 & idx_w_i[5];
  assign N5961 = N5952 & N1060;
  assign N5962 = N5952 & idx_w_i[5];
  assign N5963 = N5953 & N1060;
  assign N5964 = N5953 & idx_w_i[5];
  assign N5965 = N5954 & N1060;
  assign N5966 = N5954 & idx_w_i[5];
  assign N5967 = N5955 & N1060;
  assign N5968 = N5955 & idx_w_i[5];
  assign N5969 = N5956 & N1060;
  assign N5970 = N5956 & idx_w_i[5];
  assign N5971 = N5957 & N1060;
  assign N5972 = N5957 & idx_w_i[5];
  assign N5973 = N5958 & N1060;
  assign N5974 = N5958 & idx_w_i[5];
  assign N5975 = N2715 & N1060;
  assign N5976 = N2716 & N1060;
  assign N5977 = N2717 & N1060;
  assign N5978 = N2718 & N1060;
  assign N5979 = N2719 & N1060;
  assign N5980 = N2720 & N1060;
  assign N5981 = N2721 & N1060;
  assign N5982 = N2722 & N1060;
  assign N5983 = N5959 & N1093;
  assign N5984 = N5959 & idx_w_i[6];
  assign N5985 = N5961 & N1093;
  assign N5986 = N5961 & idx_w_i[6];
  assign N5987 = N5963 & N1093;
  assign N5988 = N5963 & idx_w_i[6];
  assign N5989 = N5965 & N1093;
  assign N5990 = N5965 & idx_w_i[6];
  assign N5991 = N5967 & N1093;
  assign N5992 = N5967 & idx_w_i[6];
  assign N5993 = N5969 & N1093;
  assign N5994 = N5969 & idx_w_i[6];
  assign N5995 = N5971 & N1093;
  assign N5996 = N5971 & idx_w_i[6];
  assign N5997 = N5973 & N1093;
  assign N5998 = N5973 & idx_w_i[6];
  assign N5999 = N5975 & N1093;
  assign N6000 = N5975 & idx_w_i[6];
  assign N6001 = N5976 & N1093;
  assign N6002 = N5976 & idx_w_i[6];
  assign N6003 = N5977 & N1093;
  assign N6004 = N5977 & idx_w_i[6];
  assign N6005 = N5978 & N1093;
  assign N6006 = N5978 & idx_w_i[6];
  assign N6007 = N5979 & N1093;
  assign N6008 = N5979 & idx_w_i[6];
  assign N6009 = N5980 & N1093;
  assign N6010 = N5980 & idx_w_i[6];
  assign N6011 = N5981 & N1093;
  assign N6012 = N5981 & idx_w_i[6];
  assign N6013 = N5982 & N1093;
  assign N6014 = N5982 & idx_w_i[6];
  assign N6015 = N5110 & N1093;
  assign N6016 = N5111 & N1093;
  assign N6017 = N5112 & N1093;
  assign N6018 = N5113 & N1093;
  assign N6019 = N5114 & N1093;
  assign N6020 = N5115 & N1093;
  assign N6021 = N5116 & N1093;
  assign N6022 = N5117 & N1093;
  assign N6023 = N5118 & N1093;
  assign N6024 = N5119 & N1093;
  assign N6025 = N5120 & N1093;
  assign N6026 = N5121 & N1093;
  assign N6027 = N5122 & N1093;
  assign N6028 = N5123 & N1093;
  assign N6029 = N5124 & N1093;
  assign N6030 = N5125 & N1093;
  assign N6031 = N5960 & N1093;
  assign N6032 = N5960 & idx_w_i[6];
  assign N6033 = N5962 & N1093;
  assign N6034 = N5962 & idx_w_i[6];
  assign N6035 = N5964 & N1093;
  assign N6036 = N5964 & idx_w_i[6];
  assign N6037 = N5966 & N1093;
  assign N6038 = N5966 & idx_w_i[6];
  assign N6039 = N5968 & N1093;
  assign N6040 = N5968 & idx_w_i[6];
  assign N6041 = N5970 & N1093;
  assign N6042 = N5970 & idx_w_i[6];
  assign N6043 = N5972 & N1093;
  assign N6044 = N5972 & idx_w_i[6];
  assign N6045 = N5974 & N1093;
  assign N6046 = N5974 & idx_w_i[6];
  assign N6047 = N2740 & N1093;
  assign N6048 = N2742 & N1093;
  assign N6049 = N2744 & N1093;
  assign N6050 = N2746 & N1093;
  assign N6051 = N2748 & N1093;
  assign N6052 = N2750 & N1093;
  assign N6053 = N2752 & N1093;
  assign N6054 = N2754 & N1093;
  assign N6055 = N11185 & N1093;
  assign N6056 = N11187 & N1093;
  assign N6057 = N11189 & N1093;
  assign N6058 = N11191 & N1093;
  assign N6059 = N11193 & N1093;
  assign N6060 = N11195 & N1093;
  assign N6061 = N11197 & N1093;
  assign N6062 = N11199 & N1093;
  assign N6063 = N11201 & N1093;
  assign N6064 = N11203 & N1093;
  assign N6065 = N11205 & N1093;
  assign N6066 = N11207 & N1093;
  assign N6067 = N11209 & N1093;
  assign N6068 = N11211 & N1093;
  assign N6069 = N11213 & N1093;
  assign N6070 = N11215 & N1093;
  assign N6071 = N5983 & N1190;
  assign N6072 = N5983 & idx_w_i[7];
  assign N6073 = N5985 & N1190;
  assign N6074 = N5985 & idx_w_i[7];
  assign N6075 = N5987 & N1190;
  assign N6076 = N5987 & idx_w_i[7];
  assign N6077 = N5989 & N1190;
  assign N6078 = N5989 & idx_w_i[7];
  assign N6079 = N5991 & N1190;
  assign N6080 = N5991 & idx_w_i[7];
  assign N6081 = N5993 & N1190;
  assign N6082 = N5993 & idx_w_i[7];
  assign N6083 = N5995 & N1190;
  assign N6084 = N5995 & idx_w_i[7];
  assign N6085 = N5997 & N1190;
  assign N6086 = N5997 & idx_w_i[7];
  assign N6087 = N5999 & N1190;
  assign N6088 = N5999 & idx_w_i[7];
  assign N6089 = N6001 & N1190;
  assign N6090 = N6001 & idx_w_i[7];
  assign N6091 = N6003 & N1190;
  assign N6092 = N6003 & idx_w_i[7];
  assign N6093 = N6005 & N1190;
  assign N6094 = N6005 & idx_w_i[7];
  assign N6095 = N6007 & N1190;
  assign N6096 = N6007 & idx_w_i[7];
  assign N6097 = N6009 & N1190;
  assign N6098 = N6009 & idx_w_i[7];
  assign N6099 = N6011 & N1190;
  assign N6100 = N6011 & idx_w_i[7];
  assign N6101 = N6013 & N1190;
  assign N6102 = N6013 & idx_w_i[7];
  assign N6103 = N6015 & N1190;
  assign N6104 = N6015 & idx_w_i[7];
  assign N6105 = N6016 & N1190;
  assign N6106 = N6016 & idx_w_i[7];
  assign N6107 = N6017 & N1190;
  assign N6108 = N6017 & idx_w_i[7];
  assign N6109 = N6018 & N1190;
  assign N6110 = N6018 & idx_w_i[7];
  assign N6111 = N6019 & N1190;
  assign N6112 = N6019 & idx_w_i[7];
  assign N6113 = N6020 & N1190;
  assign N6114 = N6020 & idx_w_i[7];
  assign N6115 = N6021 & N1190;
  assign N6116 = N6021 & idx_w_i[7];
  assign N6117 = N6022 & N1190;
  assign N6118 = N6022 & idx_w_i[7];
  assign N6119 = N6023 & N1190;
  assign N6120 = N6023 & idx_w_i[7];
  assign N6121 = N6024 & N1190;
  assign N6122 = N6024 & idx_w_i[7];
  assign N6123 = N6025 & N1190;
  assign N6124 = N6025 & idx_w_i[7];
  assign N6125 = N6026 & N1190;
  assign N6126 = N6026 & idx_w_i[7];
  assign N6127 = N6027 & N1190;
  assign N6128 = N6027 & idx_w_i[7];
  assign N6129 = N6028 & N1190;
  assign N6130 = N6028 & idx_w_i[7];
  assign N6131 = N6029 & N1190;
  assign N6132 = N6029 & idx_w_i[7];
  assign N6133 = N6030 & N1190;
  assign N6134 = N6030 & idx_w_i[7];
  assign N6135 = N6031 & N1190;
  assign N6136 = N6031 & idx_w_i[7];
  assign N6137 = N6033 & N1190;
  assign N6138 = N6033 & idx_w_i[7];
  assign N6139 = N6035 & N1190;
  assign N6140 = N6035 & idx_w_i[7];
  assign N6141 = N6037 & N1190;
  assign N6142 = N6037 & idx_w_i[7];
  assign N6143 = N6039 & N1190;
  assign N6144 = N6039 & idx_w_i[7];
  assign N6145 = N6041 & N1190;
  assign N6146 = N6041 & idx_w_i[7];
  assign N6147 = N6043 & N1190;
  assign N6148 = N6043 & idx_w_i[7];
  assign N6149 = N6045 & N1190;
  assign N6150 = N6045 & idx_w_i[7];
  assign N6151 = N6047 & N1190;
  assign N6152 = N6047 & idx_w_i[7];
  assign N6153 = N6048 & N1190;
  assign N6154 = N6048 & idx_w_i[7];
  assign N6155 = N6049 & N1190;
  assign N6156 = N6049 & idx_w_i[7];
  assign N6157 = N6050 & N1190;
  assign N6158 = N6050 & idx_w_i[7];
  assign N6159 = N6051 & N1190;
  assign N6160 = N6051 & idx_w_i[7];
  assign N6161 = N6052 & N1190;
  assign N6162 = N6052 & idx_w_i[7];
  assign N6163 = N6053 & N1190;
  assign N6164 = N6053 & idx_w_i[7];
  assign N6165 = N6054 & N1190;
  assign N6166 = N6054 & idx_w_i[7];
  assign N6167 = N6055 & N1190;
  assign N6168 = N6055 & idx_w_i[7];
  assign N6169 = N6056 & N1190;
  assign N6170 = N6056 & idx_w_i[7];
  assign N6171 = N6057 & N1190;
  assign N6172 = N6057 & idx_w_i[7];
  assign N6173 = N6058 & N1190;
  assign N6174 = N6058 & idx_w_i[7];
  assign N6175 = N6059 & N1190;
  assign N6176 = N6059 & idx_w_i[7];
  assign N6177 = N6060 & N1190;
  assign N6178 = N6060 & idx_w_i[7];
  assign N6179 = N6061 & N1190;
  assign N6180 = N6061 & idx_w_i[7];
  assign N6181 = N6062 & N1190;
  assign N6182 = N6062 & idx_w_i[7];
  assign N6183 = N6063 & N1190;
  assign N6184 = N6063 & idx_w_i[7];
  assign N6185 = N6064 & N1190;
  assign N6186 = N6064 & idx_w_i[7];
  assign N6187 = N6065 & N1190;
  assign N6188 = N6065 & idx_w_i[7];
  assign N6189 = N6066 & N1190;
  assign N6190 = N6066 & idx_w_i[7];
  assign N6191 = N6067 & N1190;
  assign N6192 = N6067 & idx_w_i[7];
  assign N6193 = N6068 & N1190;
  assign N6194 = N6068 & idx_w_i[7];
  assign N6195 = N6069 & N1190;
  assign N6196 = N6069 & idx_w_i[7];
  assign N6197 = N6070 & N1190;
  assign N6198 = N6070 & idx_w_i[7];
  assign N6199 = N5984 & N1190;
  assign N6200 = N5984 & idx_w_i[7];
  assign N6201 = N5986 & N1190;
  assign N6202 = N5986 & idx_w_i[7];
  assign N6203 = N5988 & N1190;
  assign N6204 = N5988 & idx_w_i[7];
  assign N6205 = N5990 & N1190;
  assign N6206 = N5990 & idx_w_i[7];
  assign N6207 = N5992 & N1190;
  assign N6208 = N5992 & idx_w_i[7];
  assign N6209 = N5994 & N1190;
  assign N6210 = N5994 & idx_w_i[7];
  assign N6211 = N5996 & N1190;
  assign N6212 = N5996 & idx_w_i[7];
  assign N6213 = N5998 & N1190;
  assign N6214 = N5998 & idx_w_i[7];
  assign N6215 = N6000 & N1190;
  assign N6216 = N6000 & idx_w_i[7];
  assign N6217 = N6002 & N1190;
  assign N6218 = N6002 & idx_w_i[7];
  assign N6219 = N6004 & N1190;
  assign N6220 = N6004 & idx_w_i[7];
  assign N6221 = N6006 & N1190;
  assign N6222 = N6006 & idx_w_i[7];
  assign N6223 = N6008 & N1190;
  assign N6224 = N6008 & idx_w_i[7];
  assign N6225 = N6010 & N1190;
  assign N6226 = N6010 & idx_w_i[7];
  assign N6227 = N6012 & N1190;
  assign N6228 = N6012 & idx_w_i[7];
  assign N6229 = N6014 & N1190;
  assign N6230 = N6014 & idx_w_i[7];
  assign N6231 = N5159 & N1190;
  assign N6232 = N5161 & N1190;
  assign N6233 = N5163 & N1190;
  assign N6234 = N5165 & N1190;
  assign N6235 = N5167 & N1190;
  assign N6236 = N5169 & N1190;
  assign N6237 = N5171 & N1190;
  assign N6238 = N5173 & N1190;
  assign N6239 = N5175 & N1190;
  assign N6240 = N5177 & N1190;
  assign N6241 = N5179 & N1190;
  assign N6242 = N5181 & N1190;
  assign N6243 = N5183 & N1190;
  assign N6244 = N5185 & N1190;
  assign N6245 = N5187 & N1190;
  assign N6246 = N5189 & N1190;
  assign N6247 = N6032 & N1190;
  assign N6248 = N6032 & idx_w_i[7];
  assign N6249 = N6034 & N1190;
  assign N6250 = N6034 & idx_w_i[7];
  assign N6251 = N6036 & N1190;
  assign N6252 = N6036 & idx_w_i[7];
  assign N6253 = N6038 & N1190;
  assign N6254 = N6038 & idx_w_i[7];
  assign N6255 = N6040 & N1190;
  assign N6256 = N6040 & idx_w_i[7];
  assign N6257 = N6042 & N1190;
  assign N6258 = N6042 & idx_w_i[7];
  assign N6259 = N6044 & N1190;
  assign N6260 = N6044 & idx_w_i[7];
  assign N6261 = N6046 & N1190;
  assign N6262 = N6046 & idx_w_i[7];
  assign N6263 = N2860 & N1190;
  assign N6264 = N2862 & N1190;
  assign N6265 = N2864 & N1190;
  assign N6266 = N2866 & N1190;
  assign N6267 = N2868 & N1190;
  assign N6268 = N2870 & N1190;
  assign N6269 = N2872 & N1190;
  assign N6270 = N2874 & N1190;
  assign N6271 = N11313 & N1190;
  assign N6272 = N11315 & N1190;
  assign N6273 = N11317 & N1190;
  assign N6274 = N11319 & N1190;
  assign N6275 = N11321 & N1190;
  assign N6276 = N11323 & N1190;
  assign N6277 = N11325 & N1190;
  assign N6278 = N11327 & N1190;
  assign N6279 = N11329 & N1190;
  assign N6280 = N11331 & N1190;
  assign N6281 = N11333 & N1190;
  assign N6282 = N11335 & N1190;
  assign N6283 = N11337 & N1190;
  assign N6284 = N11339 & N1190;
  assign N6285 = N11341 & N1190;
  assign N6286 = N11343 & N1190;
  assign N6287 = N6071 & N1415;
  assign N6288 = N6071 & idx_w_i[8];
  assign N6289 = N6073 & N1415;
  assign N6290 = N6073 & idx_w_i[8];
  assign N6291 = N6075 & N1415;
  assign N6292 = N6075 & idx_w_i[8];
  assign N6293 = N6077 & N1415;
  assign N6294 = N6077 & idx_w_i[8];
  assign N6295 = N6079 & N1415;
  assign N6296 = N6079 & idx_w_i[8];
  assign N6297 = N6081 & N1415;
  assign N6298 = N6081 & idx_w_i[8];
  assign N6299 = N6083 & N1415;
  assign N6300 = N6083 & idx_w_i[8];
  assign N6301 = N6085 & N1415;
  assign N6302 = N6085 & idx_w_i[8];
  assign N6303 = N6087 & N1415;
  assign N6304 = N6087 & idx_w_i[8];
  assign N6305 = N6089 & N1415;
  assign N6306 = N6089 & idx_w_i[8];
  assign N6307 = N6091 & N1415;
  assign N6308 = N6091 & idx_w_i[8];
  assign N6309 = N6093 & N1415;
  assign N6310 = N6093 & idx_w_i[8];
  assign N6311 = N6095 & N1415;
  assign N6312 = N6095 & idx_w_i[8];
  assign N6313 = N6097 & N1415;
  assign N6314 = N6097 & idx_w_i[8];
  assign N6315 = N6099 & N1415;
  assign N6316 = N6099 & idx_w_i[8];
  assign N6317 = N6101 & N1415;
  assign N6318 = N6101 & idx_w_i[8];
  assign N6319 = N6103 & N1415;
  assign N6320 = N6103 & idx_w_i[8];
  assign N6321 = N6105 & N1415;
  assign N6322 = N6105 & idx_w_i[8];
  assign N6323 = N6107 & N1415;
  assign N6324 = N6107 & idx_w_i[8];
  assign N6325 = N6109 & N1415;
  assign N6326 = N6109 & idx_w_i[8];
  assign N6327 = N6111 & N1415;
  assign N6328 = N6111 & idx_w_i[8];
  assign N6329 = N6113 & N1415;
  assign N6330 = N6113 & idx_w_i[8];
  assign N6331 = N6115 & N1415;
  assign N6332 = N6115 & idx_w_i[8];
  assign N6333 = N6117 & N1415;
  assign N6334 = N6117 & idx_w_i[8];
  assign N6335 = N6119 & N1415;
  assign N6336 = N6119 & idx_w_i[8];
  assign N6337 = N6121 & N1415;
  assign N6338 = N6121 & idx_w_i[8];
  assign N6339 = N6123 & N1415;
  assign N6340 = N6123 & idx_w_i[8];
  assign N6341 = N6125 & N1415;
  assign N6342 = N6125 & idx_w_i[8];
  assign N6343 = N6127 & N1415;
  assign N6344 = N6127 & idx_w_i[8];
  assign N6345 = N6129 & N1415;
  assign N6346 = N6129 & idx_w_i[8];
  assign N6347 = N6131 & N1415;
  assign N6348 = N6131 & idx_w_i[8];
  assign N6349 = N6133 & N1415;
  assign N6350 = N6133 & idx_w_i[8];
  assign N6351 = N6135 & N1415;
  assign N6352 = N6135 & idx_w_i[8];
  assign N6353 = N6137 & N1415;
  assign N6354 = N6137 & idx_w_i[8];
  assign N6355 = N6139 & N1415;
  assign N6356 = N6139 & idx_w_i[8];
  assign N6357 = N6141 & N1415;
  assign N6358 = N6141 & idx_w_i[8];
  assign N6359 = N6143 & N1415;
  assign N6360 = N6143 & idx_w_i[8];
  assign N6361 = N6145 & N1415;
  assign N6362 = N6145 & idx_w_i[8];
  assign N6363 = N6147 & N1415;
  assign N6364 = N6147 & idx_w_i[8];
  assign N6365 = N6149 & N1415;
  assign N6366 = N6149 & idx_w_i[8];
  assign N6367 = N6151 & N1415;
  assign N6368 = N6151 & idx_w_i[8];
  assign N6369 = N6153 & N1415;
  assign N6370 = N6153 & idx_w_i[8];
  assign N6371 = N6155 & N1415;
  assign N6372 = N6155 & idx_w_i[8];
  assign N6373 = N6157 & N1415;
  assign N6374 = N6157 & idx_w_i[8];
  assign N6375 = N6159 & N1415;
  assign N6376 = N6159 & idx_w_i[8];
  assign N6377 = N6161 & N1415;
  assign N6378 = N6161 & idx_w_i[8];
  assign N6379 = N6163 & N1415;
  assign N6380 = N6163 & idx_w_i[8];
  assign N6381 = N6165 & N1415;
  assign N6382 = N6165 & idx_w_i[8];
  assign N6383 = N6167 & N1415;
  assign N6384 = N6167 & idx_w_i[8];
  assign N6385 = N6169 & N1415;
  assign N6386 = N6169 & idx_w_i[8];
  assign N6387 = N6171 & N1415;
  assign N6388 = N6171 & idx_w_i[8];
  assign N6389 = N6173 & N1415;
  assign N6390 = N6173 & idx_w_i[8];
  assign N6391 = N6175 & N1415;
  assign N6392 = N6175 & idx_w_i[8];
  assign N6393 = N6177 & N1415;
  assign N6394 = N6177 & idx_w_i[8];
  assign N6395 = N6179 & N1415;
  assign N6396 = N6179 & idx_w_i[8];
  assign N6397 = N6181 & N1415;
  assign N6398 = N6181 & idx_w_i[8];
  assign N6399 = N6183 & N1415;
  assign N6400 = N6183 & idx_w_i[8];
  assign N6401 = N6185 & N1415;
  assign N6402 = N6185 & idx_w_i[8];
  assign N6403 = N6187 & N1415;
  assign N6404 = N6187 & idx_w_i[8];
  assign N6405 = N6189 & N1415;
  assign N6406 = N6189 & idx_w_i[8];
  assign N6407 = N6191 & N1415;
  assign N6408 = N6191 & idx_w_i[8];
  assign N6409 = N6193 & N1415;
  assign N6410 = N6193 & idx_w_i[8];
  assign N6411 = N6195 & N1415;
  assign N6412 = N6195 & idx_w_i[8];
  assign N6413 = N6197 & N1415;
  assign N6414 = N6197 & idx_w_i[8];
  assign N6415 = N6199 & N1415;
  assign N6416 = N6199 & idx_w_i[8];
  assign N6417 = N6201 & N1415;
  assign N6418 = N6201 & idx_w_i[8];
  assign N6419 = N6203 & N1415;
  assign N6420 = N6203 & idx_w_i[8];
  assign N6421 = N6205 & N1415;
  assign N6422 = N6205 & idx_w_i[8];
  assign N6423 = N6207 & N1415;
  assign N6424 = N6207 & idx_w_i[8];
  assign N6425 = N6209 & N1415;
  assign N6426 = N6209 & idx_w_i[8];
  assign N6427 = N6211 & N1415;
  assign N6428 = N6211 & idx_w_i[8];
  assign N6429 = N6213 & N1415;
  assign N6430 = N6213 & idx_w_i[8];
  assign N6431 = N6215 & N1415;
  assign N6432 = N6215 & idx_w_i[8];
  assign N6433 = N6217 & N1415;
  assign N6434 = N6217 & idx_w_i[8];
  assign N6435 = N6219 & N1415;
  assign N6436 = N6219 & idx_w_i[8];
  assign N6437 = N6221 & N1415;
  assign N6438 = N6221 & idx_w_i[8];
  assign N6439 = N6223 & N1415;
  assign N6440 = N6223 & idx_w_i[8];
  assign N6441 = N6225 & N1415;
  assign N6442 = N6225 & idx_w_i[8];
  assign N6443 = N6227 & N1415;
  assign N6444 = N6227 & idx_w_i[8];
  assign N6445 = N6229 & N1415;
  assign N6446 = N6229 & idx_w_i[8];
  assign N6447 = N6231 & N1415;
  assign N6448 = N6231 & idx_w_i[8];
  assign N6449 = N6232 & N1415;
  assign N6450 = N6232 & idx_w_i[8];
  assign N6451 = N6233 & N1415;
  assign N6452 = N6233 & idx_w_i[8];
  assign N6453 = N6234 & N1415;
  assign N6454 = N6234 & idx_w_i[8];
  assign N6455 = N6235 & N1415;
  assign N6456 = N6235 & idx_w_i[8];
  assign N6457 = N6236 & N1415;
  assign N6458 = N6236 & idx_w_i[8];
  assign N6459 = N6237 & N1415;
  assign N6460 = N6237 & idx_w_i[8];
  assign N6461 = N6238 & N1415;
  assign N6462 = N6238 & idx_w_i[8];
  assign N6463 = N6239 & N1415;
  assign N6464 = N6239 & idx_w_i[8];
  assign N6465 = N6240 & N1415;
  assign N6466 = N6240 & idx_w_i[8];
  assign N6467 = N6241 & N1415;
  assign N6468 = N6241 & idx_w_i[8];
  assign N6469 = N6242 & N1415;
  assign N6470 = N6242 & idx_w_i[8];
  assign N6471 = N6243 & N1415;
  assign N6472 = N6243 & idx_w_i[8];
  assign N6473 = N6244 & N1415;
  assign N6474 = N6244 & idx_w_i[8];
  assign N6475 = N6245 & N1415;
  assign N6476 = N6245 & idx_w_i[8];
  assign N6477 = N6246 & N1415;
  assign N6478 = N6246 & idx_w_i[8];
  assign N6479 = N6247 & N1415;
  assign N6480 = N6247 & idx_w_i[8];
  assign N6481 = N6249 & N1415;
  assign N6482 = N6249 & idx_w_i[8];
  assign N6483 = N6251 & N1415;
  assign N6484 = N6251 & idx_w_i[8];
  assign N6485 = N6253 & N1415;
  assign N6486 = N6253 & idx_w_i[8];
  assign N6487 = N6255 & N1415;
  assign N6488 = N6255 & idx_w_i[8];
  assign N6489 = N6257 & N1415;
  assign N6490 = N6257 & idx_w_i[8];
  assign N6491 = N6259 & N1415;
  assign N6492 = N6259 & idx_w_i[8];
  assign N6493 = N6261 & N1415;
  assign N6494 = N6261 & idx_w_i[8];
  assign N6495 = N6263 & N1415;
  assign N6496 = N6263 & idx_w_i[8];
  assign N6497 = N6264 & N1415;
  assign N6498 = N6264 & idx_w_i[8];
  assign N6499 = N6265 & N1415;
  assign N6500 = N6265 & idx_w_i[8];
  assign N6501 = N6266 & N1415;
  assign N6502 = N6266 & idx_w_i[8];
  assign N6503 = N6267 & N1415;
  assign N6504 = N6267 & idx_w_i[8];
  assign N6505 = N6268 & N1415;
  assign N6506 = N6268 & idx_w_i[8];
  assign N6507 = N6269 & N1415;
  assign N6508 = N6269 & idx_w_i[8];
  assign N6509 = N6270 & N1415;
  assign N6510 = N6270 & idx_w_i[8];
  assign N6511 = N6271 & N1415;
  assign N6512 = N6271 & idx_w_i[8];
  assign N6513 = N6272 & N1415;
  assign N6514 = N6272 & idx_w_i[8];
  assign N6515 = N6273 & N1415;
  assign N6516 = N6273 & idx_w_i[8];
  assign N6517 = N6274 & N1415;
  assign N6518 = N6274 & idx_w_i[8];
  assign N6519 = N6275 & N1415;
  assign N6520 = N6275 & idx_w_i[8];
  assign N6521 = N6276 & N1415;
  assign N6522 = N6276 & idx_w_i[8];
  assign N6523 = N6277 & N1415;
  assign N6524 = N6277 & idx_w_i[8];
  assign N6525 = N6278 & N1415;
  assign N6526 = N6278 & idx_w_i[8];
  assign N6527 = N6279 & N1415;
  assign N6528 = N6279 & idx_w_i[8];
  assign N6529 = N6280 & N1415;
  assign N6530 = N6280 & idx_w_i[8];
  assign N6531 = N6281 & N1415;
  assign N6532 = N6281 & idx_w_i[8];
  assign N6533 = N6282 & N1415;
  assign N6534 = N6282 & idx_w_i[8];
  assign N6535 = N6283 & N1415;
  assign N6536 = N6283 & idx_w_i[8];
  assign N6537 = N6284 & N1415;
  assign N6538 = N6284 & idx_w_i[8];
  assign N6539 = N6285 & N1415;
  assign N6540 = N6285 & idx_w_i[8];
  assign N6541 = N6286 & N1415;
  assign N6542 = N6286 & idx_w_i[8];
  assign N6543 = N6072 & N1415;
  assign N6544 = N6072 & idx_w_i[8];
  assign N6545 = N6074 & N1415;
  assign N6546 = N6074 & idx_w_i[8];
  assign N6547 = N6076 & N1415;
  assign N6548 = N6076 & idx_w_i[8];
  assign N6549 = N6078 & N1415;
  assign N6550 = N6078 & idx_w_i[8];
  assign N6551 = N6080 & N1415;
  assign N6552 = N6080 & idx_w_i[8];
  assign N6553 = N6082 & N1415;
  assign N6554 = N6082 & idx_w_i[8];
  assign N6555 = N6084 & N1415;
  assign N6556 = N6084 & idx_w_i[8];
  assign N6557 = N6086 & N1415;
  assign N6558 = N6086 & idx_w_i[8];
  assign N6559 = N6088 & N1415;
  assign N6560 = N6088 & idx_w_i[8];
  assign N6561 = N6090 & N1415;
  assign N6562 = N6090 & idx_w_i[8];
  assign N6563 = N6092 & N1415;
  assign N6564 = N6092 & idx_w_i[8];
  assign N6565 = N6094 & N1415;
  assign N6566 = N6094 & idx_w_i[8];
  assign N6567 = N6096 & N1415;
  assign N6568 = N6096 & idx_w_i[8];
  assign N6569 = N6098 & N1415;
  assign N6570 = N6098 & idx_w_i[8];
  assign N6571 = N6100 & N1415;
  assign N6572 = N6100 & idx_w_i[8];
  assign N6573 = N6102 & N1415;
  assign N6574 = N6102 & idx_w_i[8];
  assign N6575 = N6104 & N1415;
  assign N6576 = N6104 & idx_w_i[8];
  assign N6577 = N6106 & N1415;
  assign N6578 = N6106 & idx_w_i[8];
  assign N6579 = N6108 & N1415;
  assign N6580 = N6108 & idx_w_i[8];
  assign N6581 = N6110 & N1415;
  assign N6582 = N6110 & idx_w_i[8];
  assign N6583 = N6112 & N1415;
  assign N6584 = N6112 & idx_w_i[8];
  assign N6585 = N6114 & N1415;
  assign N6586 = N6114 & idx_w_i[8];
  assign N6587 = N6116 & N1415;
  assign N6588 = N6116 & idx_w_i[8];
  assign N6589 = N6118 & N1415;
  assign N6590 = N6118 & idx_w_i[8];
  assign N6591 = N6120 & N1415;
  assign N6592 = N6120 & idx_w_i[8];
  assign N6593 = N6122 & N1415;
  assign N6594 = N6122 & idx_w_i[8];
  assign N6595 = N6124 & N1415;
  assign N6596 = N6124 & idx_w_i[8];
  assign N6597 = N6126 & N1415;
  assign N6598 = N6126 & idx_w_i[8];
  assign N6599 = N6128 & N1415;
  assign N6600 = N6128 & idx_w_i[8];
  assign N6601 = N6130 & N1415;
  assign N6602 = N6130 & idx_w_i[8];
  assign N6603 = N6132 & N1415;
  assign N6604 = N6132 & idx_w_i[8];
  assign N6605 = N6134 & N1415;
  assign N6606 = N6134 & idx_w_i[8];
  assign N6607 = N6136 & N1415;
  assign N6608 = N6136 & idx_w_i[8];
  assign N6609 = N6138 & N1415;
  assign N6610 = N6138 & idx_w_i[8];
  assign N6611 = N6140 & N1415;
  assign N6612 = N6140 & idx_w_i[8];
  assign N6613 = N6142 & N1415;
  assign N6614 = N6142 & idx_w_i[8];
  assign N6615 = N6144 & N1415;
  assign N6616 = N6144 & idx_w_i[8];
  assign N6617 = N6146 & N1415;
  assign N6618 = N6146 & idx_w_i[8];
  assign N6619 = N6148 & N1415;
  assign N6620 = N6148 & idx_w_i[8];
  assign N6621 = N6150 & N1415;
  assign N6622 = N6150 & idx_w_i[8];
  assign N6623 = N6152 & N1415;
  assign N6624 = N6152 & idx_w_i[8];
  assign N6625 = N6154 & N1415;
  assign N6626 = N6154 & idx_w_i[8];
  assign N6627 = N6156 & N1415;
  assign N6628 = N6156 & idx_w_i[8];
  assign N6629 = N6158 & N1415;
  assign N6630 = N6158 & idx_w_i[8];
  assign N6631 = N6160 & N1415;
  assign N6632 = N6160 & idx_w_i[8];
  assign N6633 = N6162 & N1415;
  assign N6634 = N6162 & idx_w_i[8];
  assign N6635 = N6164 & N1415;
  assign N6636 = N6164 & idx_w_i[8];
  assign N6637 = N6166 & N1415;
  assign N6638 = N6166 & idx_w_i[8];
  assign N6639 = N6168 & N1415;
  assign N6640 = N6168 & idx_w_i[8];
  assign N6641 = N6170 & N1415;
  assign N6642 = N6170 & idx_w_i[8];
  assign N6643 = N6172 & N1415;
  assign N6644 = N6172 & idx_w_i[8];
  assign N6645 = N6174 & N1415;
  assign N6646 = N6174 & idx_w_i[8];
  assign N6647 = N6176 & N1415;
  assign N6648 = N6176 & idx_w_i[8];
  assign N6649 = N6178 & N1415;
  assign N6650 = N6178 & idx_w_i[8];
  assign N6651 = N6180 & N1415;
  assign N6652 = N6180 & idx_w_i[8];
  assign N6653 = N6182 & N1415;
  assign N6654 = N6182 & idx_w_i[8];
  assign N6655 = N6184 & N1415;
  assign N6656 = N6184 & idx_w_i[8];
  assign N6657 = N6186 & N1415;
  assign N6658 = N6186 & idx_w_i[8];
  assign N6659 = N6188 & N1415;
  assign N6660 = N6188 & idx_w_i[8];
  assign N6661 = N6190 & N1415;
  assign N6662 = N6190 & idx_w_i[8];
  assign N6663 = N6192 & N1415;
  assign N6664 = N6192 & idx_w_i[8];
  assign N6665 = N6194 & N1415;
  assign N6666 = N6194 & idx_w_i[8];
  assign N6667 = N6196 & N1415;
  assign N6668 = N6196 & idx_w_i[8];
  assign N6669 = N6198 & N1415;
  assign N6670 = N6198 & idx_w_i[8];
  assign N6671 = N6200 & N1415;
  assign N6672 = N6200 & idx_w_i[8];
  assign N6673 = N6202 & N1415;
  assign N6674 = N6202 & idx_w_i[8];
  assign N6675 = N6204 & N1415;
  assign N6676 = N6204 & idx_w_i[8];
  assign N6677 = N6206 & N1415;
  assign N6678 = N6206 & idx_w_i[8];
  assign N6679 = N6208 & N1415;
  assign N6680 = N6208 & idx_w_i[8];
  assign N6681 = N6210 & N1415;
  assign N6682 = N6210 & idx_w_i[8];
  assign N6683 = N6212 & N1415;
  assign N6684 = N6212 & idx_w_i[8];
  assign N6685 = N6214 & N1415;
  assign N6686 = N6214 & idx_w_i[8];
  assign N6687 = N6216 & N1415;
  assign N6688 = N6216 & idx_w_i[8];
  assign N6689 = N6218 & N1415;
  assign N6690 = N6218 & idx_w_i[8];
  assign N6691 = N6220 & N1415;
  assign N6692 = N6220 & idx_w_i[8];
  assign N6693 = N6222 & N1415;
  assign N6694 = N6222 & idx_w_i[8];
  assign N6695 = N6224 & N1415;
  assign N6696 = N6224 & idx_w_i[8];
  assign N6697 = N6226 & N1415;
  assign N6698 = N6226 & idx_w_i[8];
  assign N6699 = N6228 & N1415;
  assign N6700 = N6228 & idx_w_i[8];
  assign N6701 = N6230 & N1415;
  assign N6702 = N6230 & idx_w_i[8];
  assign N6703 = N5391 & N1415;
  assign N6704 = N5393 & N1415;
  assign N6705 = N5395 & N1415;
  assign N6706 = N5397 & N1415;
  assign N6707 = N5399 & N1415;
  assign N6708 = N5401 & N1415;
  assign N6709 = N5403 & N1415;
  assign N6710 = N5405 & N1415;
  assign N6711 = N5407 & N1415;
  assign N6712 = N5409 & N1415;
  assign N6713 = N5411 & N1415;
  assign N6714 = N5413 & N1415;
  assign N6715 = N5415 & N1415;
  assign N6716 = N5417 & N1415;
  assign N6717 = N5419 & N1415;
  assign N6718 = N5421 & N1415;
  assign N6719 = N6248 & N1415;
  assign N6720 = N6248 & idx_w_i[8];
  assign N6721 = N6250 & N1415;
  assign N6722 = N6250 & idx_w_i[8];
  assign N6723 = N6252 & N1415;
  assign N6724 = N6252 & idx_w_i[8];
  assign N6725 = N6254 & N1415;
  assign N6726 = N6254 & idx_w_i[8];
  assign N6727 = N6256 & N1415;
  assign N6728 = N6256 & idx_w_i[8];
  assign N6729 = N6258 & N1415;
  assign N6730 = N6258 & idx_w_i[8];
  assign N6731 = N6260 & N1415;
  assign N6732 = N6260 & idx_w_i[8];
  assign N6733 = N6262 & N1415;
  assign N6734 = N6262 & idx_w_i[8];
  assign N6735 = N3108 & N1415;
  assign N6736 = N3110 & N1415;
  assign N6737 = N3112 & N1415;
  assign N6738 = N3114 & N1415;
  assign N6739 = N3116 & N1415;
  assign N6740 = N3118 & N1415;
  assign N6741 = N3120 & N1415;
  assign N6742 = N3122 & N1415;
  assign N6743 = N11569 & N1415;
  assign N6744 = N11571 & N1415;
  assign N6745 = N11573 & N1415;
  assign N6746 = N11575 & N1415;
  assign N6747 = N11577 & N1415;
  assign N6748 = N11579 & N1415;
  assign N6749 = N11581 & N1415;
  assign N6750 = N11583 & N1415;
  assign N6751 = N11585 & N1415;
  assign N6752 = N11587 & N1415;
  assign N6753 = N11589 & N1415;
  assign N6754 = N11591 & N1415;
  assign N6755 = N11593 & N1415;
  assign N6756 = N11595 & N1415;
  assign N6757 = N11597 & N1415;
  assign N6758 = N11599 & N1415;
  assign N6760 = N5950 ^ N6759;
  assign N6761 = N5951 & N1060;
  assign N6762 = N5952 & N1060;
  assign N6763 = N5953 & N1060;
  assign N6764 = N5954 & N1060;
  assign N6765 = N5955 & N1060;
  assign N6766 = N5956 & N1060;
  assign N6767 = N5957 & N1060;
  assign N6768 = N5958 & N1060;
  assign N6769 = N2715 & N1060;
  assign N6770 = N2716 & N1060;
  assign N6771 = N2717 & N1060;
  assign N6772 = N2718 & N1060;
  assign N6773 = N2719 & N1060;
  assign N6774 = N2720 & N1060;
  assign N6775 = N2721 & N1060;
  assign N6776 = N2722 & N1060;
  assign N6777 = N11121 & N1060;
  assign N6778 = N11123 & N1060;
  assign N6779 = N11125 & N1060;
  assign N6780 = N11127 & N1060;
  assign N6781 = N11129 & N1060;
  assign N6782 = N11131 & N1060;
  assign N6783 = N11133 & N1060;
  assign N6784 = N11135 & N1060;
  assign N6785 = N6761 & N1093;
  assign N6786 = N6761 & idx_w_i[6];
  assign N6787 = N6762 & N1093;
  assign N6788 = N6762 & idx_w_i[6];
  assign N6789 = N6763 & N1093;
  assign N6790 = N6763 & idx_w_i[6];
  assign N6791 = N6764 & N1093;
  assign N6792 = N6764 & idx_w_i[6];
  assign N6793 = N6765 & N1093;
  assign N6794 = N6765 & idx_w_i[6];
  assign N6795 = N6766 & N1093;
  assign N6796 = N6766 & idx_w_i[6];
  assign N6797 = N6767 & N1093;
  assign N6798 = N6767 & idx_w_i[6];
  assign N6799 = N6768 & N1093;
  assign N6800 = N6768 & idx_w_i[6];
  assign N6801 = N6769 & N1093;
  assign N6802 = N6769 & idx_w_i[6];
  assign N6803 = N6770 & N1093;
  assign N6804 = N6770 & idx_w_i[6];
  assign N6805 = N6771 & N1093;
  assign N6806 = N6771 & idx_w_i[6];
  assign N6807 = N6772 & N1093;
  assign N6808 = N6772 & idx_w_i[6];
  assign N6809 = N6773 & N1093;
  assign N6810 = N6773 & idx_w_i[6];
  assign N6811 = N6774 & N1093;
  assign N6812 = N6774 & idx_w_i[6];
  assign N6813 = N6775 & N1093;
  assign N6814 = N6775 & idx_w_i[6];
  assign N6815 = N6776 & N1093;
  assign N6816 = N6776 & idx_w_i[6];
  assign N6817 = N6777 & N1093;
  assign N6818 = N6777 & idx_w_i[6];
  assign N6819 = N6778 & N1093;
  assign N6820 = N6778 & idx_w_i[6];
  assign N6821 = N6779 & N1093;
  assign N6822 = N6779 & idx_w_i[6];
  assign N6823 = N6780 & N1093;
  assign N6824 = N6780 & idx_w_i[6];
  assign N6825 = N6781 & N1093;
  assign N6826 = N6781 & idx_w_i[6];
  assign N6827 = N6782 & N1093;
  assign N6828 = N6782 & idx_w_i[6];
  assign N6829 = N6783 & N1093;
  assign N6830 = N6783 & idx_w_i[6];
  assign N6831 = N6784 & N1093;
  assign N6832 = N6784 & idx_w_i[6];
  assign N6833 = N3708 & N1093;
  assign N6834 = N3709 & N1093;
  assign N6835 = N3710 & N1093;
  assign N6836 = N3711 & N1093;
  assign N6837 = N3712 & N1093;
  assign N6838 = N3713 & N1093;
  assign N6839 = N3714 & N1093;
  assign N6840 = N3715 & N1093;
  assign N6841 = N5960 & N1093;
  assign N6842 = N5962 & N1093;
  assign N6843 = N5964 & N1093;
  assign N6844 = N5966 & N1093;
  assign N6845 = N5968 & N1093;
  assign N6846 = N5970 & N1093;
  assign N6847 = N5972 & N1093;
  assign N6848 = N5974 & N1093;
  assign N6849 = N2740 & N1093;
  assign N6850 = N2742 & N1093;
  assign N6851 = N2744 & N1093;
  assign N6852 = N2746 & N1093;
  assign N6853 = N2748 & N1093;
  assign N6854 = N2750 & N1093;
  assign N6855 = N2752 & N1093;
  assign N6856 = N2754 & N1093;
  assign N6857 = N11185 & N1093;
  assign N6858 = N11187 & N1093;
  assign N6859 = N11189 & N1093;
  assign N6860 = N11191 & N1093;
  assign N6861 = N11193 & N1093;
  assign N6862 = N11195 & N1093;
  assign N6863 = N11197 & N1093;
  assign N6864 = N11199 & N1093;
  assign N6865 = N11201 & N1093;
  assign N6866 = N11203 & N1093;
  assign N6867 = N11205 & N1093;
  assign N6868 = N11207 & N1093;
  assign N6869 = N11209 & N1093;
  assign N6870 = N11211 & N1093;
  assign N6871 = N11213 & N1093;
  assign N6872 = N11215 & N1093;
  assign N6873 = N6785 & N1190;
  assign N6874 = N6785 & idx_w_i[7];
  assign N6875 = N6787 & N1190;
  assign N6876 = N6787 & idx_w_i[7];
  assign N6877 = N6789 & N1190;
  assign N6878 = N6789 & idx_w_i[7];
  assign N6879 = N6791 & N1190;
  assign N6880 = N6791 & idx_w_i[7];
  assign N6881 = N6793 & N1190;
  assign N6882 = N6793 & idx_w_i[7];
  assign N6883 = N6795 & N1190;
  assign N6884 = N6795 & idx_w_i[7];
  assign N6885 = N6797 & N1190;
  assign N6886 = N6797 & idx_w_i[7];
  assign N6887 = N6799 & N1190;
  assign N6888 = N6799 & idx_w_i[7];
  assign N6889 = N6801 & N1190;
  assign N6890 = N6801 & idx_w_i[7];
  assign N6891 = N6803 & N1190;
  assign N6892 = N6803 & idx_w_i[7];
  assign N6893 = N6805 & N1190;
  assign N6894 = N6805 & idx_w_i[7];
  assign N6895 = N6807 & N1190;
  assign N6896 = N6807 & idx_w_i[7];
  assign N6897 = N6809 & N1190;
  assign N6898 = N6809 & idx_w_i[7];
  assign N6899 = N6811 & N1190;
  assign N6900 = N6811 & idx_w_i[7];
  assign N6901 = N6813 & N1190;
  assign N6902 = N6813 & idx_w_i[7];
  assign N6903 = N6815 & N1190;
  assign N6904 = N6815 & idx_w_i[7];
  assign N6905 = N6817 & N1190;
  assign N6906 = N6817 & idx_w_i[7];
  assign N6907 = N6819 & N1190;
  assign N6908 = N6819 & idx_w_i[7];
  assign N6909 = N6821 & N1190;
  assign N6910 = N6821 & idx_w_i[7];
  assign N6911 = N6823 & N1190;
  assign N6912 = N6823 & idx_w_i[7];
  assign N6913 = N6825 & N1190;
  assign N6914 = N6825 & idx_w_i[7];
  assign N6915 = N6827 & N1190;
  assign N6916 = N6827 & idx_w_i[7];
  assign N6917 = N6829 & N1190;
  assign N6918 = N6829 & idx_w_i[7];
  assign N6919 = N6831 & N1190;
  assign N6920 = N6831 & idx_w_i[7];
  assign N6921 = N6833 & N1190;
  assign N6922 = N6833 & idx_w_i[7];
  assign N6923 = N6834 & N1190;
  assign N6924 = N6834 & idx_w_i[7];
  assign N6925 = N6835 & N1190;
  assign N6926 = N6835 & idx_w_i[7];
  assign N6927 = N6836 & N1190;
  assign N6928 = N6836 & idx_w_i[7];
  assign N6929 = N6837 & N1190;
  assign N6930 = N6837 & idx_w_i[7];
  assign N6931 = N6838 & N1190;
  assign N6932 = N6838 & idx_w_i[7];
  assign N6933 = N6839 & N1190;
  assign N6934 = N6839 & idx_w_i[7];
  assign N6935 = N6840 & N1190;
  assign N6936 = N6840 & idx_w_i[7];
  assign N6937 = N6841 & N1190;
  assign N6938 = N6841 & idx_w_i[7];
  assign N6939 = N6842 & N1190;
  assign N6940 = N6842 & idx_w_i[7];
  assign N6941 = N6843 & N1190;
  assign N6942 = N6843 & idx_w_i[7];
  assign N6943 = N6844 & N1190;
  assign N6944 = N6844 & idx_w_i[7];
  assign N6945 = N6845 & N1190;
  assign N6946 = N6845 & idx_w_i[7];
  assign N6947 = N6846 & N1190;
  assign N6948 = N6846 & idx_w_i[7];
  assign N6949 = N6847 & N1190;
  assign N6950 = N6847 & idx_w_i[7];
  assign N6951 = N6848 & N1190;
  assign N6952 = N6848 & idx_w_i[7];
  assign N6953 = N6849 & N1190;
  assign N6954 = N6849 & idx_w_i[7];
  assign N6955 = N6850 & N1190;
  assign N6956 = N6850 & idx_w_i[7];
  assign N6957 = N6851 & N1190;
  assign N6958 = N6851 & idx_w_i[7];
  assign N6959 = N6852 & N1190;
  assign N6960 = N6852 & idx_w_i[7];
  assign N6961 = N6853 & N1190;
  assign N6962 = N6853 & idx_w_i[7];
  assign N6963 = N6854 & N1190;
  assign N6964 = N6854 & idx_w_i[7];
  assign N6965 = N6855 & N1190;
  assign N6966 = N6855 & idx_w_i[7];
  assign N6967 = N6856 & N1190;
  assign N6968 = N6856 & idx_w_i[7];
  assign N6969 = N6857 & N1190;
  assign N6970 = N6857 & idx_w_i[7];
  assign N6971 = N6858 & N1190;
  assign N6972 = N6858 & idx_w_i[7];
  assign N6973 = N6859 & N1190;
  assign N6974 = N6859 & idx_w_i[7];
  assign N6975 = N6860 & N1190;
  assign N6976 = N6860 & idx_w_i[7];
  assign N6977 = N6861 & N1190;
  assign N6978 = N6861 & idx_w_i[7];
  assign N6979 = N6862 & N1190;
  assign N6980 = N6862 & idx_w_i[7];
  assign N6981 = N6863 & N1190;
  assign N6982 = N6863 & idx_w_i[7];
  assign N6983 = N6864 & N1190;
  assign N6984 = N6864 & idx_w_i[7];
  assign N6985 = N6865 & N1190;
  assign N6986 = N6865 & idx_w_i[7];
  assign N6987 = N6866 & N1190;
  assign N6988 = N6866 & idx_w_i[7];
  assign N6989 = N6867 & N1190;
  assign N6990 = N6867 & idx_w_i[7];
  assign N6991 = N6868 & N1190;
  assign N6992 = N6868 & idx_w_i[7];
  assign N6993 = N6869 & N1190;
  assign N6994 = N6869 & idx_w_i[7];
  assign N6995 = N6870 & N1190;
  assign N6996 = N6870 & idx_w_i[7];
  assign N6997 = N6871 & N1190;
  assign N6998 = N6871 & idx_w_i[7];
  assign N6999 = N6872 & N1190;
  assign N7000 = N6872 & idx_w_i[7];
  assign N7001 = N6786 & N1190;
  assign N7002 = N6786 & idx_w_i[7];
  assign N7003 = N6788 & N1190;
  assign N7004 = N6788 & idx_w_i[7];
  assign N7005 = N6790 & N1190;
  assign N7006 = N6790 & idx_w_i[7];
  assign N7007 = N6792 & N1190;
  assign N7008 = N6792 & idx_w_i[7];
  assign N7009 = N6794 & N1190;
  assign N7010 = N6794 & idx_w_i[7];
  assign N7011 = N6796 & N1190;
  assign N7012 = N6796 & idx_w_i[7];
  assign N7013 = N6798 & N1190;
  assign N7014 = N6798 & idx_w_i[7];
  assign N7015 = N6800 & N1190;
  assign N7016 = N6800 & idx_w_i[7];
  assign N7017 = N6802 & N1190;
  assign N7018 = N6802 & idx_w_i[7];
  assign N7019 = N6804 & N1190;
  assign N7020 = N6804 & idx_w_i[7];
  assign N7021 = N6806 & N1190;
  assign N7022 = N6806 & idx_w_i[7];
  assign N7023 = N6808 & N1190;
  assign N7024 = N6808 & idx_w_i[7];
  assign N7025 = N6810 & N1190;
  assign N7026 = N6810 & idx_w_i[7];
  assign N7027 = N6812 & N1190;
  assign N7028 = N6812 & idx_w_i[7];
  assign N7029 = N6814 & N1190;
  assign N7030 = N6814 & idx_w_i[7];
  assign N7031 = N6816 & N1190;
  assign N7032 = N6816 & idx_w_i[7];
  assign N7033 = N6818 & N1190;
  assign N7034 = N6818 & idx_w_i[7];
  assign N7035 = N6820 & N1190;
  assign N7036 = N6820 & idx_w_i[7];
  assign N7037 = N6822 & N1190;
  assign N7038 = N6822 & idx_w_i[7];
  assign N7039 = N6824 & N1190;
  assign N7040 = N6824 & idx_w_i[7];
  assign N7041 = N6826 & N1190;
  assign N7042 = N6826 & idx_w_i[7];
  assign N7043 = N6828 & N1190;
  assign N7044 = N6828 & idx_w_i[7];
  assign N7045 = N6830 & N1190;
  assign N7046 = N6830 & idx_w_i[7];
  assign N7047 = N6832 & N1190;
  assign N7048 = N6832 & idx_w_i[7];
  assign N7049 = N3765 & N1190;
  assign N7050 = N3767 & N1190;
  assign N7051 = N3769 & N1190;
  assign N7052 = N3771 & N1190;
  assign N7053 = N3773 & N1190;
  assign N7054 = N3775 & N1190;
  assign N7055 = N3777 & N1190;
  assign N7056 = N3779 & N1190;
  assign N7057 = N6032 & N1190;
  assign N7058 = N6034 & N1190;
  assign N7059 = N6036 & N1190;
  assign N7060 = N6038 & N1190;
  assign N7061 = N6040 & N1190;
  assign N7062 = N6042 & N1190;
  assign N7063 = N6044 & N1190;
  assign N7064 = N6046 & N1190;
  assign N7065 = N2860 & N1190;
  assign N7066 = N2862 & N1190;
  assign N7067 = N2864 & N1190;
  assign N7068 = N2866 & N1190;
  assign N7069 = N2868 & N1190;
  assign N7070 = N2870 & N1190;
  assign N7071 = N2872 & N1190;
  assign N7072 = N2874 & N1190;
  assign N7073 = N11313 & N1190;
  assign N7074 = N11315 & N1190;
  assign N7075 = N11317 & N1190;
  assign N7076 = N11319 & N1190;
  assign N7077 = N11321 & N1190;
  assign N7078 = N11323 & N1190;
  assign N7079 = N11325 & N1190;
  assign N7080 = N11327 & N1190;
  assign N7081 = N11329 & N1190;
  assign N7082 = N11331 & N1190;
  assign N7083 = N11333 & N1190;
  assign N7084 = N11335 & N1190;
  assign N7085 = N11337 & N1190;
  assign N7086 = N11339 & N1190;
  assign N7087 = N11341 & N1190;
  assign N7088 = N11343 & N1190;
  assign N7089 = N6873 & N1415;
  assign N7090 = N6873 & idx_w_i[8];
  assign N7091 = N6875 & N1415;
  assign N7092 = N6875 & idx_w_i[8];
  assign N7093 = N6877 & N1415;
  assign N7094 = N6877 & idx_w_i[8];
  assign N7095 = N6879 & N1415;
  assign N7096 = N6879 & idx_w_i[8];
  assign N7097 = N6881 & N1415;
  assign N7098 = N6881 & idx_w_i[8];
  assign N7099 = N6883 & N1415;
  assign N7100 = N6883 & idx_w_i[8];
  assign N7101 = N6885 & N1415;
  assign N7102 = N6885 & idx_w_i[8];
  assign N7103 = N6887 & N1415;
  assign N7104 = N6887 & idx_w_i[8];
  assign N7105 = N6889 & N1415;
  assign N7106 = N6889 & idx_w_i[8];
  assign N7107 = N6891 & N1415;
  assign N7108 = N6891 & idx_w_i[8];
  assign N7109 = N6893 & N1415;
  assign N7110 = N6893 & idx_w_i[8];
  assign N7111 = N6895 & N1415;
  assign N7112 = N6895 & idx_w_i[8];
  assign N7113 = N6897 & N1415;
  assign N7114 = N6897 & idx_w_i[8];
  assign N7115 = N6899 & N1415;
  assign N7116 = N6899 & idx_w_i[8];
  assign N7117 = N6901 & N1415;
  assign N7118 = N6901 & idx_w_i[8];
  assign N7119 = N6903 & N1415;
  assign N7120 = N6903 & idx_w_i[8];
  assign N7121 = N6905 & N1415;
  assign N7122 = N6905 & idx_w_i[8];
  assign N7123 = N6907 & N1415;
  assign N7124 = N6907 & idx_w_i[8];
  assign N7125 = N6909 & N1415;
  assign N7126 = N6909 & idx_w_i[8];
  assign N7127 = N6911 & N1415;
  assign N7128 = N6911 & idx_w_i[8];
  assign N7129 = N6913 & N1415;
  assign N7130 = N6913 & idx_w_i[8];
  assign N7131 = N6915 & N1415;
  assign N7132 = N6915 & idx_w_i[8];
  assign N7133 = N6917 & N1415;
  assign N7134 = N6917 & idx_w_i[8];
  assign N7135 = N6919 & N1415;
  assign N7136 = N6919 & idx_w_i[8];
  assign N7137 = N6921 & N1415;
  assign N7138 = N6921 & idx_w_i[8];
  assign N7139 = N6923 & N1415;
  assign N7140 = N6923 & idx_w_i[8];
  assign N7141 = N6925 & N1415;
  assign N7142 = N6925 & idx_w_i[8];
  assign N7143 = N6927 & N1415;
  assign N7144 = N6927 & idx_w_i[8];
  assign N7145 = N6929 & N1415;
  assign N7146 = N6929 & idx_w_i[8];
  assign N7147 = N6931 & N1415;
  assign N7148 = N6931 & idx_w_i[8];
  assign N7149 = N6933 & N1415;
  assign N7150 = N6933 & idx_w_i[8];
  assign N7151 = N6935 & N1415;
  assign N7152 = N6935 & idx_w_i[8];
  assign N7153 = N6937 & N1415;
  assign N7154 = N6937 & idx_w_i[8];
  assign N7155 = N6939 & N1415;
  assign N7156 = N6939 & idx_w_i[8];
  assign N7157 = N6941 & N1415;
  assign N7158 = N6941 & idx_w_i[8];
  assign N7159 = N6943 & N1415;
  assign N7160 = N6943 & idx_w_i[8];
  assign N7161 = N6945 & N1415;
  assign N7162 = N6945 & idx_w_i[8];
  assign N7163 = N6947 & N1415;
  assign N7164 = N6947 & idx_w_i[8];
  assign N7165 = N6949 & N1415;
  assign N7166 = N6949 & idx_w_i[8];
  assign N7167 = N6951 & N1415;
  assign N7168 = N6951 & idx_w_i[8];
  assign N7169 = N6953 & N1415;
  assign N7170 = N6953 & idx_w_i[8];
  assign N7171 = N6955 & N1415;
  assign N7172 = N6955 & idx_w_i[8];
  assign N7173 = N6957 & N1415;
  assign N7174 = N6957 & idx_w_i[8];
  assign N7175 = N6959 & N1415;
  assign N7176 = N6959 & idx_w_i[8];
  assign N7177 = N6961 & N1415;
  assign N7178 = N6961 & idx_w_i[8];
  assign N7179 = N6963 & N1415;
  assign N7180 = N6963 & idx_w_i[8];
  assign N7181 = N6965 & N1415;
  assign N7182 = N6965 & idx_w_i[8];
  assign N7183 = N6967 & N1415;
  assign N7184 = N6967 & idx_w_i[8];
  assign N7185 = N6969 & N1415;
  assign N7186 = N6969 & idx_w_i[8];
  assign N7187 = N6971 & N1415;
  assign N7188 = N6971 & idx_w_i[8];
  assign N7189 = N6973 & N1415;
  assign N7190 = N6973 & idx_w_i[8];
  assign N7191 = N6975 & N1415;
  assign N7192 = N6975 & idx_w_i[8];
  assign N7193 = N6977 & N1415;
  assign N7194 = N6977 & idx_w_i[8];
  assign N7195 = N6979 & N1415;
  assign N7196 = N6979 & idx_w_i[8];
  assign N7197 = N6981 & N1415;
  assign N7198 = N6981 & idx_w_i[8];
  assign N7199 = N6983 & N1415;
  assign N7200 = N6983 & idx_w_i[8];
  assign N7201 = N6985 & N1415;
  assign N7202 = N6985 & idx_w_i[8];
  assign N7203 = N6987 & N1415;
  assign N7204 = N6987 & idx_w_i[8];
  assign N7205 = N6989 & N1415;
  assign N7206 = N6989 & idx_w_i[8];
  assign N7207 = N6991 & N1415;
  assign N7208 = N6991 & idx_w_i[8];
  assign N7209 = N6993 & N1415;
  assign N7210 = N6993 & idx_w_i[8];
  assign N7211 = N6995 & N1415;
  assign N7212 = N6995 & idx_w_i[8];
  assign N7213 = N6997 & N1415;
  assign N7214 = N6997 & idx_w_i[8];
  assign N7215 = N6999 & N1415;
  assign N7216 = N6999 & idx_w_i[8];
  assign N7217 = N7001 & N1415;
  assign N7218 = N7001 & idx_w_i[8];
  assign N7219 = N7003 & N1415;
  assign N7220 = N7003 & idx_w_i[8];
  assign N7221 = N7005 & N1415;
  assign N7222 = N7005 & idx_w_i[8];
  assign N7223 = N7007 & N1415;
  assign N7224 = N7007 & idx_w_i[8];
  assign N7225 = N7009 & N1415;
  assign N7226 = N7009 & idx_w_i[8];
  assign N7227 = N7011 & N1415;
  assign N7228 = N7011 & idx_w_i[8];
  assign N7229 = N7013 & N1415;
  assign N7230 = N7013 & idx_w_i[8];
  assign N7231 = N7015 & N1415;
  assign N7232 = N7015 & idx_w_i[8];
  assign N7233 = N7017 & N1415;
  assign N7234 = N7017 & idx_w_i[8];
  assign N7235 = N7019 & N1415;
  assign N7236 = N7019 & idx_w_i[8];
  assign N7237 = N7021 & N1415;
  assign N7238 = N7021 & idx_w_i[8];
  assign N7239 = N7023 & N1415;
  assign N7240 = N7023 & idx_w_i[8];
  assign N7241 = N7025 & N1415;
  assign N7242 = N7025 & idx_w_i[8];
  assign N7243 = N7027 & N1415;
  assign N7244 = N7027 & idx_w_i[8];
  assign N7245 = N7029 & N1415;
  assign N7246 = N7029 & idx_w_i[8];
  assign N7247 = N7031 & N1415;
  assign N7248 = N7031 & idx_w_i[8];
  assign N7249 = N7033 & N1415;
  assign N7250 = N7033 & idx_w_i[8];
  assign N7251 = N7035 & N1415;
  assign N7252 = N7035 & idx_w_i[8];
  assign N7253 = N7037 & N1415;
  assign N7254 = N7037 & idx_w_i[8];
  assign N7255 = N7039 & N1415;
  assign N7256 = N7039 & idx_w_i[8];
  assign N7257 = N7041 & N1415;
  assign N7258 = N7041 & idx_w_i[8];
  assign N7259 = N7043 & N1415;
  assign N7260 = N7043 & idx_w_i[8];
  assign N7261 = N7045 & N1415;
  assign N7262 = N7045 & idx_w_i[8];
  assign N7263 = N7047 & N1415;
  assign N7264 = N7047 & idx_w_i[8];
  assign N7265 = N7049 & N1415;
  assign N7266 = N7049 & idx_w_i[8];
  assign N7267 = N7050 & N1415;
  assign N7268 = N7050 & idx_w_i[8];
  assign N7269 = N7051 & N1415;
  assign N7270 = N7051 & idx_w_i[8];
  assign N7271 = N7052 & N1415;
  assign N7272 = N7052 & idx_w_i[8];
  assign N7273 = N7053 & N1415;
  assign N7274 = N7053 & idx_w_i[8];
  assign N7275 = N7054 & N1415;
  assign N7276 = N7054 & idx_w_i[8];
  assign N7277 = N7055 & N1415;
  assign N7278 = N7055 & idx_w_i[8];
  assign N7279 = N7056 & N1415;
  assign N7280 = N7056 & idx_w_i[8];
  assign N7281 = N7057 & N1415;
  assign N7282 = N7057 & idx_w_i[8];
  assign N7283 = N7058 & N1415;
  assign N7284 = N7058 & idx_w_i[8];
  assign N7285 = N7059 & N1415;
  assign N7286 = N7059 & idx_w_i[8];
  assign N7287 = N7060 & N1415;
  assign N7288 = N7060 & idx_w_i[8];
  assign N7289 = N7061 & N1415;
  assign N7290 = N7061 & idx_w_i[8];
  assign N7291 = N7062 & N1415;
  assign N7292 = N7062 & idx_w_i[8];
  assign N7293 = N7063 & N1415;
  assign N7294 = N7063 & idx_w_i[8];
  assign N7295 = N7064 & N1415;
  assign N7296 = N7064 & idx_w_i[8];
  assign N7297 = N7065 & N1415;
  assign N7298 = N7065 & idx_w_i[8];
  assign N7299 = N7066 & N1415;
  assign N7300 = N7066 & idx_w_i[8];
  assign N7301 = N7067 & N1415;
  assign N7302 = N7067 & idx_w_i[8];
  assign N7303 = N7068 & N1415;
  assign N7304 = N7068 & idx_w_i[8];
  assign N7305 = N7069 & N1415;
  assign N7306 = N7069 & idx_w_i[8];
  assign N7307 = N7070 & N1415;
  assign N7308 = N7070 & idx_w_i[8];
  assign N7309 = N7071 & N1415;
  assign N7310 = N7071 & idx_w_i[8];
  assign N7311 = N7072 & N1415;
  assign N7312 = N7072 & idx_w_i[8];
  assign N7313 = N7073 & N1415;
  assign N7314 = N7073 & idx_w_i[8];
  assign N7315 = N7074 & N1415;
  assign N7316 = N7074 & idx_w_i[8];
  assign N7317 = N7075 & N1415;
  assign N7318 = N7075 & idx_w_i[8];
  assign N7319 = N7076 & N1415;
  assign N7320 = N7076 & idx_w_i[8];
  assign N7321 = N7077 & N1415;
  assign N7322 = N7077 & idx_w_i[8];
  assign N7323 = N7078 & N1415;
  assign N7324 = N7078 & idx_w_i[8];
  assign N7325 = N7079 & N1415;
  assign N7326 = N7079 & idx_w_i[8];
  assign N7327 = N7080 & N1415;
  assign N7328 = N7080 & idx_w_i[8];
  assign N7329 = N7081 & N1415;
  assign N7330 = N7081 & idx_w_i[8];
  assign N7331 = N7082 & N1415;
  assign N7332 = N7082 & idx_w_i[8];
  assign N7333 = N7083 & N1415;
  assign N7334 = N7083 & idx_w_i[8];
  assign N7335 = N7084 & N1415;
  assign N7336 = N7084 & idx_w_i[8];
  assign N7337 = N7085 & N1415;
  assign N7338 = N7085 & idx_w_i[8];
  assign N7339 = N7086 & N1415;
  assign N7340 = N7086 & idx_w_i[8];
  assign N7341 = N7087 & N1415;
  assign N7342 = N7087 & idx_w_i[8];
  assign N7343 = N7088 & N1415;
  assign N7344 = N7088 & idx_w_i[8];
  assign N7345 = N6874 & N1415;
  assign N7346 = N6874 & idx_w_i[8];
  assign N7347 = N6876 & N1415;
  assign N7348 = N6876 & idx_w_i[8];
  assign N7349 = N6878 & N1415;
  assign N7350 = N6878 & idx_w_i[8];
  assign N7351 = N6880 & N1415;
  assign N7352 = N6880 & idx_w_i[8];
  assign N7353 = N6882 & N1415;
  assign N7354 = N6882 & idx_w_i[8];
  assign N7355 = N6884 & N1415;
  assign N7356 = N6884 & idx_w_i[8];
  assign N7357 = N6886 & N1415;
  assign N7358 = N6886 & idx_w_i[8];
  assign N7359 = N6888 & N1415;
  assign N7360 = N6888 & idx_w_i[8];
  assign N7361 = N6890 & N1415;
  assign N7362 = N6890 & idx_w_i[8];
  assign N7363 = N6892 & N1415;
  assign N7364 = N6892 & idx_w_i[8];
  assign N7365 = N6894 & N1415;
  assign N7366 = N6894 & idx_w_i[8];
  assign N7367 = N6896 & N1415;
  assign N7368 = N6896 & idx_w_i[8];
  assign N7369 = N6898 & N1415;
  assign N7370 = N6898 & idx_w_i[8];
  assign N7371 = N6900 & N1415;
  assign N7372 = N6900 & idx_w_i[8];
  assign N7373 = N6902 & N1415;
  assign N7374 = N6902 & idx_w_i[8];
  assign N7375 = N6904 & N1415;
  assign N7376 = N6904 & idx_w_i[8];
  assign N7377 = N6906 & N1415;
  assign N7378 = N6906 & idx_w_i[8];
  assign N7379 = N6908 & N1415;
  assign N7380 = N6908 & idx_w_i[8];
  assign N7381 = N6910 & N1415;
  assign N7382 = N6910 & idx_w_i[8];
  assign N7383 = N6912 & N1415;
  assign N7384 = N6912 & idx_w_i[8];
  assign N7385 = N6914 & N1415;
  assign N7386 = N6914 & idx_w_i[8];
  assign N7387 = N6916 & N1415;
  assign N7388 = N6916 & idx_w_i[8];
  assign N7389 = N6918 & N1415;
  assign N7390 = N6918 & idx_w_i[8];
  assign N7391 = N6920 & N1415;
  assign N7392 = N6920 & idx_w_i[8];
  assign N7393 = N6922 & N1415;
  assign N7394 = N6922 & idx_w_i[8];
  assign N7395 = N6924 & N1415;
  assign N7396 = N6924 & idx_w_i[8];
  assign N7397 = N6926 & N1415;
  assign N7398 = N6926 & idx_w_i[8];
  assign N7399 = N6928 & N1415;
  assign N7400 = N6928 & idx_w_i[8];
  assign N7401 = N6930 & N1415;
  assign N7402 = N6930 & idx_w_i[8];
  assign N7403 = N6932 & N1415;
  assign N7404 = N6932 & idx_w_i[8];
  assign N7405 = N6934 & N1415;
  assign N7406 = N6934 & idx_w_i[8];
  assign N7407 = N6936 & N1415;
  assign N7408 = N6936 & idx_w_i[8];
  assign N7409 = N6938 & N1415;
  assign N7410 = N6938 & idx_w_i[8];
  assign N7411 = N6940 & N1415;
  assign N7412 = N6940 & idx_w_i[8];
  assign N7413 = N6942 & N1415;
  assign N7414 = N6942 & idx_w_i[8];
  assign N7415 = N6944 & N1415;
  assign N7416 = N6944 & idx_w_i[8];
  assign N7417 = N6946 & N1415;
  assign N7418 = N6946 & idx_w_i[8];
  assign N7419 = N6948 & N1415;
  assign N7420 = N6948 & idx_w_i[8];
  assign N7421 = N6950 & N1415;
  assign N7422 = N6950 & idx_w_i[8];
  assign N7423 = N6952 & N1415;
  assign N7424 = N6952 & idx_w_i[8];
  assign N7425 = N6954 & N1415;
  assign N7426 = N6954 & idx_w_i[8];
  assign N7427 = N6956 & N1415;
  assign N7428 = N6956 & idx_w_i[8];
  assign N7429 = N6958 & N1415;
  assign N7430 = N6958 & idx_w_i[8];
  assign N7431 = N6960 & N1415;
  assign N7432 = N6960 & idx_w_i[8];
  assign N7433 = N6962 & N1415;
  assign N7434 = N6962 & idx_w_i[8];
  assign N7435 = N6964 & N1415;
  assign N7436 = N6964 & idx_w_i[8];
  assign N7437 = N6966 & N1415;
  assign N7438 = N6966 & idx_w_i[8];
  assign N7439 = N6968 & N1415;
  assign N7440 = N6968 & idx_w_i[8];
  assign N7441 = N6970 & N1415;
  assign N7442 = N6970 & idx_w_i[8];
  assign N7443 = N6972 & N1415;
  assign N7444 = N6972 & idx_w_i[8];
  assign N7445 = N6974 & N1415;
  assign N7446 = N6974 & idx_w_i[8];
  assign N7447 = N6976 & N1415;
  assign N7448 = N6976 & idx_w_i[8];
  assign N7449 = N6978 & N1415;
  assign N7450 = N6978 & idx_w_i[8];
  assign N7451 = N6980 & N1415;
  assign N7452 = N6980 & idx_w_i[8];
  assign N7453 = N6982 & N1415;
  assign N7454 = N6982 & idx_w_i[8];
  assign N7455 = N6984 & N1415;
  assign N7456 = N6984 & idx_w_i[8];
  assign N7457 = N6986 & N1415;
  assign N7458 = N6986 & idx_w_i[8];
  assign N7459 = N6988 & N1415;
  assign N7460 = N6988 & idx_w_i[8];
  assign N7461 = N6990 & N1415;
  assign N7462 = N6990 & idx_w_i[8];
  assign N7463 = N6992 & N1415;
  assign N7464 = N6992 & idx_w_i[8];
  assign N7465 = N6994 & N1415;
  assign N7466 = N6994 & idx_w_i[8];
  assign N7467 = N6996 & N1415;
  assign N7468 = N6996 & idx_w_i[8];
  assign N7469 = N6998 & N1415;
  assign N7470 = N6998 & idx_w_i[8];
  assign N7471 = N7000 & N1415;
  assign N7472 = N7000 & idx_w_i[8];
  assign N7473 = N7002 & N1415;
  assign N7474 = N7002 & idx_w_i[8];
  assign N7475 = N7004 & N1415;
  assign N7476 = N7004 & idx_w_i[8];
  assign N7477 = N7006 & N1415;
  assign N7478 = N7006 & idx_w_i[8];
  assign N7479 = N7008 & N1415;
  assign N7480 = N7008 & idx_w_i[8];
  assign N7481 = N7010 & N1415;
  assign N7482 = N7010 & idx_w_i[8];
  assign N7483 = N7012 & N1415;
  assign N7484 = N7012 & idx_w_i[8];
  assign N7485 = N7014 & N1415;
  assign N7486 = N7014 & idx_w_i[8];
  assign N7487 = N7016 & N1415;
  assign N7488 = N7016 & idx_w_i[8];
  assign N7489 = N7018 & N1415;
  assign N7490 = N7018 & idx_w_i[8];
  assign N7491 = N7020 & N1415;
  assign N7492 = N7020 & idx_w_i[8];
  assign N7493 = N7022 & N1415;
  assign N7494 = N7022 & idx_w_i[8];
  assign N7495 = N7024 & N1415;
  assign N7496 = N7024 & idx_w_i[8];
  assign N7497 = N7026 & N1415;
  assign N7498 = N7026 & idx_w_i[8];
  assign N7499 = N7028 & N1415;
  assign N7500 = N7028 & idx_w_i[8];
  assign N7501 = N7030 & N1415;
  assign N7502 = N7030 & idx_w_i[8];
  assign N7503 = N7032 & N1415;
  assign N7504 = N7032 & idx_w_i[8];
  assign N7505 = N7034 & N1415;
  assign N7506 = N7034 & idx_w_i[8];
  assign N7507 = N7036 & N1415;
  assign N7508 = N7036 & idx_w_i[8];
  assign N7509 = N7038 & N1415;
  assign N7510 = N7038 & idx_w_i[8];
  assign N7511 = N7040 & N1415;
  assign N7512 = N7040 & idx_w_i[8];
  assign N7513 = N7042 & N1415;
  assign N7514 = N7042 & idx_w_i[8];
  assign N7515 = N7044 & N1415;
  assign N7516 = N7044 & idx_w_i[8];
  assign N7517 = N7046 & N1415;
  assign N7518 = N7046 & idx_w_i[8];
  assign N7519 = N7048 & N1415;
  assign N7520 = N7048 & idx_w_i[8];
  assign N7521 = N4005 & N1415;
  assign N7522 = N4007 & N1415;
  assign N7523 = N4009 & N1415;
  assign N7524 = N4011 & N1415;
  assign N7525 = N4013 & N1415;
  assign N7526 = N4015 & N1415;
  assign N7527 = N4017 & N1415;
  assign N7528 = N4019 & N1415;
  assign N7529 = N6248 & N1415;
  assign N7530 = N6250 & N1415;
  assign N7531 = N6252 & N1415;
  assign N7532 = N6254 & N1415;
  assign N7533 = N6256 & N1415;
  assign N7534 = N6258 & N1415;
  assign N7535 = N6260 & N1415;
  assign N7536 = N6262 & N1415;
  assign N7537 = N3108 & N1415;
  assign N7538 = N3110 & N1415;
  assign N7539 = N3112 & N1415;
  assign N7540 = N3114 & N1415;
  assign N7541 = N3116 & N1415;
  assign N7542 = N3118 & N1415;
  assign N7543 = N3120 & N1415;
  assign N7544 = N3122 & N1415;
  assign N7545 = N11569 & N1415;
  assign N7546 = N11571 & N1415;
  assign N7547 = N11573 & N1415;
  assign N7548 = N11575 & N1415;
  assign N7549 = N11577 & N1415;
  assign N7550 = N11579 & N1415;
  assign N7551 = N11581 & N1415;
  assign N7552 = N11583 & N1415;
  assign N7553 = N11585 & N1415;
  assign N7554 = N11587 & N1415;
  assign N7555 = N11589 & N1415;
  assign N7556 = N11591 & N1415;
  assign N7557 = N11593 & N1415;
  assign N7558 = N11595 & N1415;
  assign N7559 = N11597 & N1415;
  assign N7560 = N11599 & N1415;
  assign N7562 = N6761 & N1093;
  assign N7563 = N6762 & N1093;
  assign N7564 = N6763 & N1093;
  assign N7565 = N6764 & N1093;
  assign N7566 = N6765 & N1093;
  assign N7567 = N6766 & N1093;
  assign N7568 = N6767 & N1093;
  assign N7569 = N6768 & N1093;
  assign N7570 = N6769 & N1093;
  assign N7571 = N6770 & N1093;
  assign N7572 = N6771 & N1093;
  assign N7573 = N6772 & N1093;
  assign N7574 = N6773 & N1093;
  assign N7575 = N6774 & N1093;
  assign N7576 = N6775 & N1093;
  assign N7577 = N6776 & N1093;
  assign N7578 = N6777 & N1093;
  assign N7579 = N6778 & N1093;
  assign N7580 = N6779 & N1093;
  assign N7581 = N6780 & N1093;
  assign N7582 = N6781 & N1093;
  assign N7583 = N6782 & N1093;
  assign N7584 = N6783 & N1093;
  assign N7585 = N6784 & N1093;
  assign N7586 = N3708 & N1093;
  assign N7587 = N3709 & N1093;
  assign N7588 = N3710 & N1093;
  assign N7589 = N3711 & N1093;
  assign N7590 = N3712 & N1093;
  assign N7591 = N3713 & N1093;
  assign N7592 = N3714 & N1093;
  assign N7593 = N3715 & N1093;
  assign N7594 = N5960 & N1093;
  assign N7595 = N5962 & N1093;
  assign N7596 = N5964 & N1093;
  assign N7597 = N5966 & N1093;
  assign N7598 = N5968 & N1093;
  assign N7599 = N5970 & N1093;
  assign N7600 = N5972 & N1093;
  assign N7601 = N5974 & N1093;
  assign N7602 = N2740 & N1093;
  assign N7603 = N2742 & N1093;
  assign N7604 = N2744 & N1093;
  assign N7605 = N2746 & N1093;
  assign N7606 = N2748 & N1093;
  assign N7607 = N2750 & N1093;
  assign N7608 = N2752 & N1093;
  assign N7609 = N2754 & N1093;
  assign N7610 = N11185 & N1093;
  assign N7611 = N11187 & N1093;
  assign N7612 = N11189 & N1093;
  assign N7613 = N11191 & N1093;
  assign N7614 = N11193 & N1093;
  assign N7615 = N11195 & N1093;
  assign N7616 = N11197 & N1093;
  assign N7617 = N11199 & N1093;
  assign N7618 = N11201 & N1093;
  assign N7619 = N11203 & N1093;
  assign N7620 = N11205 & N1093;
  assign N7621 = N11207 & N1093;
  assign N7622 = N11209 & N1093;
  assign N7623 = N11211 & N1093;
  assign N7624 = N11213 & N1093;
  assign N7625 = N11215 & N1093;
  assign N7626 = N7562 & N1190;
  assign N7627 = N7562 & idx_w_i[7];
  assign N7628 = N7563 & N1190;
  assign N7629 = N7563 & idx_w_i[7];
  assign N7630 = N7564 & N1190;
  assign N7631 = N7564 & idx_w_i[7];
  assign N7632 = N7565 & N1190;
  assign N7633 = N7565 & idx_w_i[7];
  assign N7634 = N7566 & N1190;
  assign N7635 = N7566 & idx_w_i[7];
  assign N7636 = N7567 & N1190;
  assign N7637 = N7567 & idx_w_i[7];
  assign N7638 = N7568 & N1190;
  assign N7639 = N7568 & idx_w_i[7];
  assign N7640 = N7569 & N1190;
  assign N7641 = N7569 & idx_w_i[7];
  assign N7642 = N7570 & N1190;
  assign N7643 = N7570 & idx_w_i[7];
  assign N7644 = N7571 & N1190;
  assign N7645 = N7571 & idx_w_i[7];
  assign N7646 = N7572 & N1190;
  assign N7647 = N7572 & idx_w_i[7];
  assign N7648 = N7573 & N1190;
  assign N7649 = N7573 & idx_w_i[7];
  assign N7650 = N7574 & N1190;
  assign N7651 = N7574 & idx_w_i[7];
  assign N7652 = N7575 & N1190;
  assign N7653 = N7575 & idx_w_i[7];
  assign N7654 = N7576 & N1190;
  assign N7655 = N7576 & idx_w_i[7];
  assign N7656 = N7577 & N1190;
  assign N7657 = N7577 & idx_w_i[7];
  assign N7658 = N7578 & N1190;
  assign N7659 = N7578 & idx_w_i[7];
  assign N7660 = N7579 & N1190;
  assign N7661 = N7579 & idx_w_i[7];
  assign N7662 = N7580 & N1190;
  assign N7663 = N7580 & idx_w_i[7];
  assign N7664 = N7581 & N1190;
  assign N7665 = N7581 & idx_w_i[7];
  assign N7666 = N7582 & N1190;
  assign N7667 = N7582 & idx_w_i[7];
  assign N7668 = N7583 & N1190;
  assign N7669 = N7583 & idx_w_i[7];
  assign N7670 = N7584 & N1190;
  assign N7671 = N7584 & idx_w_i[7];
  assign N7672 = N7585 & N1190;
  assign N7673 = N7585 & idx_w_i[7];
  assign N7674 = N7586 & N1190;
  assign N7675 = N7586 & idx_w_i[7];
  assign N7676 = N7587 & N1190;
  assign N7677 = N7587 & idx_w_i[7];
  assign N7678 = N7588 & N1190;
  assign N7679 = N7588 & idx_w_i[7];
  assign N7680 = N7589 & N1190;
  assign N7681 = N7589 & idx_w_i[7];
  assign N7682 = N7590 & N1190;
  assign N7683 = N7590 & idx_w_i[7];
  assign N7684 = N7591 & N1190;
  assign N7685 = N7591 & idx_w_i[7];
  assign N7686 = N7592 & N1190;
  assign N7687 = N7592 & idx_w_i[7];
  assign N7688 = N7593 & N1190;
  assign N7689 = N7593 & idx_w_i[7];
  assign N7690 = N7594 & N1190;
  assign N7691 = N7594 & idx_w_i[7];
  assign N7692 = N7595 & N1190;
  assign N7693 = N7595 & idx_w_i[7];
  assign N7694 = N7596 & N1190;
  assign N7695 = N7596 & idx_w_i[7];
  assign N7696 = N7597 & N1190;
  assign N7697 = N7597 & idx_w_i[7];
  assign N7698 = N7598 & N1190;
  assign N7699 = N7598 & idx_w_i[7];
  assign N7700 = N7599 & N1190;
  assign N7701 = N7599 & idx_w_i[7];
  assign N7702 = N7600 & N1190;
  assign N7703 = N7600 & idx_w_i[7];
  assign N7704 = N7601 & N1190;
  assign N7705 = N7601 & idx_w_i[7];
  assign N7706 = N7602 & N1190;
  assign N7707 = N7602 & idx_w_i[7];
  assign N7708 = N7603 & N1190;
  assign N7709 = N7603 & idx_w_i[7];
  assign N7710 = N7604 & N1190;
  assign N7711 = N7604 & idx_w_i[7];
  assign N7712 = N7605 & N1190;
  assign N7713 = N7605 & idx_w_i[7];
  assign N7714 = N7606 & N1190;
  assign N7715 = N7606 & idx_w_i[7];
  assign N7716 = N7607 & N1190;
  assign N7717 = N7607 & idx_w_i[7];
  assign N7718 = N7608 & N1190;
  assign N7719 = N7608 & idx_w_i[7];
  assign N7720 = N7609 & N1190;
  assign N7721 = N7609 & idx_w_i[7];
  assign N7722 = N7610 & N1190;
  assign N7723 = N7610 & idx_w_i[7];
  assign N7724 = N7611 & N1190;
  assign N7725 = N7611 & idx_w_i[7];
  assign N7726 = N7612 & N1190;
  assign N7727 = N7612 & idx_w_i[7];
  assign N7728 = N7613 & N1190;
  assign N7729 = N7613 & idx_w_i[7];
  assign N7730 = N7614 & N1190;
  assign N7731 = N7614 & idx_w_i[7];
  assign N7732 = N7615 & N1190;
  assign N7733 = N7615 & idx_w_i[7];
  assign N7734 = N7616 & N1190;
  assign N7735 = N7616 & idx_w_i[7];
  assign N7736 = N7617 & N1190;
  assign N7737 = N7617 & idx_w_i[7];
  assign N7738 = N7618 & N1190;
  assign N7739 = N7618 & idx_w_i[7];
  assign N7740 = N7619 & N1190;
  assign N7741 = N7619 & idx_w_i[7];
  assign N7742 = N7620 & N1190;
  assign N7743 = N7620 & idx_w_i[7];
  assign N7744 = N7621 & N1190;
  assign N7745 = N7621 & idx_w_i[7];
  assign N7746 = N7622 & N1190;
  assign N7747 = N7622 & idx_w_i[7];
  assign N7748 = N7623 & N1190;
  assign N7749 = N7623 & idx_w_i[7];
  assign N7750 = N7624 & N1190;
  assign N7751 = N7624 & idx_w_i[7];
  assign N7752 = N7625 & N1190;
  assign N7753 = N7625 & idx_w_i[7];
  assign N7754 = N6786 & N1190;
  assign N7755 = N6788 & N1190;
  assign N7756 = N6790 & N1190;
  assign N7757 = N6792 & N1190;
  assign N7758 = N6794 & N1190;
  assign N7759 = N6796 & N1190;
  assign N7760 = N6798 & N1190;
  assign N7761 = N6800 & N1190;
  assign N7762 = N6802 & N1190;
  assign N7763 = N6804 & N1190;
  assign N7764 = N6806 & N1190;
  assign N7765 = N6808 & N1190;
  assign N7766 = N6810 & N1190;
  assign N7767 = N6812 & N1190;
  assign N7768 = N6814 & N1190;
  assign N7769 = N6816 & N1190;
  assign N7770 = N6818 & N1190;
  assign N7771 = N6820 & N1190;
  assign N7772 = N6822 & N1190;
  assign N7773 = N6824 & N1190;
  assign N7774 = N6826 & N1190;
  assign N7775 = N6828 & N1190;
  assign N7776 = N6830 & N1190;
  assign N7777 = N6832 & N1190;
  assign N7778 = N3765 & N1190;
  assign N7779 = N3767 & N1190;
  assign N7780 = N3769 & N1190;
  assign N7781 = N3771 & N1190;
  assign N7782 = N3773 & N1190;
  assign N7783 = N3775 & N1190;
  assign N7784 = N3777 & N1190;
  assign N7785 = N3779 & N1190;
  assign N7786 = N6032 & N1190;
  assign N7787 = N6034 & N1190;
  assign N7788 = N6036 & N1190;
  assign N7789 = N6038 & N1190;
  assign N7790 = N6040 & N1190;
  assign N7791 = N6042 & N1190;
  assign N7792 = N6044 & N1190;
  assign N7793 = N6046 & N1190;
  assign N7794 = N2860 & N1190;
  assign N7795 = N2862 & N1190;
  assign N7796 = N2864 & N1190;
  assign N7797 = N2866 & N1190;
  assign N7798 = N2868 & N1190;
  assign N7799 = N2870 & N1190;
  assign N7800 = N2872 & N1190;
  assign N7801 = N2874 & N1190;
  assign N7802 = N11313 & N1190;
  assign N7803 = N11315 & N1190;
  assign N7804 = N11317 & N1190;
  assign N7805 = N11319 & N1190;
  assign N7806 = N11321 & N1190;
  assign N7807 = N11323 & N1190;
  assign N7808 = N11325 & N1190;
  assign N7809 = N11327 & N1190;
  assign N7810 = N11329 & N1190;
  assign N7811 = N11331 & N1190;
  assign N7812 = N11333 & N1190;
  assign N7813 = N11335 & N1190;
  assign N7814 = N11337 & N1190;
  assign N7815 = N11339 & N1190;
  assign N7816 = N11341 & N1190;
  assign N7817 = N11343 & N1190;
  assign N7818 = N7626 & N1415;
  assign N7819 = N7626 & idx_w_i[8];
  assign N7820 = N7628 & N1415;
  assign N7821 = N7628 & idx_w_i[8];
  assign N7822 = N7630 & N1415;
  assign N7823 = N7630 & idx_w_i[8];
  assign N7824 = N7632 & N1415;
  assign N7825 = N7632 & idx_w_i[8];
  assign N7826 = N7634 & N1415;
  assign N7827 = N7634 & idx_w_i[8];
  assign N7828 = N7636 & N1415;
  assign N7829 = N7636 & idx_w_i[8];
  assign N7830 = N7638 & N1415;
  assign N7831 = N7638 & idx_w_i[8];
  assign N7832 = N7640 & N1415;
  assign N7833 = N7640 & idx_w_i[8];
  assign N7834 = N7642 & N1415;
  assign N7835 = N7642 & idx_w_i[8];
  assign N7836 = N7644 & N1415;
  assign N7837 = N7644 & idx_w_i[8];
  assign N7838 = N7646 & N1415;
  assign N7839 = N7646 & idx_w_i[8];
  assign N7840 = N7648 & N1415;
  assign N7841 = N7648 & idx_w_i[8];
  assign N7842 = N7650 & N1415;
  assign N7843 = N7650 & idx_w_i[8];
  assign N7844 = N7652 & N1415;
  assign N7845 = N7652 & idx_w_i[8];
  assign N7846 = N7654 & N1415;
  assign N7847 = N7654 & idx_w_i[8];
  assign N7848 = N7656 & N1415;
  assign N7849 = N7656 & idx_w_i[8];
  assign N7850 = N7658 & N1415;
  assign N7851 = N7658 & idx_w_i[8];
  assign N7852 = N7660 & N1415;
  assign N7853 = N7660 & idx_w_i[8];
  assign N7854 = N7662 & N1415;
  assign N7855 = N7662 & idx_w_i[8];
  assign N7856 = N7664 & N1415;
  assign N7857 = N7664 & idx_w_i[8];
  assign N7858 = N7666 & N1415;
  assign N7859 = N7666 & idx_w_i[8];
  assign N7860 = N7668 & N1415;
  assign N7861 = N7668 & idx_w_i[8];
  assign N7862 = N7670 & N1415;
  assign N7863 = N7670 & idx_w_i[8];
  assign N7864 = N7672 & N1415;
  assign N7865 = N7672 & idx_w_i[8];
  assign N7866 = N7674 & N1415;
  assign N7867 = N7674 & idx_w_i[8];
  assign N7868 = N7676 & N1415;
  assign N7869 = N7676 & idx_w_i[8];
  assign N7870 = N7678 & N1415;
  assign N7871 = N7678 & idx_w_i[8];
  assign N7872 = N7680 & N1415;
  assign N7873 = N7680 & idx_w_i[8];
  assign N7874 = N7682 & N1415;
  assign N7875 = N7682 & idx_w_i[8];
  assign N7876 = N7684 & N1415;
  assign N7877 = N7684 & idx_w_i[8];
  assign N7878 = N7686 & N1415;
  assign N7879 = N7686 & idx_w_i[8];
  assign N7880 = N7688 & N1415;
  assign N7881 = N7688 & idx_w_i[8];
  assign N7882 = N7690 & N1415;
  assign N7883 = N7690 & idx_w_i[8];
  assign N7884 = N7692 & N1415;
  assign N7885 = N7692 & idx_w_i[8];
  assign N7886 = N7694 & N1415;
  assign N7887 = N7694 & idx_w_i[8];
  assign N7888 = N7696 & N1415;
  assign N7889 = N7696 & idx_w_i[8];
  assign N7890 = N7698 & N1415;
  assign N7891 = N7698 & idx_w_i[8];
  assign N7892 = N7700 & N1415;
  assign N7893 = N7700 & idx_w_i[8];
  assign N7894 = N7702 & N1415;
  assign N7895 = N7702 & idx_w_i[8];
  assign N7896 = N7704 & N1415;
  assign N7897 = N7704 & idx_w_i[8];
  assign N7898 = N7706 & N1415;
  assign N7899 = N7706 & idx_w_i[8];
  assign N7900 = N7708 & N1415;
  assign N7901 = N7708 & idx_w_i[8];
  assign N7902 = N7710 & N1415;
  assign N7903 = N7710 & idx_w_i[8];
  assign N7904 = N7712 & N1415;
  assign N7905 = N7712 & idx_w_i[8];
  assign N7906 = N7714 & N1415;
  assign N7907 = N7714 & idx_w_i[8];
  assign N7908 = N7716 & N1415;
  assign N7909 = N7716 & idx_w_i[8];
  assign N7910 = N7718 & N1415;
  assign N7911 = N7718 & idx_w_i[8];
  assign N7912 = N7720 & N1415;
  assign N7913 = N7720 & idx_w_i[8];
  assign N7914 = N7722 & N1415;
  assign N7915 = N7722 & idx_w_i[8];
  assign N7916 = N7724 & N1415;
  assign N7917 = N7724 & idx_w_i[8];
  assign N7918 = N7726 & N1415;
  assign N7919 = N7726 & idx_w_i[8];
  assign N7920 = N7728 & N1415;
  assign N7921 = N7728 & idx_w_i[8];
  assign N7922 = N7730 & N1415;
  assign N7923 = N7730 & idx_w_i[8];
  assign N7924 = N7732 & N1415;
  assign N7925 = N7732 & idx_w_i[8];
  assign N7926 = N7734 & N1415;
  assign N7927 = N7734 & idx_w_i[8];
  assign N7928 = N7736 & N1415;
  assign N7929 = N7736 & idx_w_i[8];
  assign N7930 = N7738 & N1415;
  assign N7931 = N7738 & idx_w_i[8];
  assign N7932 = N7740 & N1415;
  assign N7933 = N7740 & idx_w_i[8];
  assign N7934 = N7742 & N1415;
  assign N7935 = N7742 & idx_w_i[8];
  assign N7936 = N7744 & N1415;
  assign N7937 = N7744 & idx_w_i[8];
  assign N7938 = N7746 & N1415;
  assign N7939 = N7746 & idx_w_i[8];
  assign N7940 = N7748 & N1415;
  assign N7941 = N7748 & idx_w_i[8];
  assign N7942 = N7750 & N1415;
  assign N7943 = N7750 & idx_w_i[8];
  assign N7944 = N7752 & N1415;
  assign N7945 = N7752 & idx_w_i[8];
  assign N7946 = N7754 & N1415;
  assign N7947 = N7754 & idx_w_i[8];
  assign N7948 = N7755 & N1415;
  assign N7949 = N7755 & idx_w_i[8];
  assign N7950 = N7756 & N1415;
  assign N7951 = N7756 & idx_w_i[8];
  assign N7952 = N7757 & N1415;
  assign N7953 = N7757 & idx_w_i[8];
  assign N7954 = N7758 & N1415;
  assign N7955 = N7758 & idx_w_i[8];
  assign N7956 = N7759 & N1415;
  assign N7957 = N7759 & idx_w_i[8];
  assign N7958 = N7760 & N1415;
  assign N7959 = N7760 & idx_w_i[8];
  assign N7960 = N7761 & N1415;
  assign N7961 = N7761 & idx_w_i[8];
  assign N7962 = N7762 & N1415;
  assign N7963 = N7762 & idx_w_i[8];
  assign N7964 = N7763 & N1415;
  assign N7965 = N7763 & idx_w_i[8];
  assign N7966 = N7764 & N1415;
  assign N7967 = N7764 & idx_w_i[8];
  assign N7968 = N7765 & N1415;
  assign N7969 = N7765 & idx_w_i[8];
  assign N7970 = N7766 & N1415;
  assign N7971 = N7766 & idx_w_i[8];
  assign N7972 = N7767 & N1415;
  assign N7973 = N7767 & idx_w_i[8];
  assign N7974 = N7768 & N1415;
  assign N7975 = N7768 & idx_w_i[8];
  assign N7976 = N7769 & N1415;
  assign N7977 = N7769 & idx_w_i[8];
  assign N7978 = N7770 & N1415;
  assign N7979 = N7770 & idx_w_i[8];
  assign N7980 = N7771 & N1415;
  assign N7981 = N7771 & idx_w_i[8];
  assign N7982 = N7772 & N1415;
  assign N7983 = N7772 & idx_w_i[8];
  assign N7984 = N7773 & N1415;
  assign N7985 = N7773 & idx_w_i[8];
  assign N7986 = N7774 & N1415;
  assign N7987 = N7774 & idx_w_i[8];
  assign N7988 = N7775 & N1415;
  assign N7989 = N7775 & idx_w_i[8];
  assign N7990 = N7776 & N1415;
  assign N7991 = N7776 & idx_w_i[8];
  assign N7992 = N7777 & N1415;
  assign N7993 = N7777 & idx_w_i[8];
  assign N7994 = N7778 & N1415;
  assign N7995 = N7778 & idx_w_i[8];
  assign N7996 = N7779 & N1415;
  assign N7997 = N7779 & idx_w_i[8];
  assign N7998 = N7780 & N1415;
  assign N7999 = N7780 & idx_w_i[8];
  assign N8000 = N7781 & N1415;
  assign N8001 = N7781 & idx_w_i[8];
  assign N8002 = N7782 & N1415;
  assign N8003 = N7782 & idx_w_i[8];
  assign N8004 = N7783 & N1415;
  assign N8005 = N7783 & idx_w_i[8];
  assign N8006 = N7784 & N1415;
  assign N8007 = N7784 & idx_w_i[8];
  assign N8008 = N7785 & N1415;
  assign N8009 = N7785 & idx_w_i[8];
  assign N8010 = N7786 & N1415;
  assign N8011 = N7786 & idx_w_i[8];
  assign N8012 = N7787 & N1415;
  assign N8013 = N7787 & idx_w_i[8];
  assign N8014 = N7788 & N1415;
  assign N8015 = N7788 & idx_w_i[8];
  assign N8016 = N7789 & N1415;
  assign N8017 = N7789 & idx_w_i[8];
  assign N8018 = N7790 & N1415;
  assign N8019 = N7790 & idx_w_i[8];
  assign N8020 = N7791 & N1415;
  assign N8021 = N7791 & idx_w_i[8];
  assign N8022 = N7792 & N1415;
  assign N8023 = N7792 & idx_w_i[8];
  assign N8024 = N7793 & N1415;
  assign N8025 = N7793 & idx_w_i[8];
  assign N8026 = N7794 & N1415;
  assign N8027 = N7794 & idx_w_i[8];
  assign N8028 = N7795 & N1415;
  assign N8029 = N7795 & idx_w_i[8];
  assign N8030 = N7796 & N1415;
  assign N8031 = N7796 & idx_w_i[8];
  assign N8032 = N7797 & N1415;
  assign N8033 = N7797 & idx_w_i[8];
  assign N8034 = N7798 & N1415;
  assign N8035 = N7798 & idx_w_i[8];
  assign N8036 = N7799 & N1415;
  assign N8037 = N7799 & idx_w_i[8];
  assign N8038 = N7800 & N1415;
  assign N8039 = N7800 & idx_w_i[8];
  assign N8040 = N7801 & N1415;
  assign N8041 = N7801 & idx_w_i[8];
  assign N8042 = N7802 & N1415;
  assign N8043 = N7802 & idx_w_i[8];
  assign N8044 = N7803 & N1415;
  assign N8045 = N7803 & idx_w_i[8];
  assign N8046 = N7804 & N1415;
  assign N8047 = N7804 & idx_w_i[8];
  assign N8048 = N7805 & N1415;
  assign N8049 = N7805 & idx_w_i[8];
  assign N8050 = N7806 & N1415;
  assign N8051 = N7806 & idx_w_i[8];
  assign N8052 = N7807 & N1415;
  assign N8053 = N7807 & idx_w_i[8];
  assign N8054 = N7808 & N1415;
  assign N8055 = N7808 & idx_w_i[8];
  assign N8056 = N7809 & N1415;
  assign N8057 = N7809 & idx_w_i[8];
  assign N8058 = N7810 & N1415;
  assign N8059 = N7810 & idx_w_i[8];
  assign N8060 = N7811 & N1415;
  assign N8061 = N7811 & idx_w_i[8];
  assign N8062 = N7812 & N1415;
  assign N8063 = N7812 & idx_w_i[8];
  assign N8064 = N7813 & N1415;
  assign N8065 = N7813 & idx_w_i[8];
  assign N8066 = N7814 & N1415;
  assign N8067 = N7814 & idx_w_i[8];
  assign N8068 = N7815 & N1415;
  assign N8069 = N7815 & idx_w_i[8];
  assign N8070 = N7816 & N1415;
  assign N8071 = N7816 & idx_w_i[8];
  assign N8072 = N7817 & N1415;
  assign N8073 = N7817 & idx_w_i[8];
  assign N8074 = N7627 & N1415;
  assign N8075 = N7627 & idx_w_i[8];
  assign N8076 = N7629 & N1415;
  assign N8077 = N7629 & idx_w_i[8];
  assign N8078 = N7631 & N1415;
  assign N8079 = N7631 & idx_w_i[8];
  assign N8080 = N7633 & N1415;
  assign N8081 = N7633 & idx_w_i[8];
  assign N8082 = N7635 & N1415;
  assign N8083 = N7635 & idx_w_i[8];
  assign N8084 = N7637 & N1415;
  assign N8085 = N7637 & idx_w_i[8];
  assign N8086 = N7639 & N1415;
  assign N8087 = N7639 & idx_w_i[8];
  assign N8088 = N7641 & N1415;
  assign N8089 = N7641 & idx_w_i[8];
  assign N8090 = N7643 & N1415;
  assign N8091 = N7643 & idx_w_i[8];
  assign N8092 = N7645 & N1415;
  assign N8093 = N7645 & idx_w_i[8];
  assign N8094 = N7647 & N1415;
  assign N8095 = N7647 & idx_w_i[8];
  assign N8096 = N7649 & N1415;
  assign N8097 = N7649 & idx_w_i[8];
  assign N8098 = N7651 & N1415;
  assign N8099 = N7651 & idx_w_i[8];
  assign N8100 = N7653 & N1415;
  assign N8101 = N7653 & idx_w_i[8];
  assign N8102 = N7655 & N1415;
  assign N8103 = N7655 & idx_w_i[8];
  assign N8104 = N7657 & N1415;
  assign N8105 = N7657 & idx_w_i[8];
  assign N8106 = N7659 & N1415;
  assign N8107 = N7659 & idx_w_i[8];
  assign N8108 = N7661 & N1415;
  assign N8109 = N7661 & idx_w_i[8];
  assign N8110 = N7663 & N1415;
  assign N8111 = N7663 & idx_w_i[8];
  assign N8112 = N7665 & N1415;
  assign N8113 = N7665 & idx_w_i[8];
  assign N8114 = N7667 & N1415;
  assign N8115 = N7667 & idx_w_i[8];
  assign N8116 = N7669 & N1415;
  assign N8117 = N7669 & idx_w_i[8];
  assign N8118 = N7671 & N1415;
  assign N8119 = N7671 & idx_w_i[8];
  assign N8120 = N7673 & N1415;
  assign N8121 = N7673 & idx_w_i[8];
  assign N8122 = N7675 & N1415;
  assign N8123 = N7675 & idx_w_i[8];
  assign N8124 = N7677 & N1415;
  assign N8125 = N7677 & idx_w_i[8];
  assign N8126 = N7679 & N1415;
  assign N8127 = N7679 & idx_w_i[8];
  assign N8128 = N7681 & N1415;
  assign N8129 = N7681 & idx_w_i[8];
  assign N8130 = N7683 & N1415;
  assign N8131 = N7683 & idx_w_i[8];
  assign N8132 = N7685 & N1415;
  assign N8133 = N7685 & idx_w_i[8];
  assign N8134 = N7687 & N1415;
  assign N8135 = N7687 & idx_w_i[8];
  assign N8136 = N7689 & N1415;
  assign N8137 = N7689 & idx_w_i[8];
  assign N8138 = N7691 & N1415;
  assign N8139 = N7691 & idx_w_i[8];
  assign N8140 = N7693 & N1415;
  assign N8141 = N7693 & idx_w_i[8];
  assign N8142 = N7695 & N1415;
  assign N8143 = N7695 & idx_w_i[8];
  assign N8144 = N7697 & N1415;
  assign N8145 = N7697 & idx_w_i[8];
  assign N8146 = N7699 & N1415;
  assign N8147 = N7699 & idx_w_i[8];
  assign N8148 = N7701 & N1415;
  assign N8149 = N7701 & idx_w_i[8];
  assign N8150 = N7703 & N1415;
  assign N8151 = N7703 & idx_w_i[8];
  assign N8152 = N7705 & N1415;
  assign N8153 = N7705 & idx_w_i[8];
  assign N8154 = N7707 & N1415;
  assign N8155 = N7707 & idx_w_i[8];
  assign N8156 = N7709 & N1415;
  assign N8157 = N7709 & idx_w_i[8];
  assign N8158 = N7711 & N1415;
  assign N8159 = N7711 & idx_w_i[8];
  assign N8160 = N7713 & N1415;
  assign N8161 = N7713 & idx_w_i[8];
  assign N8162 = N7715 & N1415;
  assign N8163 = N7715 & idx_w_i[8];
  assign N8164 = N7717 & N1415;
  assign N8165 = N7717 & idx_w_i[8];
  assign N8166 = N7719 & N1415;
  assign N8167 = N7719 & idx_w_i[8];
  assign N8168 = N7721 & N1415;
  assign N8169 = N7721 & idx_w_i[8];
  assign N8170 = N7723 & N1415;
  assign N8171 = N7723 & idx_w_i[8];
  assign N8172 = N7725 & N1415;
  assign N8173 = N7725 & idx_w_i[8];
  assign N8174 = N7727 & N1415;
  assign N8175 = N7727 & idx_w_i[8];
  assign N8176 = N7729 & N1415;
  assign N8177 = N7729 & idx_w_i[8];
  assign N8178 = N7731 & N1415;
  assign N8179 = N7731 & idx_w_i[8];
  assign N8180 = N7733 & N1415;
  assign N8181 = N7733 & idx_w_i[8];
  assign N8182 = N7735 & N1415;
  assign N8183 = N7735 & idx_w_i[8];
  assign N8184 = N7737 & N1415;
  assign N8185 = N7737 & idx_w_i[8];
  assign N8186 = N7739 & N1415;
  assign N8187 = N7739 & idx_w_i[8];
  assign N8188 = N7741 & N1415;
  assign N8189 = N7741 & idx_w_i[8];
  assign N8190 = N7743 & N1415;
  assign N8191 = N7743 & idx_w_i[8];
  assign N8192 = N7745 & N1415;
  assign N8193 = N7745 & idx_w_i[8];
  assign N8194 = N7747 & N1415;
  assign N8195 = N7747 & idx_w_i[8];
  assign N8196 = N7749 & N1415;
  assign N8197 = N7749 & idx_w_i[8];
  assign N8198 = N7751 & N1415;
  assign N8199 = N7751 & idx_w_i[8];
  assign N8200 = N7753 & N1415;
  assign N8201 = N7753 & idx_w_i[8];
  assign N8202 = N7002 & N1415;
  assign N8203 = N7004 & N1415;
  assign N8204 = N7006 & N1415;
  assign N8205 = N7008 & N1415;
  assign N8206 = N7010 & N1415;
  assign N8207 = N7012 & N1415;
  assign N8208 = N7014 & N1415;
  assign N8209 = N7016 & N1415;
  assign N8210 = N7018 & N1415;
  assign N8211 = N7020 & N1415;
  assign N8212 = N7022 & N1415;
  assign N8213 = N7024 & N1415;
  assign N8214 = N7026 & N1415;
  assign N8215 = N7028 & N1415;
  assign N8216 = N7030 & N1415;
  assign N8217 = N7032 & N1415;
  assign N8218 = N7034 & N1415;
  assign N8219 = N7036 & N1415;
  assign N8220 = N7038 & N1415;
  assign N8221 = N7040 & N1415;
  assign N8222 = N7042 & N1415;
  assign N8223 = N7044 & N1415;
  assign N8224 = N7046 & N1415;
  assign N8225 = N7048 & N1415;
  assign N8226 = N4005 & N1415;
  assign N8227 = N4007 & N1415;
  assign N8228 = N4009 & N1415;
  assign N8229 = N4011 & N1415;
  assign N8230 = N4013 & N1415;
  assign N8231 = N4015 & N1415;
  assign N8232 = N4017 & N1415;
  assign N8233 = N4019 & N1415;
  assign N8234 = N6248 & N1415;
  assign N8235 = N6250 & N1415;
  assign N8236 = N6252 & N1415;
  assign N8237 = N6254 & N1415;
  assign N8238 = N6256 & N1415;
  assign N8239 = N6258 & N1415;
  assign N8240 = N6260 & N1415;
  assign N8241 = N6262 & N1415;
  assign N8242 = N3108 & N1415;
  assign N8243 = N3110 & N1415;
  assign N8244 = N3112 & N1415;
  assign N8245 = N3114 & N1415;
  assign N8246 = N3116 & N1415;
  assign N8247 = N3118 & N1415;
  assign N8248 = N3120 & N1415;
  assign N8249 = N3122 & N1415;
  assign N8250 = N11569 & N1415;
  assign N8251 = N11571 & N1415;
  assign N8252 = N11573 & N1415;
  assign N8253 = N11575 & N1415;
  assign N8254 = N11577 & N1415;
  assign N8255 = N11579 & N1415;
  assign N8256 = N11581 & N1415;
  assign N8257 = N11583 & N1415;
  assign N8258 = N11585 & N1415;
  assign N8259 = N11587 & N1415;
  assign N8260 = N11589 & N1415;
  assign N8261 = N11591 & N1415;
  assign N8262 = N11593 & N1415;
  assign N8263 = N11595 & N1415;
  assign N8264 = N11597 & N1415;
  assign N8265 = N11599 & N1415;
  assign N8267 = N7561 ^ N8266;
  assign N8268 = N5951 & N1060;
  assign N8269 = N5952 & N1060;
  assign N8270 = N5953 & N1060;
  assign N8271 = N5954 & N1060;
  assign N8272 = N5955 & N1060;
  assign N8273 = N5956 & N1060;
  assign N8274 = N5957 & N1060;
  assign N8275 = N5958 & N1060;
  assign N8276 = N11121 & N1060;
  assign N8277 = N11123 & N1060;
  assign N8278 = N11125 & N1060;
  assign N8279 = N11127 & N1060;
  assign N8280 = N11129 & N1060;
  assign N8281 = N11131 & N1060;
  assign N8282 = N11133 & N1060;
  assign N8283 = N11135 & N1060;
  assign N8284 = N8268 & N1093;
  assign N8285 = N8268 & idx_w_i[6];
  assign N8286 = N8269 & N1093;
  assign N8287 = N8269 & idx_w_i[6];
  assign N8288 = N8270 & N1093;
  assign N8289 = N8270 & idx_w_i[6];
  assign N8290 = N8271 & N1093;
  assign N8291 = N8271 & idx_w_i[6];
  assign N8292 = N8272 & N1093;
  assign N8293 = N8272 & idx_w_i[6];
  assign N8294 = N8273 & N1093;
  assign N8295 = N8273 & idx_w_i[6];
  assign N8296 = N8274 & N1093;
  assign N8297 = N8274 & idx_w_i[6];
  assign N8298 = N8275 & N1093;
  assign N8299 = N8275 & idx_w_i[6];
  assign N8300 = N2739 & N1093;
  assign N8301 = N2741 & N1093;
  assign N8302 = N2743 & N1093;
  assign N8303 = N2745 & N1093;
  assign N8304 = N2747 & N1093;
  assign N8305 = N2749 & N1093;
  assign N8306 = N2751 & N1093;
  assign N8307 = N2753 & N1093;
  assign N8308 = N8276 & N1093;
  assign N8309 = N8276 & idx_w_i[6];
  assign N8310 = N8277 & N1093;
  assign N8311 = N8277 & idx_w_i[6];
  assign N8312 = N8278 & N1093;
  assign N8313 = N8278 & idx_w_i[6];
  assign N8314 = N8279 & N1093;
  assign N8315 = N8279 & idx_w_i[6];
  assign N8316 = N8280 & N1093;
  assign N8317 = N8280 & idx_w_i[6];
  assign N8318 = N8281 & N1093;
  assign N8319 = N8281 & idx_w_i[6];
  assign N8320 = N8282 & N1093;
  assign N8321 = N8282 & idx_w_i[6];
  assign N8322 = N8283 & N1093;
  assign N8323 = N8283 & idx_w_i[6];
  assign N8324 = N2771 & N1093;
  assign N8325 = N2772 & N1093;
  assign N8326 = N2773 & N1093;
  assign N8327 = N2774 & N1093;
  assign N8328 = N2775 & N1093;
  assign N8329 = N2776 & N1093;
  assign N8330 = N2777 & N1093;
  assign N8331 = N2778 & N1093;
  assign N8332 = N5960 & N1093;
  assign N8333 = N5962 & N1093;
  assign N8334 = N5964 & N1093;
  assign N8335 = N5966 & N1093;
  assign N8336 = N5968 & N1093;
  assign N8337 = N5970 & N1093;
  assign N8338 = N5972 & N1093;
  assign N8339 = N5974 & N1093;
  assign N8340 = N2740 & N1093;
  assign N8341 = N2742 & N1093;
  assign N8342 = N2744 & N1093;
  assign N8343 = N2746 & N1093;
  assign N8344 = N2748 & N1093;
  assign N8345 = N2750 & N1093;
  assign N8346 = N2752 & N1093;
  assign N8347 = N2754 & N1093;
  assign N8348 = N11185 & N1093;
  assign N8349 = N11187 & N1093;
  assign N8350 = N11189 & N1093;
  assign N8351 = N11191 & N1093;
  assign N8352 = N11193 & N1093;
  assign N8353 = N11195 & N1093;
  assign N8354 = N11197 & N1093;
  assign N8355 = N11199 & N1093;
  assign N8356 = N11201 & N1093;
  assign N8357 = N11203 & N1093;
  assign N8358 = N11205 & N1093;
  assign N8359 = N11207 & N1093;
  assign N8360 = N11209 & N1093;
  assign N8361 = N11211 & N1093;
  assign N8362 = N11213 & N1093;
  assign N8363 = N11215 & N1093;
  assign N8364 = N8284 & N1190;
  assign N8365 = N8284 & idx_w_i[7];
  assign N8366 = N8286 & N1190;
  assign N8367 = N8286 & idx_w_i[7];
  assign N8368 = N8288 & N1190;
  assign N8369 = N8288 & idx_w_i[7];
  assign N8370 = N8290 & N1190;
  assign N8371 = N8290 & idx_w_i[7];
  assign N8372 = N8292 & N1190;
  assign N8373 = N8292 & idx_w_i[7];
  assign N8374 = N8294 & N1190;
  assign N8375 = N8294 & idx_w_i[7];
  assign N8376 = N8296 & N1190;
  assign N8377 = N8296 & idx_w_i[7];
  assign N8378 = N8298 & N1190;
  assign N8379 = N8298 & idx_w_i[7];
  assign N8380 = N8300 & N1190;
  assign N8381 = N8300 & idx_w_i[7];
  assign N8382 = N8301 & N1190;
  assign N8383 = N8301 & idx_w_i[7];
  assign N8384 = N8302 & N1190;
  assign N8385 = N8302 & idx_w_i[7];
  assign N8386 = N8303 & N1190;
  assign N8387 = N8303 & idx_w_i[7];
  assign N8388 = N8304 & N1190;
  assign N8389 = N8304 & idx_w_i[7];
  assign N8390 = N8305 & N1190;
  assign N8391 = N8305 & idx_w_i[7];
  assign N8392 = N8306 & N1190;
  assign N8393 = N8306 & idx_w_i[7];
  assign N8394 = N8307 & N1190;
  assign N8395 = N8307 & idx_w_i[7];
  assign N8396 = N8308 & N1190;
  assign N8397 = N8308 & idx_w_i[7];
  assign N8398 = N8310 & N1190;
  assign N8399 = N8310 & idx_w_i[7];
  assign N8400 = N8312 & N1190;
  assign N8401 = N8312 & idx_w_i[7];
  assign N8402 = N8314 & N1190;
  assign N8403 = N8314 & idx_w_i[7];
  assign N8404 = N8316 & N1190;
  assign N8405 = N8316 & idx_w_i[7];
  assign N8406 = N8318 & N1190;
  assign N8407 = N8318 & idx_w_i[7];
  assign N8408 = N8320 & N1190;
  assign N8409 = N8320 & idx_w_i[7];
  assign N8410 = N8322 & N1190;
  assign N8411 = N8322 & idx_w_i[7];
  assign N8412 = N8324 & N1190;
  assign N8413 = N8324 & idx_w_i[7];
  assign N8414 = N8325 & N1190;
  assign N8415 = N8325 & idx_w_i[7];
  assign N8416 = N8326 & N1190;
  assign N8417 = N8326 & idx_w_i[7];
  assign N8418 = N8327 & N1190;
  assign N8419 = N8327 & idx_w_i[7];
  assign N8420 = N8328 & N1190;
  assign N8421 = N8328 & idx_w_i[7];
  assign N8422 = N8329 & N1190;
  assign N8423 = N8329 & idx_w_i[7];
  assign N8424 = N8330 & N1190;
  assign N8425 = N8330 & idx_w_i[7];
  assign N8426 = N8331 & N1190;
  assign N8427 = N8331 & idx_w_i[7];
  assign N8428 = N8332 & N1190;
  assign N8429 = N8332 & idx_w_i[7];
  assign N8430 = N8333 & N1190;
  assign N8431 = N8333 & idx_w_i[7];
  assign N8432 = N8334 & N1190;
  assign N8433 = N8334 & idx_w_i[7];
  assign N8434 = N8335 & N1190;
  assign N8435 = N8335 & idx_w_i[7];
  assign N8436 = N8336 & N1190;
  assign N8437 = N8336 & idx_w_i[7];
  assign N8438 = N8337 & N1190;
  assign N8439 = N8337 & idx_w_i[7];
  assign N8440 = N8338 & N1190;
  assign N8441 = N8338 & idx_w_i[7];
  assign N8442 = N8339 & N1190;
  assign N8443 = N8339 & idx_w_i[7];
  assign N8444 = N8340 & N1190;
  assign N8445 = N8340 & idx_w_i[7];
  assign N8446 = N8341 & N1190;
  assign N8447 = N8341 & idx_w_i[7];
  assign N8448 = N8342 & N1190;
  assign N8449 = N8342 & idx_w_i[7];
  assign N8450 = N8343 & N1190;
  assign N8451 = N8343 & idx_w_i[7];
  assign N8452 = N8344 & N1190;
  assign N8453 = N8344 & idx_w_i[7];
  assign N8454 = N8345 & N1190;
  assign N8455 = N8345 & idx_w_i[7];
  assign N8456 = N8346 & N1190;
  assign N8457 = N8346 & idx_w_i[7];
  assign N8458 = N8347 & N1190;
  assign N8459 = N8347 & idx_w_i[7];
  assign N8460 = N8348 & N1190;
  assign N8461 = N8348 & idx_w_i[7];
  assign N8462 = N8349 & N1190;
  assign N8463 = N8349 & idx_w_i[7];
  assign N8464 = N8350 & N1190;
  assign N8465 = N8350 & idx_w_i[7];
  assign N8466 = N8351 & N1190;
  assign N8467 = N8351 & idx_w_i[7];
  assign N8468 = N8352 & N1190;
  assign N8469 = N8352 & idx_w_i[7];
  assign N8470 = N8353 & N1190;
  assign N8471 = N8353 & idx_w_i[7];
  assign N8472 = N8354 & N1190;
  assign N8473 = N8354 & idx_w_i[7];
  assign N8474 = N8355 & N1190;
  assign N8475 = N8355 & idx_w_i[7];
  assign N8476 = N8356 & N1190;
  assign N8477 = N8356 & idx_w_i[7];
  assign N8478 = N8357 & N1190;
  assign N8479 = N8357 & idx_w_i[7];
  assign N8480 = N8358 & N1190;
  assign N8481 = N8358 & idx_w_i[7];
  assign N8482 = N8359 & N1190;
  assign N8483 = N8359 & idx_w_i[7];
  assign N8484 = N8360 & N1190;
  assign N8485 = N8360 & idx_w_i[7];
  assign N8486 = N8361 & N1190;
  assign N8487 = N8361 & idx_w_i[7];
  assign N8488 = N8362 & N1190;
  assign N8489 = N8362 & idx_w_i[7];
  assign N8490 = N8363 & N1190;
  assign N8491 = N8363 & idx_w_i[7];
  assign N8492 = N8285 & N1190;
  assign N8493 = N8285 & idx_w_i[7];
  assign N8494 = N8287 & N1190;
  assign N8495 = N8287 & idx_w_i[7];
  assign N8496 = N8289 & N1190;
  assign N8497 = N8289 & idx_w_i[7];
  assign N8498 = N8291 & N1190;
  assign N8499 = N8291 & idx_w_i[7];
  assign N8500 = N8293 & N1190;
  assign N8501 = N8293 & idx_w_i[7];
  assign N8502 = N8295 & N1190;
  assign N8503 = N8295 & idx_w_i[7];
  assign N8504 = N8297 & N1190;
  assign N8505 = N8297 & idx_w_i[7];
  assign N8506 = N8299 & N1190;
  assign N8507 = N8299 & idx_w_i[7];
  assign N8508 = N2796 & N1190;
  assign N8509 = N2798 & N1190;
  assign N8510 = N2800 & N1190;
  assign N8511 = N2802 & N1190;
  assign N8512 = N2804 & N1190;
  assign N8513 = N2806 & N1190;
  assign N8514 = N2808 & N1190;
  assign N8515 = N2810 & N1190;
  assign N8516 = N8309 & N1190;
  assign N8517 = N8309 & idx_w_i[7];
  assign N8518 = N8311 & N1190;
  assign N8519 = N8311 & idx_w_i[7];
  assign N8520 = N8313 & N1190;
  assign N8521 = N8313 & idx_w_i[7];
  assign N8522 = N8315 & N1190;
  assign N8523 = N8315 & idx_w_i[7];
  assign N8524 = N8317 & N1190;
  assign N8525 = N8317 & idx_w_i[7];
  assign N8526 = N8319 & N1190;
  assign N8527 = N8319 & idx_w_i[7];
  assign N8528 = N8321 & N1190;
  assign N8529 = N8321 & idx_w_i[7];
  assign N8530 = N8323 & N1190;
  assign N8531 = N8323 & idx_w_i[7];
  assign N8532 = N2828 & N1190;
  assign N8533 = N2830 & N1190;
  assign N8534 = N2832 & N1190;
  assign N8535 = N2834 & N1190;
  assign N8536 = N2836 & N1190;
  assign N8537 = N2838 & N1190;
  assign N8538 = N2840 & N1190;
  assign N8539 = N2842 & N1190;
  assign N8540 = N6032 & N1190;
  assign N8541 = N6034 & N1190;
  assign N8542 = N6036 & N1190;
  assign N8543 = N6038 & N1190;
  assign N8544 = N6040 & N1190;
  assign N8545 = N6042 & N1190;
  assign N8546 = N6044 & N1190;
  assign N8547 = N6046 & N1190;
  assign N8548 = N2860 & N1190;
  assign N8549 = N2862 & N1190;
  assign N8550 = N2864 & N1190;
  assign N8551 = N2866 & N1190;
  assign N8552 = N2868 & N1190;
  assign N8553 = N2870 & N1190;
  assign N8554 = N2872 & N1190;
  assign N8555 = N2874 & N1190;
  assign N8556 = N11313 & N1190;
  assign N8557 = N11315 & N1190;
  assign N8558 = N11317 & N1190;
  assign N8559 = N11319 & N1190;
  assign N8560 = N11321 & N1190;
  assign N8561 = N11323 & N1190;
  assign N8562 = N11325 & N1190;
  assign N8563 = N11327 & N1190;
  assign N8564 = N11329 & N1190;
  assign N8565 = N11331 & N1190;
  assign N8566 = N11333 & N1190;
  assign N8567 = N11335 & N1190;
  assign N8568 = N11337 & N1190;
  assign N8569 = N11339 & N1190;
  assign N8570 = N11341 & N1190;
  assign N8571 = N11343 & N1190;
  assign N8572 = N8364 & N1415;
  assign N8573 = N8364 & idx_w_i[8];
  assign N8574 = N8366 & N1415;
  assign N8575 = N8366 & idx_w_i[8];
  assign N8576 = N8368 & N1415;
  assign N8577 = N8368 & idx_w_i[8];
  assign N8578 = N8370 & N1415;
  assign N8579 = N8370 & idx_w_i[8];
  assign N8580 = N8372 & N1415;
  assign N8581 = N8372 & idx_w_i[8];
  assign N8582 = N8374 & N1415;
  assign N8583 = N8374 & idx_w_i[8];
  assign N8584 = N8376 & N1415;
  assign N8585 = N8376 & idx_w_i[8];
  assign N8586 = N8378 & N1415;
  assign N8587 = N8378 & idx_w_i[8];
  assign N8588 = N8380 & N1415;
  assign N8589 = N8380 & idx_w_i[8];
  assign N8590 = N8382 & N1415;
  assign N8591 = N8382 & idx_w_i[8];
  assign N8592 = N8384 & N1415;
  assign N8593 = N8384 & idx_w_i[8];
  assign N8594 = N8386 & N1415;
  assign N8595 = N8386 & idx_w_i[8];
  assign N8596 = N8388 & N1415;
  assign N8597 = N8388 & idx_w_i[8];
  assign N8598 = N8390 & N1415;
  assign N8599 = N8390 & idx_w_i[8];
  assign N8600 = N8392 & N1415;
  assign N8601 = N8392 & idx_w_i[8];
  assign N8602 = N8394 & N1415;
  assign N8603 = N8394 & idx_w_i[8];
  assign N8604 = N8396 & N1415;
  assign N8605 = N8396 & idx_w_i[8];
  assign N8606 = N8398 & N1415;
  assign N8607 = N8398 & idx_w_i[8];
  assign N8608 = N8400 & N1415;
  assign N8609 = N8400 & idx_w_i[8];
  assign N8610 = N8402 & N1415;
  assign N8611 = N8402 & idx_w_i[8];
  assign N8612 = N8404 & N1415;
  assign N8613 = N8404 & idx_w_i[8];
  assign N8614 = N8406 & N1415;
  assign N8615 = N8406 & idx_w_i[8];
  assign N8616 = N8408 & N1415;
  assign N8617 = N8408 & idx_w_i[8];
  assign N8618 = N8410 & N1415;
  assign N8619 = N8410 & idx_w_i[8];
  assign N8620 = N8412 & N1415;
  assign N8621 = N8412 & idx_w_i[8];
  assign N8622 = N8414 & N1415;
  assign N8623 = N8414 & idx_w_i[8];
  assign N8624 = N8416 & N1415;
  assign N8625 = N8416 & idx_w_i[8];
  assign N8626 = N8418 & N1415;
  assign N8627 = N8418 & idx_w_i[8];
  assign N8628 = N8420 & N1415;
  assign N8629 = N8420 & idx_w_i[8];
  assign N8630 = N8422 & N1415;
  assign N8631 = N8422 & idx_w_i[8];
  assign N8632 = N8424 & N1415;
  assign N8633 = N8424 & idx_w_i[8];
  assign N8634 = N8426 & N1415;
  assign N8635 = N8426 & idx_w_i[8];
  assign N8636 = N8428 & N1415;
  assign N8637 = N8428 & idx_w_i[8];
  assign N8638 = N8430 & N1415;
  assign N8639 = N8430 & idx_w_i[8];
  assign N8640 = N8432 & N1415;
  assign N8641 = N8432 & idx_w_i[8];
  assign N8642 = N8434 & N1415;
  assign N8643 = N8434 & idx_w_i[8];
  assign N8644 = N8436 & N1415;
  assign N8645 = N8436 & idx_w_i[8];
  assign N8646 = N8438 & N1415;
  assign N8647 = N8438 & idx_w_i[8];
  assign N8648 = N8440 & N1415;
  assign N8649 = N8440 & idx_w_i[8];
  assign N8650 = N8442 & N1415;
  assign N8651 = N8442 & idx_w_i[8];
  assign N8652 = N8444 & N1415;
  assign N8653 = N8444 & idx_w_i[8];
  assign N8654 = N8446 & N1415;
  assign N8655 = N8446 & idx_w_i[8];
  assign N8656 = N8448 & N1415;
  assign N8657 = N8448 & idx_w_i[8];
  assign N8658 = N8450 & N1415;
  assign N8659 = N8450 & idx_w_i[8];
  assign N8660 = N8452 & N1415;
  assign N8661 = N8452 & idx_w_i[8];
  assign N8662 = N8454 & N1415;
  assign N8663 = N8454 & idx_w_i[8];
  assign N8664 = N8456 & N1415;
  assign N8665 = N8456 & idx_w_i[8];
  assign N8666 = N8458 & N1415;
  assign N8667 = N8458 & idx_w_i[8];
  assign N8668 = N8460 & N1415;
  assign N8669 = N8460 & idx_w_i[8];
  assign N8670 = N8462 & N1415;
  assign N8671 = N8462 & idx_w_i[8];
  assign N8672 = N8464 & N1415;
  assign N8673 = N8464 & idx_w_i[8];
  assign N8674 = N8466 & N1415;
  assign N8675 = N8466 & idx_w_i[8];
  assign N8676 = N8468 & N1415;
  assign N8677 = N8468 & idx_w_i[8];
  assign N8678 = N8470 & N1415;
  assign N8679 = N8470 & idx_w_i[8];
  assign N8680 = N8472 & N1415;
  assign N8681 = N8472 & idx_w_i[8];
  assign N8682 = N8474 & N1415;
  assign N8683 = N8474 & idx_w_i[8];
  assign N8684 = N8476 & N1415;
  assign N8685 = N8476 & idx_w_i[8];
  assign N8686 = N8478 & N1415;
  assign N8687 = N8478 & idx_w_i[8];
  assign N8688 = N8480 & N1415;
  assign N8689 = N8480 & idx_w_i[8];
  assign N8690 = N8482 & N1415;
  assign N8691 = N8482 & idx_w_i[8];
  assign N8692 = N8484 & N1415;
  assign N8693 = N8484 & idx_w_i[8];
  assign N8694 = N8486 & N1415;
  assign N8695 = N8486 & idx_w_i[8];
  assign N8696 = N8488 & N1415;
  assign N8697 = N8488 & idx_w_i[8];
  assign N8698 = N8490 & N1415;
  assign N8699 = N8490 & idx_w_i[8];
  assign N8700 = N8492 & N1415;
  assign N8701 = N8492 & idx_w_i[8];
  assign N8702 = N8494 & N1415;
  assign N8703 = N8494 & idx_w_i[8];
  assign N8704 = N8496 & N1415;
  assign N8705 = N8496 & idx_w_i[8];
  assign N8706 = N8498 & N1415;
  assign N8707 = N8498 & idx_w_i[8];
  assign N8708 = N8500 & N1415;
  assign N8709 = N8500 & idx_w_i[8];
  assign N8710 = N8502 & N1415;
  assign N8711 = N8502 & idx_w_i[8];
  assign N8712 = N8504 & N1415;
  assign N8713 = N8504 & idx_w_i[8];
  assign N8714 = N8506 & N1415;
  assign N8715 = N8506 & idx_w_i[8];
  assign N8716 = N8508 & N1415;
  assign N8717 = N8508 & idx_w_i[8];
  assign N8718 = N8509 & N1415;
  assign N8719 = N8509 & idx_w_i[8];
  assign N8720 = N8510 & N1415;
  assign N8721 = N8510 & idx_w_i[8];
  assign N8722 = N8511 & N1415;
  assign N8723 = N8511 & idx_w_i[8];
  assign N8724 = N8512 & N1415;
  assign N8725 = N8512 & idx_w_i[8];
  assign N8726 = N8513 & N1415;
  assign N8727 = N8513 & idx_w_i[8];
  assign N8728 = N8514 & N1415;
  assign N8729 = N8514 & idx_w_i[8];
  assign N8730 = N8515 & N1415;
  assign N8731 = N8515 & idx_w_i[8];
  assign N8732 = N8516 & N1415;
  assign N8733 = N8516 & idx_w_i[8];
  assign N8734 = N8518 & N1415;
  assign N8735 = N8518 & idx_w_i[8];
  assign N8736 = N8520 & N1415;
  assign N8737 = N8520 & idx_w_i[8];
  assign N8738 = N8522 & N1415;
  assign N8739 = N8522 & idx_w_i[8];
  assign N8740 = N8524 & N1415;
  assign N8741 = N8524 & idx_w_i[8];
  assign N8742 = N8526 & N1415;
  assign N8743 = N8526 & idx_w_i[8];
  assign N8744 = N8528 & N1415;
  assign N8745 = N8528 & idx_w_i[8];
  assign N8746 = N8530 & N1415;
  assign N8747 = N8530 & idx_w_i[8];
  assign N8748 = N8532 & N1415;
  assign N8749 = N8532 & idx_w_i[8];
  assign N8750 = N8533 & N1415;
  assign N8751 = N8533 & idx_w_i[8];
  assign N8752 = N8534 & N1415;
  assign N8753 = N8534 & idx_w_i[8];
  assign N8754 = N8535 & N1415;
  assign N8755 = N8535 & idx_w_i[8];
  assign N8756 = N8536 & N1415;
  assign N8757 = N8536 & idx_w_i[8];
  assign N8758 = N8537 & N1415;
  assign N8759 = N8537 & idx_w_i[8];
  assign N8760 = N8538 & N1415;
  assign N8761 = N8538 & idx_w_i[8];
  assign N8762 = N8539 & N1415;
  assign N8763 = N8539 & idx_w_i[8];
  assign N8764 = N8540 & N1415;
  assign N8765 = N8540 & idx_w_i[8];
  assign N8766 = N8541 & N1415;
  assign N8767 = N8541 & idx_w_i[8];
  assign N8768 = N8542 & N1415;
  assign N8769 = N8542 & idx_w_i[8];
  assign N8770 = N8543 & N1415;
  assign N8771 = N8543 & idx_w_i[8];
  assign N8772 = N8544 & N1415;
  assign N8773 = N8544 & idx_w_i[8];
  assign N8774 = N8545 & N1415;
  assign N8775 = N8545 & idx_w_i[8];
  assign N8776 = N8546 & N1415;
  assign N8777 = N8546 & idx_w_i[8];
  assign N8778 = N8547 & N1415;
  assign N8779 = N8547 & idx_w_i[8];
  assign N8780 = N8548 & N1415;
  assign N8781 = N8548 & idx_w_i[8];
  assign N8782 = N8549 & N1415;
  assign N8783 = N8549 & idx_w_i[8];
  assign N8784 = N8550 & N1415;
  assign N8785 = N8550 & idx_w_i[8];
  assign N8786 = N8551 & N1415;
  assign N8787 = N8551 & idx_w_i[8];
  assign N8788 = N8552 & N1415;
  assign N8789 = N8552 & idx_w_i[8];
  assign N8790 = N8553 & N1415;
  assign N8791 = N8553 & idx_w_i[8];
  assign N8792 = N8554 & N1415;
  assign N8793 = N8554 & idx_w_i[8];
  assign N8794 = N8555 & N1415;
  assign N8795 = N8555 & idx_w_i[8];
  assign N8796 = N8556 & N1415;
  assign N8797 = N8556 & idx_w_i[8];
  assign N8798 = N8557 & N1415;
  assign N8799 = N8557 & idx_w_i[8];
  assign N8800 = N8558 & N1415;
  assign N8801 = N8558 & idx_w_i[8];
  assign N8802 = N8559 & N1415;
  assign N8803 = N8559 & idx_w_i[8];
  assign N8804 = N8560 & N1415;
  assign N8805 = N8560 & idx_w_i[8];
  assign N8806 = N8561 & N1415;
  assign N8807 = N8561 & idx_w_i[8];
  assign N8808 = N8562 & N1415;
  assign N8809 = N8562 & idx_w_i[8];
  assign N8810 = N8563 & N1415;
  assign N8811 = N8563 & idx_w_i[8];
  assign N8812 = N8564 & N1415;
  assign N8813 = N8564 & idx_w_i[8];
  assign N8814 = N8565 & N1415;
  assign N8815 = N8565 & idx_w_i[8];
  assign N8816 = N8566 & N1415;
  assign N8817 = N8566 & idx_w_i[8];
  assign N8818 = N8567 & N1415;
  assign N8819 = N8567 & idx_w_i[8];
  assign N8820 = N8568 & N1415;
  assign N8821 = N8568 & idx_w_i[8];
  assign N8822 = N8569 & N1415;
  assign N8823 = N8569 & idx_w_i[8];
  assign N8824 = N8570 & N1415;
  assign N8825 = N8570 & idx_w_i[8];
  assign N8826 = N8571 & N1415;
  assign N8827 = N8571 & idx_w_i[8];
  assign N8828 = N8365 & N1415;
  assign N8829 = N8365 & idx_w_i[8];
  assign N8830 = N8367 & N1415;
  assign N8831 = N8367 & idx_w_i[8];
  assign N8832 = N8369 & N1415;
  assign N8833 = N8369 & idx_w_i[8];
  assign N8834 = N8371 & N1415;
  assign N8835 = N8371 & idx_w_i[8];
  assign N8836 = N8373 & N1415;
  assign N8837 = N8373 & idx_w_i[8];
  assign N8838 = N8375 & N1415;
  assign N8839 = N8375 & idx_w_i[8];
  assign N8840 = N8377 & N1415;
  assign N8841 = N8377 & idx_w_i[8];
  assign N8842 = N8379 & N1415;
  assign N8843 = N8379 & idx_w_i[8];
  assign N8844 = N8381 & N1415;
  assign N8845 = N8381 & idx_w_i[8];
  assign N8846 = N8383 & N1415;
  assign N8847 = N8383 & idx_w_i[8];
  assign N8848 = N8385 & N1415;
  assign N8849 = N8385 & idx_w_i[8];
  assign N8850 = N8387 & N1415;
  assign N8851 = N8387 & idx_w_i[8];
  assign N8852 = N8389 & N1415;
  assign N8853 = N8389 & idx_w_i[8];
  assign N8854 = N8391 & N1415;
  assign N8855 = N8391 & idx_w_i[8];
  assign N8856 = N8393 & N1415;
  assign N8857 = N8393 & idx_w_i[8];
  assign N8858 = N8395 & N1415;
  assign N8859 = N8395 & idx_w_i[8];
  assign N8860 = N8397 & N1415;
  assign N8861 = N8397 & idx_w_i[8];
  assign N8862 = N8399 & N1415;
  assign N8863 = N8399 & idx_w_i[8];
  assign N8864 = N8401 & N1415;
  assign N8865 = N8401 & idx_w_i[8];
  assign N8866 = N8403 & N1415;
  assign N8867 = N8403 & idx_w_i[8];
  assign N8868 = N8405 & N1415;
  assign N8869 = N8405 & idx_w_i[8];
  assign N8870 = N8407 & N1415;
  assign N8871 = N8407 & idx_w_i[8];
  assign N8872 = N8409 & N1415;
  assign N8873 = N8409 & idx_w_i[8];
  assign N8874 = N8411 & N1415;
  assign N8875 = N8411 & idx_w_i[8];
  assign N8876 = N8413 & N1415;
  assign N8877 = N8413 & idx_w_i[8];
  assign N8878 = N8415 & N1415;
  assign N8879 = N8415 & idx_w_i[8];
  assign N8880 = N8417 & N1415;
  assign N8881 = N8417 & idx_w_i[8];
  assign N8882 = N8419 & N1415;
  assign N8883 = N8419 & idx_w_i[8];
  assign N8884 = N8421 & N1415;
  assign N8885 = N8421 & idx_w_i[8];
  assign N8886 = N8423 & N1415;
  assign N8887 = N8423 & idx_w_i[8];
  assign N8888 = N8425 & N1415;
  assign N8889 = N8425 & idx_w_i[8];
  assign N8890 = N8427 & N1415;
  assign N8891 = N8427 & idx_w_i[8];
  assign N8892 = N8429 & N1415;
  assign N8893 = N8429 & idx_w_i[8];
  assign N8894 = N8431 & N1415;
  assign N8895 = N8431 & idx_w_i[8];
  assign N8896 = N8433 & N1415;
  assign N8897 = N8433 & idx_w_i[8];
  assign N8898 = N8435 & N1415;
  assign N8899 = N8435 & idx_w_i[8];
  assign N8900 = N8437 & N1415;
  assign N8901 = N8437 & idx_w_i[8];
  assign N8902 = N8439 & N1415;
  assign N8903 = N8439 & idx_w_i[8];
  assign N8904 = N8441 & N1415;
  assign N8905 = N8441 & idx_w_i[8];
  assign N8906 = N8443 & N1415;
  assign N8907 = N8443 & idx_w_i[8];
  assign N8908 = N8445 & N1415;
  assign N8909 = N8445 & idx_w_i[8];
  assign N8910 = N8447 & N1415;
  assign N8911 = N8447 & idx_w_i[8];
  assign N8912 = N8449 & N1415;
  assign N8913 = N8449 & idx_w_i[8];
  assign N8914 = N8451 & N1415;
  assign N8915 = N8451 & idx_w_i[8];
  assign N8916 = N8453 & N1415;
  assign N8917 = N8453 & idx_w_i[8];
  assign N8918 = N8455 & N1415;
  assign N8919 = N8455 & idx_w_i[8];
  assign N8920 = N8457 & N1415;
  assign N8921 = N8457 & idx_w_i[8];
  assign N8922 = N8459 & N1415;
  assign N8923 = N8459 & idx_w_i[8];
  assign N8924 = N8461 & N1415;
  assign N8925 = N8461 & idx_w_i[8];
  assign N8926 = N8463 & N1415;
  assign N8927 = N8463 & idx_w_i[8];
  assign N8928 = N8465 & N1415;
  assign N8929 = N8465 & idx_w_i[8];
  assign N8930 = N8467 & N1415;
  assign N8931 = N8467 & idx_w_i[8];
  assign N8932 = N8469 & N1415;
  assign N8933 = N8469 & idx_w_i[8];
  assign N8934 = N8471 & N1415;
  assign N8935 = N8471 & idx_w_i[8];
  assign N8936 = N8473 & N1415;
  assign N8937 = N8473 & idx_w_i[8];
  assign N8938 = N8475 & N1415;
  assign N8939 = N8475 & idx_w_i[8];
  assign N8940 = N8477 & N1415;
  assign N8941 = N8477 & idx_w_i[8];
  assign N8942 = N8479 & N1415;
  assign N8943 = N8479 & idx_w_i[8];
  assign N8944 = N8481 & N1415;
  assign N8945 = N8481 & idx_w_i[8];
  assign N8946 = N8483 & N1415;
  assign N8947 = N8483 & idx_w_i[8];
  assign N8948 = N8485 & N1415;
  assign N8949 = N8485 & idx_w_i[8];
  assign N8950 = N8487 & N1415;
  assign N8951 = N8487 & idx_w_i[8];
  assign N8952 = N8489 & N1415;
  assign N8953 = N8489 & idx_w_i[8];
  assign N8954 = N8491 & N1415;
  assign N8955 = N8491 & idx_w_i[8];
  assign N8956 = N8493 & N1415;
  assign N8957 = N8493 & idx_w_i[8];
  assign N8958 = N8495 & N1415;
  assign N8959 = N8495 & idx_w_i[8];
  assign N8960 = N8497 & N1415;
  assign N8961 = N8497 & idx_w_i[8];
  assign N8962 = N8499 & N1415;
  assign N8963 = N8499 & idx_w_i[8];
  assign N8964 = N8501 & N1415;
  assign N8965 = N8501 & idx_w_i[8];
  assign N8966 = N8503 & N1415;
  assign N8967 = N8503 & idx_w_i[8];
  assign N8968 = N8505 & N1415;
  assign N8969 = N8505 & idx_w_i[8];
  assign N8970 = N8507 & N1415;
  assign N8971 = N8507 & idx_w_i[8];
  assign N8972 = N3044 & N1415;
  assign N8973 = N3046 & N1415;
  assign N8974 = N3048 & N1415;
  assign N8975 = N3050 & N1415;
  assign N8976 = N3052 & N1415;
  assign N8977 = N3054 & N1415;
  assign N8978 = N3056 & N1415;
  assign N8979 = N3058 & N1415;
  assign N8980 = N8517 & N1415;
  assign N8981 = N8517 & idx_w_i[8];
  assign N8982 = N8519 & N1415;
  assign N8983 = N8519 & idx_w_i[8];
  assign N8984 = N8521 & N1415;
  assign N8985 = N8521 & idx_w_i[8];
  assign N8986 = N8523 & N1415;
  assign N8987 = N8523 & idx_w_i[8];
  assign N8988 = N8525 & N1415;
  assign N8989 = N8525 & idx_w_i[8];
  assign N8990 = N8527 & N1415;
  assign N8991 = N8527 & idx_w_i[8];
  assign N8992 = N8529 & N1415;
  assign N8993 = N8529 & idx_w_i[8];
  assign N8994 = N8531 & N1415;
  assign N8995 = N8531 & idx_w_i[8];
  assign N8996 = N3076 & N1415;
  assign N8997 = N3078 & N1415;
  assign N8998 = N3080 & N1415;
  assign N8999 = N3082 & N1415;
  assign N9000 = N3084 & N1415;
  assign N9001 = N3086 & N1415;
  assign N9002 = N3088 & N1415;
  assign N9003 = N3090 & N1415;
  assign N9004 = N6248 & N1415;
  assign N9005 = N6250 & N1415;
  assign N9006 = N6252 & N1415;
  assign N9007 = N6254 & N1415;
  assign N9008 = N6256 & N1415;
  assign N9009 = N6258 & N1415;
  assign N9010 = N6260 & N1415;
  assign N9011 = N6262 & N1415;
  assign N9012 = N3108 & N1415;
  assign N9013 = N3110 & N1415;
  assign N9014 = N3112 & N1415;
  assign N9015 = N3114 & N1415;
  assign N9016 = N3116 & N1415;
  assign N9017 = N3118 & N1415;
  assign N9018 = N3120 & N1415;
  assign N9019 = N3122 & N1415;
  assign N9020 = N11569 & N1415;
  assign N9021 = N11571 & N1415;
  assign N9022 = N11573 & N1415;
  assign N9023 = N11575 & N1415;
  assign N9024 = N11577 & N1415;
  assign N9025 = N11579 & N1415;
  assign N9026 = N11581 & N1415;
  assign N9027 = N11583 & N1415;
  assign N9028 = N11585 & N1415;
  assign N9029 = N11587 & N1415;
  assign N9030 = N11589 & N1415;
  assign N9031 = N11591 & N1415;
  assign N9032 = N11593 & N1415;
  assign N9033 = N11595 & N1415;
  assign N9034 = N11597 & N1415;
  assign N9035 = N11599 & N1415;
  assign N9037 = N8268 & N1093;
  assign N9038 = N8269 & N1093;
  assign N9039 = N8270 & N1093;
  assign N9040 = N8271 & N1093;
  assign N9041 = N8272 & N1093;
  assign N9042 = N8273 & N1093;
  assign N9043 = N8274 & N1093;
  assign N9044 = N8275 & N1093;
  assign N9045 = N2739 & N1093;
  assign N9046 = N2741 & N1093;
  assign N9047 = N2743 & N1093;
  assign N9048 = N2745 & N1093;
  assign N9049 = N2747 & N1093;
  assign N9050 = N2749 & N1093;
  assign N9051 = N2751 & N1093;
  assign N9052 = N2753 & N1093;
  assign N9053 = N8276 & N1093;
  assign N9054 = N8277 & N1093;
  assign N9055 = N8278 & N1093;
  assign N9056 = N8279 & N1093;
  assign N9057 = N8280 & N1093;
  assign N9058 = N8281 & N1093;
  assign N9059 = N8282 & N1093;
  assign N9060 = N8283 & N1093;
  assign N9061 = N2771 & N1093;
  assign N9062 = N2772 & N1093;
  assign N9063 = N2773 & N1093;
  assign N9064 = N2774 & N1093;
  assign N9065 = N2775 & N1093;
  assign N9066 = N2776 & N1093;
  assign N9067 = N2777 & N1093;
  assign N9068 = N2778 & N1093;
  assign N9069 = N5960 & N1093;
  assign N9070 = N5962 & N1093;
  assign N9071 = N5964 & N1093;
  assign N9072 = N5966 & N1093;
  assign N9073 = N5968 & N1093;
  assign N9074 = N5970 & N1093;
  assign N9075 = N5972 & N1093;
  assign N9076 = N5974 & N1093;
  assign N9077 = N2740 & N1093;
  assign N9078 = N2742 & N1093;
  assign N9079 = N2744 & N1093;
  assign N9080 = N2746 & N1093;
  assign N9081 = N2748 & N1093;
  assign N9082 = N2750 & N1093;
  assign N9083 = N2752 & N1093;
  assign N9084 = N2754 & N1093;
  assign N9085 = N11185 & N1093;
  assign N9086 = N11187 & N1093;
  assign N9087 = N11189 & N1093;
  assign N9088 = N11191 & N1093;
  assign N9089 = N11193 & N1093;
  assign N9090 = N11195 & N1093;
  assign N9091 = N11197 & N1093;
  assign N9092 = N11199 & N1093;
  assign N9093 = N11201 & N1093;
  assign N9094 = N11203 & N1093;
  assign N9095 = N11205 & N1093;
  assign N9096 = N11207 & N1093;
  assign N9097 = N11209 & N1093;
  assign N9098 = N11211 & N1093;
  assign N9099 = N11213 & N1093;
  assign N9100 = N11215 & N1093;
  assign N9101 = N9037 & N1190;
  assign N9102 = N9037 & idx_w_i[7];
  assign N9103 = N9038 & N1190;
  assign N9104 = N9038 & idx_w_i[7];
  assign N9105 = N9039 & N1190;
  assign N9106 = N9039 & idx_w_i[7];
  assign N9107 = N9040 & N1190;
  assign N9108 = N9040 & idx_w_i[7];
  assign N9109 = N9041 & N1190;
  assign N9110 = N9041 & idx_w_i[7];
  assign N9111 = N9042 & N1190;
  assign N9112 = N9042 & idx_w_i[7];
  assign N9113 = N9043 & N1190;
  assign N9114 = N9043 & idx_w_i[7];
  assign N9115 = N9044 & N1190;
  assign N9116 = N9044 & idx_w_i[7];
  assign N9117 = N9045 & N1190;
  assign N9118 = N9045 & idx_w_i[7];
  assign N9119 = N9046 & N1190;
  assign N9120 = N9046 & idx_w_i[7];
  assign N9121 = N9047 & N1190;
  assign N9122 = N9047 & idx_w_i[7];
  assign N9123 = N9048 & N1190;
  assign N9124 = N9048 & idx_w_i[7];
  assign N9125 = N9049 & N1190;
  assign N9126 = N9049 & idx_w_i[7];
  assign N9127 = N9050 & N1190;
  assign N9128 = N9050 & idx_w_i[7];
  assign N9129 = N9051 & N1190;
  assign N9130 = N9051 & idx_w_i[7];
  assign N9131 = N9052 & N1190;
  assign N9132 = N9052 & idx_w_i[7];
  assign N9133 = N9053 & N1190;
  assign N9134 = N9053 & idx_w_i[7];
  assign N9135 = N9054 & N1190;
  assign N9136 = N9054 & idx_w_i[7];
  assign N9137 = N9055 & N1190;
  assign N9138 = N9055 & idx_w_i[7];
  assign N9139 = N9056 & N1190;
  assign N9140 = N9056 & idx_w_i[7];
  assign N9141 = N9057 & N1190;
  assign N9142 = N9057 & idx_w_i[7];
  assign N9143 = N9058 & N1190;
  assign N9144 = N9058 & idx_w_i[7];
  assign N9145 = N9059 & N1190;
  assign N9146 = N9059 & idx_w_i[7];
  assign N9147 = N9060 & N1190;
  assign N9148 = N9060 & idx_w_i[7];
  assign N9149 = N9061 & N1190;
  assign N9150 = N9061 & idx_w_i[7];
  assign N9151 = N9062 & N1190;
  assign N9152 = N9062 & idx_w_i[7];
  assign N9153 = N9063 & N1190;
  assign N9154 = N9063 & idx_w_i[7];
  assign N9155 = N9064 & N1190;
  assign N9156 = N9064 & idx_w_i[7];
  assign N9157 = N9065 & N1190;
  assign N9158 = N9065 & idx_w_i[7];
  assign N9159 = N9066 & N1190;
  assign N9160 = N9066 & idx_w_i[7];
  assign N9161 = N9067 & N1190;
  assign N9162 = N9067 & idx_w_i[7];
  assign N9163 = N9068 & N1190;
  assign N9164 = N9068 & idx_w_i[7];
  assign N9165 = N9069 & N1190;
  assign N9166 = N9069 & idx_w_i[7];
  assign N9167 = N9070 & N1190;
  assign N9168 = N9070 & idx_w_i[7];
  assign N9169 = N9071 & N1190;
  assign N9170 = N9071 & idx_w_i[7];
  assign N9171 = N9072 & N1190;
  assign N9172 = N9072 & idx_w_i[7];
  assign N9173 = N9073 & N1190;
  assign N9174 = N9073 & idx_w_i[7];
  assign N9175 = N9074 & N1190;
  assign N9176 = N9074 & idx_w_i[7];
  assign N9177 = N9075 & N1190;
  assign N9178 = N9075 & idx_w_i[7];
  assign N9179 = N9076 & N1190;
  assign N9180 = N9076 & idx_w_i[7];
  assign N9181 = N9077 & N1190;
  assign N9182 = N9077 & idx_w_i[7];
  assign N9183 = N9078 & N1190;
  assign N9184 = N9078 & idx_w_i[7];
  assign N9185 = N9079 & N1190;
  assign N9186 = N9079 & idx_w_i[7];
  assign N9187 = N9080 & N1190;
  assign N9188 = N9080 & idx_w_i[7];
  assign N9189 = N9081 & N1190;
  assign N9190 = N9081 & idx_w_i[7];
  assign N9191 = N9082 & N1190;
  assign N9192 = N9082 & idx_w_i[7];
  assign N9193 = N9083 & N1190;
  assign N9194 = N9083 & idx_w_i[7];
  assign N9195 = N9084 & N1190;
  assign N9196 = N9084 & idx_w_i[7];
  assign N9197 = N9085 & N1190;
  assign N9198 = N9085 & idx_w_i[7];
  assign N9199 = N9086 & N1190;
  assign N9200 = N9086 & idx_w_i[7];
  assign N9201 = N9087 & N1190;
  assign N9202 = N9087 & idx_w_i[7];
  assign N9203 = N9088 & N1190;
  assign N9204 = N9088 & idx_w_i[7];
  assign N9205 = N9089 & N1190;
  assign N9206 = N9089 & idx_w_i[7];
  assign N9207 = N9090 & N1190;
  assign N9208 = N9090 & idx_w_i[7];
  assign N9209 = N9091 & N1190;
  assign N9210 = N9091 & idx_w_i[7];
  assign N9211 = N9092 & N1190;
  assign N9212 = N9092 & idx_w_i[7];
  assign N9213 = N9093 & N1190;
  assign N9214 = N9093 & idx_w_i[7];
  assign N9215 = N9094 & N1190;
  assign N9216 = N9094 & idx_w_i[7];
  assign N9217 = N9095 & N1190;
  assign N9218 = N9095 & idx_w_i[7];
  assign N9219 = N9096 & N1190;
  assign N9220 = N9096 & idx_w_i[7];
  assign N9221 = N9097 & N1190;
  assign N9222 = N9097 & idx_w_i[7];
  assign N9223 = N9098 & N1190;
  assign N9224 = N9098 & idx_w_i[7];
  assign N9225 = N9099 & N1190;
  assign N9226 = N9099 & idx_w_i[7];
  assign N9227 = N9100 & N1190;
  assign N9228 = N9100 & idx_w_i[7];
  assign N9229 = N8285 & N1190;
  assign N9230 = N8287 & N1190;
  assign N9231 = N8289 & N1190;
  assign N9232 = N8291 & N1190;
  assign N9233 = N8293 & N1190;
  assign N9234 = N8295 & N1190;
  assign N9235 = N8297 & N1190;
  assign N9236 = N8299 & N1190;
  assign N9237 = N2796 & N1190;
  assign N9238 = N2798 & N1190;
  assign N9239 = N2800 & N1190;
  assign N9240 = N2802 & N1190;
  assign N9241 = N2804 & N1190;
  assign N9242 = N2806 & N1190;
  assign N9243 = N2808 & N1190;
  assign N9244 = N2810 & N1190;
  assign N9245 = N8309 & N1190;
  assign N9246 = N8311 & N1190;
  assign N9247 = N8313 & N1190;
  assign N9248 = N8315 & N1190;
  assign N9249 = N8317 & N1190;
  assign N9250 = N8319 & N1190;
  assign N9251 = N8321 & N1190;
  assign N9252 = N8323 & N1190;
  assign N9253 = N2828 & N1190;
  assign N9254 = N2830 & N1190;
  assign N9255 = N2832 & N1190;
  assign N9256 = N2834 & N1190;
  assign N9257 = N2836 & N1190;
  assign N9258 = N2838 & N1190;
  assign N9259 = N2840 & N1190;
  assign N9260 = N2842 & N1190;
  assign N9261 = N6032 & N1190;
  assign N9262 = N6034 & N1190;
  assign N9263 = N6036 & N1190;
  assign N9264 = N6038 & N1190;
  assign N9265 = N6040 & N1190;
  assign N9266 = N6042 & N1190;
  assign N9267 = N6044 & N1190;
  assign N9268 = N6046 & N1190;
  assign N9269 = N2860 & N1190;
  assign N9270 = N2862 & N1190;
  assign N9271 = N2864 & N1190;
  assign N9272 = N2866 & N1190;
  assign N9273 = N2868 & N1190;
  assign N9274 = N2870 & N1190;
  assign N9275 = N2872 & N1190;
  assign N9276 = N2874 & N1190;
  assign N9277 = N11313 & N1190;
  assign N9278 = N11315 & N1190;
  assign N9279 = N11317 & N1190;
  assign N9280 = N11319 & N1190;
  assign N9281 = N11321 & N1190;
  assign N9282 = N11323 & N1190;
  assign N9283 = N11325 & N1190;
  assign N9284 = N11327 & N1190;
  assign N9285 = N11329 & N1190;
  assign N9286 = N11331 & N1190;
  assign N9287 = N11333 & N1190;
  assign N9288 = N11335 & N1190;
  assign N9289 = N11337 & N1190;
  assign N9290 = N11339 & N1190;
  assign N9291 = N11341 & N1190;
  assign N9292 = N11343 & N1190;
  assign N9293 = N9101 & N1415;
  assign N9294 = N9101 & idx_w_i[8];
  assign N9295 = N9103 & N1415;
  assign N9296 = N9103 & idx_w_i[8];
  assign N9297 = N9105 & N1415;
  assign N9298 = N9105 & idx_w_i[8];
  assign N9299 = N9107 & N1415;
  assign N9300 = N9107 & idx_w_i[8];
  assign N9301 = N9109 & N1415;
  assign N9302 = N9109 & idx_w_i[8];
  assign N9303 = N9111 & N1415;
  assign N9304 = N9111 & idx_w_i[8];
  assign N9305 = N9113 & N1415;
  assign N9306 = N9113 & idx_w_i[8];
  assign N9307 = N9115 & N1415;
  assign N9308 = N9115 & idx_w_i[8];
  assign N9309 = N9117 & N1415;
  assign N9310 = N9117 & idx_w_i[8];
  assign N9311 = N9119 & N1415;
  assign N9312 = N9119 & idx_w_i[8];
  assign N9313 = N9121 & N1415;
  assign N9314 = N9121 & idx_w_i[8];
  assign N9315 = N9123 & N1415;
  assign N9316 = N9123 & idx_w_i[8];
  assign N9317 = N9125 & N1415;
  assign N9318 = N9125 & idx_w_i[8];
  assign N9319 = N9127 & N1415;
  assign N9320 = N9127 & idx_w_i[8];
  assign N9321 = N9129 & N1415;
  assign N9322 = N9129 & idx_w_i[8];
  assign N9323 = N9131 & N1415;
  assign N9324 = N9131 & idx_w_i[8];
  assign N9325 = N9133 & N1415;
  assign N9326 = N9133 & idx_w_i[8];
  assign N9327 = N9135 & N1415;
  assign N9328 = N9135 & idx_w_i[8];
  assign N9329 = N9137 & N1415;
  assign N9330 = N9137 & idx_w_i[8];
  assign N9331 = N9139 & N1415;
  assign N9332 = N9139 & idx_w_i[8];
  assign N9333 = N9141 & N1415;
  assign N9334 = N9141 & idx_w_i[8];
  assign N9335 = N9143 & N1415;
  assign N9336 = N9143 & idx_w_i[8];
  assign N9337 = N9145 & N1415;
  assign N9338 = N9145 & idx_w_i[8];
  assign N9339 = N9147 & N1415;
  assign N9340 = N9147 & idx_w_i[8];
  assign N9341 = N9149 & N1415;
  assign N9342 = N9149 & idx_w_i[8];
  assign N9343 = N9151 & N1415;
  assign N9344 = N9151 & idx_w_i[8];
  assign N9345 = N9153 & N1415;
  assign N9346 = N9153 & idx_w_i[8];
  assign N9347 = N9155 & N1415;
  assign N9348 = N9155 & idx_w_i[8];
  assign N9349 = N9157 & N1415;
  assign N9350 = N9157 & idx_w_i[8];
  assign N9351 = N9159 & N1415;
  assign N9352 = N9159 & idx_w_i[8];
  assign N9353 = N9161 & N1415;
  assign N9354 = N9161 & idx_w_i[8];
  assign N9355 = N9163 & N1415;
  assign N9356 = N9163 & idx_w_i[8];
  assign N9357 = N9165 & N1415;
  assign N9358 = N9165 & idx_w_i[8];
  assign N9359 = N9167 & N1415;
  assign N9360 = N9167 & idx_w_i[8];
  assign N9361 = N9169 & N1415;
  assign N9362 = N9169 & idx_w_i[8];
  assign N9363 = N9171 & N1415;
  assign N9364 = N9171 & idx_w_i[8];
  assign N9365 = N9173 & N1415;
  assign N9366 = N9173 & idx_w_i[8];
  assign N9367 = N9175 & N1415;
  assign N9368 = N9175 & idx_w_i[8];
  assign N9369 = N9177 & N1415;
  assign N9370 = N9177 & idx_w_i[8];
  assign N9371 = N9179 & N1415;
  assign N9372 = N9179 & idx_w_i[8];
  assign N9373 = N9181 & N1415;
  assign N9374 = N9181 & idx_w_i[8];
  assign N9375 = N9183 & N1415;
  assign N9376 = N9183 & idx_w_i[8];
  assign N9377 = N9185 & N1415;
  assign N9378 = N9185 & idx_w_i[8];
  assign N9379 = N9187 & N1415;
  assign N9380 = N9187 & idx_w_i[8];
  assign N9381 = N9189 & N1415;
  assign N9382 = N9189 & idx_w_i[8];
  assign N9383 = N9191 & N1415;
  assign N9384 = N9191 & idx_w_i[8];
  assign N9385 = N9193 & N1415;
  assign N9386 = N9193 & idx_w_i[8];
  assign N9387 = N9195 & N1415;
  assign N9388 = N9195 & idx_w_i[8];
  assign N9389 = N9197 & N1415;
  assign N9390 = N9197 & idx_w_i[8];
  assign N9391 = N9199 & N1415;
  assign N9392 = N9199 & idx_w_i[8];
  assign N9393 = N9201 & N1415;
  assign N9394 = N9201 & idx_w_i[8];
  assign N9395 = N9203 & N1415;
  assign N9396 = N9203 & idx_w_i[8];
  assign N9397 = N9205 & N1415;
  assign N9398 = N9205 & idx_w_i[8];
  assign N9399 = N9207 & N1415;
  assign N9400 = N9207 & idx_w_i[8];
  assign N9401 = N9209 & N1415;
  assign N9402 = N9209 & idx_w_i[8];
  assign N9403 = N9211 & N1415;
  assign N9404 = N9211 & idx_w_i[8];
  assign N9405 = N9213 & N1415;
  assign N9406 = N9213 & idx_w_i[8];
  assign N9407 = N9215 & N1415;
  assign N9408 = N9215 & idx_w_i[8];
  assign N9409 = N9217 & N1415;
  assign N9410 = N9217 & idx_w_i[8];
  assign N9411 = N9219 & N1415;
  assign N9412 = N9219 & idx_w_i[8];
  assign N9413 = N9221 & N1415;
  assign N9414 = N9221 & idx_w_i[8];
  assign N9415 = N9223 & N1415;
  assign N9416 = N9223 & idx_w_i[8];
  assign N9417 = N9225 & N1415;
  assign N9418 = N9225 & idx_w_i[8];
  assign N9419 = N9227 & N1415;
  assign N9420 = N9227 & idx_w_i[8];
  assign N9421 = N9229 & N1415;
  assign N9422 = N9229 & idx_w_i[8];
  assign N9423 = N9230 & N1415;
  assign N9424 = N9230 & idx_w_i[8];
  assign N9425 = N9231 & N1415;
  assign N9426 = N9231 & idx_w_i[8];
  assign N9427 = N9232 & N1415;
  assign N9428 = N9232 & idx_w_i[8];
  assign N9429 = N9233 & N1415;
  assign N9430 = N9233 & idx_w_i[8];
  assign N9431 = N9234 & N1415;
  assign N9432 = N9234 & idx_w_i[8];
  assign N9433 = N9235 & N1415;
  assign N9434 = N9235 & idx_w_i[8];
  assign N9435 = N9236 & N1415;
  assign N9436 = N9236 & idx_w_i[8];
  assign N9437 = N9237 & N1415;
  assign N9438 = N9237 & idx_w_i[8];
  assign N9439 = N9238 & N1415;
  assign N9440 = N9238 & idx_w_i[8];
  assign N9441 = N9239 & N1415;
  assign N9442 = N9239 & idx_w_i[8];
  assign N9443 = N9240 & N1415;
  assign N9444 = N9240 & idx_w_i[8];
  assign N9445 = N9241 & N1415;
  assign N9446 = N9241 & idx_w_i[8];
  assign N9447 = N9242 & N1415;
  assign N9448 = N9242 & idx_w_i[8];
  assign N9449 = N9243 & N1415;
  assign N9450 = N9243 & idx_w_i[8];
  assign N9451 = N9244 & N1415;
  assign N9452 = N9244 & idx_w_i[8];
  assign N9453 = N9245 & N1415;
  assign N9454 = N9245 & idx_w_i[8];
  assign N9455 = N9246 & N1415;
  assign N9456 = N9246 & idx_w_i[8];
  assign N9457 = N9247 & N1415;
  assign N9458 = N9247 & idx_w_i[8];
  assign N9459 = N9248 & N1415;
  assign N9460 = N9248 & idx_w_i[8];
  assign N9461 = N9249 & N1415;
  assign N9462 = N9249 & idx_w_i[8];
  assign N9463 = N9250 & N1415;
  assign N9464 = N9250 & idx_w_i[8];
  assign N9465 = N9251 & N1415;
  assign N9466 = N9251 & idx_w_i[8];
  assign N9467 = N9252 & N1415;
  assign N9468 = N9252 & idx_w_i[8];
  assign N9469 = N9253 & N1415;
  assign N9470 = N9253 & idx_w_i[8];
  assign N9471 = N9254 & N1415;
  assign N9472 = N9254 & idx_w_i[8];
  assign N9473 = N9255 & N1415;
  assign N9474 = N9255 & idx_w_i[8];
  assign N9475 = N9256 & N1415;
  assign N9476 = N9256 & idx_w_i[8];
  assign N9477 = N9257 & N1415;
  assign N9478 = N9257 & idx_w_i[8];
  assign N9479 = N9258 & N1415;
  assign N9480 = N9258 & idx_w_i[8];
  assign N9481 = N9259 & N1415;
  assign N9482 = N9259 & idx_w_i[8];
  assign N9483 = N9260 & N1415;
  assign N9484 = N9260 & idx_w_i[8];
  assign N9485 = N9261 & N1415;
  assign N9486 = N9261 & idx_w_i[8];
  assign N9487 = N9262 & N1415;
  assign N9488 = N9262 & idx_w_i[8];
  assign N9489 = N9263 & N1415;
  assign N9490 = N9263 & idx_w_i[8];
  assign N9491 = N9264 & N1415;
  assign N9492 = N9264 & idx_w_i[8];
  assign N9493 = N9265 & N1415;
  assign N9494 = N9265 & idx_w_i[8];
  assign N9495 = N9266 & N1415;
  assign N9496 = N9266 & idx_w_i[8];
  assign N9497 = N9267 & N1415;
  assign N9498 = N9267 & idx_w_i[8];
  assign N9499 = N9268 & N1415;
  assign N9500 = N9268 & idx_w_i[8];
  assign N9501 = N9269 & N1415;
  assign N9502 = N9269 & idx_w_i[8];
  assign N9503 = N9270 & N1415;
  assign N9504 = N9270 & idx_w_i[8];
  assign N9505 = N9271 & N1415;
  assign N9506 = N9271 & idx_w_i[8];
  assign N9507 = N9272 & N1415;
  assign N9508 = N9272 & idx_w_i[8];
  assign N9509 = N9273 & N1415;
  assign N9510 = N9273 & idx_w_i[8];
  assign N9511 = N9274 & N1415;
  assign N9512 = N9274 & idx_w_i[8];
  assign N9513 = N9275 & N1415;
  assign N9514 = N9275 & idx_w_i[8];
  assign N9515 = N9276 & N1415;
  assign N9516 = N9276 & idx_w_i[8];
  assign N9517 = N9277 & N1415;
  assign N9518 = N9277 & idx_w_i[8];
  assign N9519 = N9278 & N1415;
  assign N9520 = N9278 & idx_w_i[8];
  assign N9521 = N9279 & N1415;
  assign N9522 = N9279 & idx_w_i[8];
  assign N9523 = N9280 & N1415;
  assign N9524 = N9280 & idx_w_i[8];
  assign N9525 = N9281 & N1415;
  assign N9526 = N9281 & idx_w_i[8];
  assign N9527 = N9282 & N1415;
  assign N9528 = N9282 & idx_w_i[8];
  assign N9529 = N9283 & N1415;
  assign N9530 = N9283 & idx_w_i[8];
  assign N9531 = N9284 & N1415;
  assign N9532 = N9284 & idx_w_i[8];
  assign N9533 = N9285 & N1415;
  assign N9534 = N9285 & idx_w_i[8];
  assign N9535 = N9286 & N1415;
  assign N9536 = N9286 & idx_w_i[8];
  assign N9537 = N9287 & N1415;
  assign N9538 = N9287 & idx_w_i[8];
  assign N9539 = N9288 & N1415;
  assign N9540 = N9288 & idx_w_i[8];
  assign N9541 = N9289 & N1415;
  assign N9542 = N9289 & idx_w_i[8];
  assign N9543 = N9290 & N1415;
  assign N9544 = N9290 & idx_w_i[8];
  assign N9545 = N9291 & N1415;
  assign N9546 = N9291 & idx_w_i[8];
  assign N9547 = N9292 & N1415;
  assign N9548 = N9292 & idx_w_i[8];
  assign N9549 = N9102 & N1415;
  assign N9550 = N9102 & idx_w_i[8];
  assign N9551 = N9104 & N1415;
  assign N9552 = N9104 & idx_w_i[8];
  assign N9553 = N9106 & N1415;
  assign N9554 = N9106 & idx_w_i[8];
  assign N9555 = N9108 & N1415;
  assign N9556 = N9108 & idx_w_i[8];
  assign N9557 = N9110 & N1415;
  assign N9558 = N9110 & idx_w_i[8];
  assign N9559 = N9112 & N1415;
  assign N9560 = N9112 & idx_w_i[8];
  assign N9561 = N9114 & N1415;
  assign N9562 = N9114 & idx_w_i[8];
  assign N9563 = N9116 & N1415;
  assign N9564 = N9116 & idx_w_i[8];
  assign N9565 = N9118 & N1415;
  assign N9566 = N9118 & idx_w_i[8];
  assign N9567 = N9120 & N1415;
  assign N9568 = N9120 & idx_w_i[8];
  assign N9569 = N9122 & N1415;
  assign N9570 = N9122 & idx_w_i[8];
  assign N9571 = N9124 & N1415;
  assign N9572 = N9124 & idx_w_i[8];
  assign N9573 = N9126 & N1415;
  assign N9574 = N9126 & idx_w_i[8];
  assign N9575 = N9128 & N1415;
  assign N9576 = N9128 & idx_w_i[8];
  assign N9577 = N9130 & N1415;
  assign N9578 = N9130 & idx_w_i[8];
  assign N9579 = N9132 & N1415;
  assign N9580 = N9132 & idx_w_i[8];
  assign N9581 = N9134 & N1415;
  assign N9582 = N9134 & idx_w_i[8];
  assign N9583 = N9136 & N1415;
  assign N9584 = N9136 & idx_w_i[8];
  assign N9585 = N9138 & N1415;
  assign N9586 = N9138 & idx_w_i[8];
  assign N9587 = N9140 & N1415;
  assign N9588 = N9140 & idx_w_i[8];
  assign N9589 = N9142 & N1415;
  assign N9590 = N9142 & idx_w_i[8];
  assign N9591 = N9144 & N1415;
  assign N9592 = N9144 & idx_w_i[8];
  assign N9593 = N9146 & N1415;
  assign N9594 = N9146 & idx_w_i[8];
  assign N9595 = N9148 & N1415;
  assign N9596 = N9148 & idx_w_i[8];
  assign N9597 = N9150 & N1415;
  assign N9598 = N9150 & idx_w_i[8];
  assign N9599 = N9152 & N1415;
  assign N9600 = N9152 & idx_w_i[8];
  assign N9601 = N9154 & N1415;
  assign N9602 = N9154 & idx_w_i[8];
  assign N9603 = N9156 & N1415;
  assign N9604 = N9156 & idx_w_i[8];
  assign N9605 = N9158 & N1415;
  assign N9606 = N9158 & idx_w_i[8];
  assign N9607 = N9160 & N1415;
  assign N9608 = N9160 & idx_w_i[8];
  assign N9609 = N9162 & N1415;
  assign N9610 = N9162 & idx_w_i[8];
  assign N9611 = N9164 & N1415;
  assign N9612 = N9164 & idx_w_i[8];
  assign N9613 = N9166 & N1415;
  assign N9614 = N9166 & idx_w_i[8];
  assign N9615 = N9168 & N1415;
  assign N9616 = N9168 & idx_w_i[8];
  assign N9617 = N9170 & N1415;
  assign N9618 = N9170 & idx_w_i[8];
  assign N9619 = N9172 & N1415;
  assign N9620 = N9172 & idx_w_i[8];
  assign N9621 = N9174 & N1415;
  assign N9622 = N9174 & idx_w_i[8];
  assign N9623 = N9176 & N1415;
  assign N9624 = N9176 & idx_w_i[8];
  assign N9625 = N9178 & N1415;
  assign N9626 = N9178 & idx_w_i[8];
  assign N9627 = N9180 & N1415;
  assign N9628 = N9180 & idx_w_i[8];
  assign N9629 = N9182 & N1415;
  assign N9630 = N9182 & idx_w_i[8];
  assign N9631 = N9184 & N1415;
  assign N9632 = N9184 & idx_w_i[8];
  assign N9633 = N9186 & N1415;
  assign N9634 = N9186 & idx_w_i[8];
  assign N9635 = N9188 & N1415;
  assign N9636 = N9188 & idx_w_i[8];
  assign N9637 = N9190 & N1415;
  assign N9638 = N9190 & idx_w_i[8];
  assign N9639 = N9192 & N1415;
  assign N9640 = N9192 & idx_w_i[8];
  assign N9641 = N9194 & N1415;
  assign N9642 = N9194 & idx_w_i[8];
  assign N9643 = N9196 & N1415;
  assign N9644 = N9196 & idx_w_i[8];
  assign N9645 = N9198 & N1415;
  assign N9646 = N9198 & idx_w_i[8];
  assign N9647 = N9200 & N1415;
  assign N9648 = N9200 & idx_w_i[8];
  assign N9649 = N9202 & N1415;
  assign N9650 = N9202 & idx_w_i[8];
  assign N9651 = N9204 & N1415;
  assign N9652 = N9204 & idx_w_i[8];
  assign N9653 = N9206 & N1415;
  assign N9654 = N9206 & idx_w_i[8];
  assign N9655 = N9208 & N1415;
  assign N9656 = N9208 & idx_w_i[8];
  assign N9657 = N9210 & N1415;
  assign N9658 = N9210 & idx_w_i[8];
  assign N9659 = N9212 & N1415;
  assign N9660 = N9212 & idx_w_i[8];
  assign N9661 = N9214 & N1415;
  assign N9662 = N9214 & idx_w_i[8];
  assign N9663 = N9216 & N1415;
  assign N9664 = N9216 & idx_w_i[8];
  assign N9665 = N9218 & N1415;
  assign N9666 = N9218 & idx_w_i[8];
  assign N9667 = N9220 & N1415;
  assign N9668 = N9220 & idx_w_i[8];
  assign N9669 = N9222 & N1415;
  assign N9670 = N9222 & idx_w_i[8];
  assign N9671 = N9224 & N1415;
  assign N9672 = N9224 & idx_w_i[8];
  assign N9673 = N9226 & N1415;
  assign N9674 = N9226 & idx_w_i[8];
  assign N9675 = N9228 & N1415;
  assign N9676 = N9228 & idx_w_i[8];
  assign N9677 = N8493 & N1415;
  assign N9678 = N8495 & N1415;
  assign N9679 = N8497 & N1415;
  assign N9680 = N8499 & N1415;
  assign N9681 = N8501 & N1415;
  assign N9682 = N8503 & N1415;
  assign N9683 = N8505 & N1415;
  assign N9684 = N8507 & N1415;
  assign N9685 = N3044 & N1415;
  assign N9686 = N3046 & N1415;
  assign N9687 = N3048 & N1415;
  assign N9688 = N3050 & N1415;
  assign N9689 = N3052 & N1415;
  assign N9690 = N3054 & N1415;
  assign N9691 = N3056 & N1415;
  assign N9692 = N3058 & N1415;
  assign N9693 = N8517 & N1415;
  assign N9694 = N8519 & N1415;
  assign N9695 = N8521 & N1415;
  assign N9696 = N8523 & N1415;
  assign N9697 = N8525 & N1415;
  assign N9698 = N8527 & N1415;
  assign N9699 = N8529 & N1415;
  assign N9700 = N8531 & N1415;
  assign N9701 = N3076 & N1415;
  assign N9702 = N3078 & N1415;
  assign N9703 = N3080 & N1415;
  assign N9704 = N3082 & N1415;
  assign N9705 = N3084 & N1415;
  assign N9706 = N3086 & N1415;
  assign N9707 = N3088 & N1415;
  assign N9708 = N3090 & N1415;
  assign N9709 = N6248 & N1415;
  assign N9710 = N6250 & N1415;
  assign N9711 = N6252 & N1415;
  assign N9712 = N6254 & N1415;
  assign N9713 = N6256 & N1415;
  assign N9714 = N6258 & N1415;
  assign N9715 = N6260 & N1415;
  assign N9716 = N6262 & N1415;
  assign N9717 = N3108 & N1415;
  assign N9718 = N3110 & N1415;
  assign N9719 = N3112 & N1415;
  assign N9720 = N3114 & N1415;
  assign N9721 = N3116 & N1415;
  assign N9722 = N3118 & N1415;
  assign N9723 = N3120 & N1415;
  assign N9724 = N3122 & N1415;
  assign N9725 = N11569 & N1415;
  assign N9726 = N11571 & N1415;
  assign N9727 = N11573 & N1415;
  assign N9728 = N11575 & N1415;
  assign N9729 = N11577 & N1415;
  assign N9730 = N11579 & N1415;
  assign N9731 = N11581 & N1415;
  assign N9732 = N11583 & N1415;
  assign N9733 = N11585 & N1415;
  assign N9734 = N11587 & N1415;
  assign N9735 = N11589 & N1415;
  assign N9736 = N11591 & N1415;
  assign N9737 = N11593 & N1415;
  assign N9738 = N11595 & N1415;
  assign N9739 = N11597 & N1415;
  assign N9740 = N11599 & N1415;
  assign N10254 = N9036 ^ N9741;
  assign N10255 = N11120 & N1060;
  assign N10256 = N11122 & N1060;
  assign N10257 = N11124 & N1060;
  assign N10258 = N11126 & N1060;
  assign N10259 = N11128 & N1060;
  assign N10260 = N11130 & N1060;
  assign N10261 = N11132 & N1060;
  assign N10262 = N11134 & N1060;
  assign N10263 = N11136 & N1060;
  assign N10264 = N11138 & N1060;
  assign N10265 = N11140 & N1060;
  assign N10266 = N11142 & N1060;
  assign N10267 = N11144 & N1060;
  assign N10268 = N11146 & N1060;
  assign N10269 = N11148 & N1060;
  assign N10270 = N11150 & N1060;
  assign N10271 = N11121 & N1060;
  assign N10272 = N11123 & N1060;
  assign N10273 = N11125 & N1060;
  assign N10274 = N11127 & N1060;
  assign N10275 = N11129 & N1060;
  assign N10276 = N11131 & N1060;
  assign N10277 = N11133 & N1060;
  assign N10278 = N11135 & N1060;
  assign N10279 = N11137 & N1060;
  assign N10280 = N11139 & N1060;
  assign N10281 = N11141 & N1060;
  assign N10282 = N11143 & N1060;
  assign N10283 = N11145 & N1060;
  assign N10284 = N11147 & N1060;
  assign N10285 = N11149 & N1060;
  assign N10286 = N11151 & N1060;
  assign N10287 = N10255 & N1093;
  assign N10288 = N10255 & idx_w_i[6];
  assign N10289 = N10256 & N1093;
  assign N10290 = N10256 & idx_w_i[6];
  assign N10291 = N10257 & N1093;
  assign N10292 = N10257 & idx_w_i[6];
  assign N10293 = N10258 & N1093;
  assign N10294 = N10258 & idx_w_i[6];
  assign N10295 = N10259 & N1093;
  assign N10296 = N10259 & idx_w_i[6];
  assign N10297 = N10260 & N1093;
  assign N10298 = N10260 & idx_w_i[6];
  assign N10299 = N10261 & N1093;
  assign N10300 = N10261 & idx_w_i[6];
  assign N10301 = N10262 & N1093;
  assign N10302 = N10262 & idx_w_i[6];
  assign N10303 = N10263 & N1093;
  assign N10304 = N10263 & idx_w_i[6];
  assign N10305 = N10264 & N1093;
  assign N10306 = N10264 & idx_w_i[6];
  assign N10307 = N10265 & N1093;
  assign N10308 = N10265 & idx_w_i[6];
  assign N10309 = N10266 & N1093;
  assign N10310 = N10266 & idx_w_i[6];
  assign N10311 = N10267 & N1093;
  assign N10312 = N10267 & idx_w_i[6];
  assign N10313 = N10268 & N1093;
  assign N10314 = N10268 & idx_w_i[6];
  assign N10315 = N10269 & N1093;
  assign N10316 = N10269 & idx_w_i[6];
  assign N10317 = N10270 & N1093;
  assign N10318 = N10270 & idx_w_i[6];
  assign N10319 = N10271 & N1093;
  assign N10320 = N10271 & idx_w_i[6];
  assign N10321 = N10272 & N1093;
  assign N10322 = N10272 & idx_w_i[6];
  assign N10323 = N10273 & N1093;
  assign N10324 = N10273 & idx_w_i[6];
  assign N10325 = N10274 & N1093;
  assign N10326 = N10274 & idx_w_i[6];
  assign N10327 = N10275 & N1093;
  assign N10328 = N10275 & idx_w_i[6];
  assign N10329 = N10276 & N1093;
  assign N10330 = N10276 & idx_w_i[6];
  assign N10331 = N10277 & N1093;
  assign N10332 = N10277 & idx_w_i[6];
  assign N10333 = N10278 & N1093;
  assign N10334 = N10278 & idx_w_i[6];
  assign N10335 = N10279 & N1093;
  assign N10336 = N10279 & idx_w_i[6];
  assign N10337 = N10280 & N1093;
  assign N10338 = N10280 & idx_w_i[6];
  assign N10339 = N10281 & N1093;
  assign N10340 = N10281 & idx_w_i[6];
  assign N10341 = N10282 & N1093;
  assign N10342 = N10282 & idx_w_i[6];
  assign N10343 = N10283 & N1093;
  assign N10344 = N10283 & idx_w_i[6];
  assign N10345 = N10284 & N1093;
  assign N10346 = N10284 & idx_w_i[6];
  assign N10347 = N10285 & N1093;
  assign N10348 = N10285 & idx_w_i[6];
  assign N10349 = N10286 & N1093;
  assign N10350 = N10286 & idx_w_i[6];
  assign N10351 = N11153 & N1093;
  assign N10352 = N11155 & N1093;
  assign N10353 = N11157 & N1093;
  assign N10354 = N11159 & N1093;
  assign N10355 = N11161 & N1093;
  assign N10356 = N11163 & N1093;
  assign N10357 = N11165 & N1093;
  assign N10358 = N11167 & N1093;
  assign N10359 = N11169 & N1093;
  assign N10360 = N11171 & N1093;
  assign N10361 = N11173 & N1093;
  assign N10362 = N11175 & N1093;
  assign N10363 = N11177 & N1093;
  assign N10364 = N11179 & N1093;
  assign N10365 = N11181 & N1093;
  assign N10366 = N11183 & N1093;
  assign N10367 = N11185 & N1093;
  assign N10368 = N11187 & N1093;
  assign N10369 = N11189 & N1093;
  assign N10370 = N11191 & N1093;
  assign N10371 = N11193 & N1093;
  assign N10372 = N11195 & N1093;
  assign N10373 = N11197 & N1093;
  assign N10374 = N11199 & N1093;
  assign N10375 = N11201 & N1093;
  assign N10376 = N11203 & N1093;
  assign N10377 = N11205 & N1093;
  assign N10378 = N11207 & N1093;
  assign N10379 = N11209 & N1093;
  assign N10380 = N11211 & N1093;
  assign N10381 = N11213 & N1093;
  assign N10382 = N11215 & N1093;
  assign N10383 = N10287 & N1190;
  assign N10384 = N10287 & idx_w_i[7];
  assign N10385 = N10289 & N1190;
  assign N10386 = N10289 & idx_w_i[7];
  assign N10387 = N10291 & N1190;
  assign N10388 = N10291 & idx_w_i[7];
  assign N10389 = N10293 & N1190;
  assign N10390 = N10293 & idx_w_i[7];
  assign N10391 = N10295 & N1190;
  assign N10392 = N10295 & idx_w_i[7];
  assign N10393 = N10297 & N1190;
  assign N10394 = N10297 & idx_w_i[7];
  assign N10395 = N10299 & N1190;
  assign N10396 = N10299 & idx_w_i[7];
  assign N10397 = N10301 & N1190;
  assign N10398 = N10301 & idx_w_i[7];
  assign N10399 = N10303 & N1190;
  assign N10400 = N10303 & idx_w_i[7];
  assign N10401 = N10305 & N1190;
  assign N10402 = N10305 & idx_w_i[7];
  assign N10403 = N10307 & N1190;
  assign N10404 = N10307 & idx_w_i[7];
  assign N10405 = N10309 & N1190;
  assign N10406 = N10309 & idx_w_i[7];
  assign N10407 = N10311 & N1190;
  assign N10408 = N10311 & idx_w_i[7];
  assign N10409 = N10313 & N1190;
  assign N10410 = N10313 & idx_w_i[7];
  assign N10411 = N10315 & N1190;
  assign N10412 = N10315 & idx_w_i[7];
  assign N10413 = N10317 & N1190;
  assign N10414 = N10317 & idx_w_i[7];
  assign N10415 = N10319 & N1190;
  assign N10416 = N10319 & idx_w_i[7];
  assign N10417 = N10321 & N1190;
  assign N10418 = N10321 & idx_w_i[7];
  assign N10419 = N10323 & N1190;
  assign N10420 = N10323 & idx_w_i[7];
  assign N10421 = N10325 & N1190;
  assign N10422 = N10325 & idx_w_i[7];
  assign N10423 = N10327 & N1190;
  assign N10424 = N10327 & idx_w_i[7];
  assign N10425 = N10329 & N1190;
  assign N10426 = N10329 & idx_w_i[7];
  assign N10427 = N10331 & N1190;
  assign N10428 = N10331 & idx_w_i[7];
  assign N10429 = N10333 & N1190;
  assign N10430 = N10333 & idx_w_i[7];
  assign N10431 = N10335 & N1190;
  assign N10432 = N10335 & idx_w_i[7];
  assign N10433 = N10337 & N1190;
  assign N10434 = N10337 & idx_w_i[7];
  assign N10435 = N10339 & N1190;
  assign N10436 = N10339 & idx_w_i[7];
  assign N10437 = N10341 & N1190;
  assign N10438 = N10341 & idx_w_i[7];
  assign N10439 = N10343 & N1190;
  assign N10440 = N10343 & idx_w_i[7];
  assign N10441 = N10345 & N1190;
  assign N10442 = N10345 & idx_w_i[7];
  assign N10443 = N10347 & N1190;
  assign N10444 = N10347 & idx_w_i[7];
  assign N10445 = N10349 & N1190;
  assign N10446 = N10349 & idx_w_i[7];
  assign N10447 = N10351 & N1190;
  assign N10448 = N10351 & idx_w_i[7];
  assign N10449 = N10352 & N1190;
  assign N10450 = N10352 & idx_w_i[7];
  assign N10451 = N10353 & N1190;
  assign N10452 = N10353 & idx_w_i[7];
  assign N10453 = N10354 & N1190;
  assign N10454 = N10354 & idx_w_i[7];
  assign N10455 = N10355 & N1190;
  assign N10456 = N10355 & idx_w_i[7];
  assign N10457 = N10356 & N1190;
  assign N10458 = N10356 & idx_w_i[7];
  assign N10459 = N10357 & N1190;
  assign N10460 = N10357 & idx_w_i[7];
  assign N10461 = N10358 & N1190;
  assign N10462 = N10358 & idx_w_i[7];
  assign N10463 = N10359 & N1190;
  assign N10464 = N10359 & idx_w_i[7];
  assign N10465 = N10360 & N1190;
  assign N10466 = N10360 & idx_w_i[7];
  assign N10467 = N10361 & N1190;
  assign N10468 = N10361 & idx_w_i[7];
  assign N10469 = N10362 & N1190;
  assign N10470 = N10362 & idx_w_i[7];
  assign N10471 = N10363 & N1190;
  assign N10472 = N10363 & idx_w_i[7];
  assign N10473 = N10364 & N1190;
  assign N10474 = N10364 & idx_w_i[7];
  assign N10475 = N10365 & N1190;
  assign N10476 = N10365 & idx_w_i[7];
  assign N10477 = N10366 & N1190;
  assign N10478 = N10366 & idx_w_i[7];
  assign N10479 = N10367 & N1190;
  assign N10480 = N10367 & idx_w_i[7];
  assign N10481 = N10368 & N1190;
  assign N10482 = N10368 & idx_w_i[7];
  assign N10483 = N10369 & N1190;
  assign N10484 = N10369 & idx_w_i[7];
  assign N10485 = N10370 & N1190;
  assign N10486 = N10370 & idx_w_i[7];
  assign N10487 = N10371 & N1190;
  assign N10488 = N10371 & idx_w_i[7];
  assign N10489 = N10372 & N1190;
  assign N10490 = N10372 & idx_w_i[7];
  assign N10491 = N10373 & N1190;
  assign N10492 = N10373 & idx_w_i[7];
  assign N10493 = N10374 & N1190;
  assign N10494 = N10374 & idx_w_i[7];
  assign N10495 = N10375 & N1190;
  assign N10496 = N10375 & idx_w_i[7];
  assign N10497 = N10376 & N1190;
  assign N10498 = N10376 & idx_w_i[7];
  assign N10499 = N10377 & N1190;
  assign N10500 = N10377 & idx_w_i[7];
  assign N10501 = N10378 & N1190;
  assign N10502 = N10378 & idx_w_i[7];
  assign N10503 = N10379 & N1190;
  assign N10504 = N10379 & idx_w_i[7];
  assign N10505 = N10380 & N1190;
  assign N10506 = N10380 & idx_w_i[7];
  assign N10507 = N10381 & N1190;
  assign N10508 = N10381 & idx_w_i[7];
  assign N10509 = N10382 & N1190;
  assign N10510 = N10382 & idx_w_i[7];
  assign N10511 = N10288 & N1190;
  assign N10512 = N10288 & idx_w_i[7];
  assign N10513 = N10290 & N1190;
  assign N10514 = N10290 & idx_w_i[7];
  assign N10515 = N10292 & N1190;
  assign N10516 = N10292 & idx_w_i[7];
  assign N10517 = N10294 & N1190;
  assign N10518 = N10294 & idx_w_i[7];
  assign N10519 = N10296 & N1190;
  assign N10520 = N10296 & idx_w_i[7];
  assign N10521 = N10298 & N1190;
  assign N10522 = N10298 & idx_w_i[7];
  assign N10523 = N10300 & N1190;
  assign N10524 = N10300 & idx_w_i[7];
  assign N10525 = N10302 & N1190;
  assign N10526 = N10302 & idx_w_i[7];
  assign N10527 = N10304 & N1190;
  assign N10528 = N10304 & idx_w_i[7];
  assign N10529 = N10306 & N1190;
  assign N10530 = N10306 & idx_w_i[7];
  assign N10531 = N10308 & N1190;
  assign N10532 = N10308 & idx_w_i[7];
  assign N10533 = N10310 & N1190;
  assign N10534 = N10310 & idx_w_i[7];
  assign N10535 = N10312 & N1190;
  assign N10536 = N10312 & idx_w_i[7];
  assign N10537 = N10314 & N1190;
  assign N10538 = N10314 & idx_w_i[7];
  assign N10539 = N10316 & N1190;
  assign N10540 = N10316 & idx_w_i[7];
  assign N10541 = N10318 & N1190;
  assign N10542 = N10318 & idx_w_i[7];
  assign N10543 = N10320 & N1190;
  assign N10544 = N10320 & idx_w_i[7];
  assign N10545 = N10322 & N1190;
  assign N10546 = N10322 & idx_w_i[7];
  assign N10547 = N10324 & N1190;
  assign N10548 = N10324 & idx_w_i[7];
  assign N10549 = N10326 & N1190;
  assign N10550 = N10326 & idx_w_i[7];
  assign N10551 = N10328 & N1190;
  assign N10552 = N10328 & idx_w_i[7];
  assign N10553 = N10330 & N1190;
  assign N10554 = N10330 & idx_w_i[7];
  assign N10555 = N10332 & N1190;
  assign N10556 = N10332 & idx_w_i[7];
  assign N10557 = N10334 & N1190;
  assign N10558 = N10334 & idx_w_i[7];
  assign N10559 = N10336 & N1190;
  assign N10560 = N10336 & idx_w_i[7];
  assign N10561 = N10338 & N1190;
  assign N10562 = N10338 & idx_w_i[7];
  assign N10563 = N10340 & N1190;
  assign N10564 = N10340 & idx_w_i[7];
  assign N10565 = N10342 & N1190;
  assign N10566 = N10342 & idx_w_i[7];
  assign N10567 = N10344 & N1190;
  assign N10568 = N10344 & idx_w_i[7];
  assign N10569 = N10346 & N1190;
  assign N10570 = N10346 & idx_w_i[7];
  assign N10571 = N10348 & N1190;
  assign N10572 = N10348 & idx_w_i[7];
  assign N10573 = N10350 & N1190;
  assign N10574 = N10350 & idx_w_i[7];
  assign N10575 = N11281 & N1190;
  assign N10576 = N11283 & N1190;
  assign N10577 = N11285 & N1190;
  assign N10578 = N11287 & N1190;
  assign N10579 = N11289 & N1190;
  assign N10580 = N11291 & N1190;
  assign N10581 = N11293 & N1190;
  assign N10582 = N11295 & N1190;
  assign N10583 = N11297 & N1190;
  assign N10584 = N11299 & N1190;
  assign N10585 = N11301 & N1190;
  assign N10586 = N11303 & N1190;
  assign N10587 = N11305 & N1190;
  assign N10588 = N11307 & N1190;
  assign N10589 = N11309 & N1190;
  assign N10590 = N11311 & N1190;
  assign N10591 = N11313 & N1190;
  assign N10592 = N11315 & N1190;
  assign N10593 = N11317 & N1190;
  assign N10594 = N11319 & N1190;
  assign N10595 = N11321 & N1190;
  assign N10596 = N11323 & N1190;
  assign N10597 = N11325 & N1190;
  assign N10598 = N11327 & N1190;
  assign N10599 = N11329 & N1190;
  assign N10600 = N11331 & N1190;
  assign N10601 = N11333 & N1190;
  assign N10602 = N11335 & N1190;
  assign N10603 = N11337 & N1190;
  assign N10604 = N11339 & N1190;
  assign N10605 = N11341 & N1190;
  assign N10606 = N11343 & N1190;
  assign N10607 = N10383 & N1415;
  assign N10608 = N10383 & idx_w_i[8];
  assign N10609 = N10385 & N1415;
  assign N10610 = N10385 & idx_w_i[8];
  assign N10611 = N10387 & N1415;
  assign N10612 = N10387 & idx_w_i[8];
  assign N10613 = N10389 & N1415;
  assign N10614 = N10389 & idx_w_i[8];
  assign N10615 = N10391 & N1415;
  assign N10616 = N10391 & idx_w_i[8];
  assign N10617 = N10393 & N1415;
  assign N10618 = N10393 & idx_w_i[8];
  assign N10619 = N10395 & N1415;
  assign N10620 = N10395 & idx_w_i[8];
  assign N10621 = N10397 & N1415;
  assign N10622 = N10397 & idx_w_i[8];
  assign N10623 = N10399 & N1415;
  assign N10624 = N10399 & idx_w_i[8];
  assign N10625 = N10401 & N1415;
  assign N10626 = N10401 & idx_w_i[8];
  assign N10627 = N10403 & N1415;
  assign N10628 = N10403 & idx_w_i[8];
  assign N10629 = N10405 & N1415;
  assign N10630 = N10405 & idx_w_i[8];
  assign N10631 = N10407 & N1415;
  assign N10632 = N10407 & idx_w_i[8];
  assign N10633 = N10409 & N1415;
  assign N10634 = N10409 & idx_w_i[8];
  assign N10635 = N10411 & N1415;
  assign N10636 = N10411 & idx_w_i[8];
  assign N10637 = N10413 & N1415;
  assign N10638 = N10413 & idx_w_i[8];
  assign N10639 = N10415 & N1415;
  assign N10640 = N10415 & idx_w_i[8];
  assign N10641 = N10417 & N1415;
  assign N10642 = N10417 & idx_w_i[8];
  assign N10643 = N10419 & N1415;
  assign N10644 = N10419 & idx_w_i[8];
  assign N10645 = N10421 & N1415;
  assign N10646 = N10421 & idx_w_i[8];
  assign N10647 = N10423 & N1415;
  assign N10648 = N10423 & idx_w_i[8];
  assign N10649 = N10425 & N1415;
  assign N10650 = N10425 & idx_w_i[8];
  assign N10651 = N10427 & N1415;
  assign N10652 = N10427 & idx_w_i[8];
  assign N10653 = N10429 & N1415;
  assign N10654 = N10429 & idx_w_i[8];
  assign N10655 = N10431 & N1415;
  assign N10656 = N10431 & idx_w_i[8];
  assign N10657 = N10433 & N1415;
  assign N10658 = N10433 & idx_w_i[8];
  assign N10659 = N10435 & N1415;
  assign N10660 = N10435 & idx_w_i[8];
  assign N10661 = N10437 & N1415;
  assign N10662 = N10437 & idx_w_i[8];
  assign N10663 = N10439 & N1415;
  assign N10664 = N10439 & idx_w_i[8];
  assign N10665 = N10441 & N1415;
  assign N10666 = N10441 & idx_w_i[8];
  assign N10667 = N10443 & N1415;
  assign N10668 = N10443 & idx_w_i[8];
  assign N10669 = N10445 & N1415;
  assign N10670 = N10445 & idx_w_i[8];
  assign N10671 = N10447 & N1415;
  assign N10672 = N10447 & idx_w_i[8];
  assign N10673 = N10449 & N1415;
  assign N10674 = N10449 & idx_w_i[8];
  assign N10675 = N10451 & N1415;
  assign N10676 = N10451 & idx_w_i[8];
  assign N10677 = N10453 & N1415;
  assign N10678 = N10453 & idx_w_i[8];
  assign N10679 = N10455 & N1415;
  assign N10680 = N10455 & idx_w_i[8];
  assign N10681 = N10457 & N1415;
  assign N10682 = N10457 & idx_w_i[8];
  assign N10683 = N10459 & N1415;
  assign N10684 = N10459 & idx_w_i[8];
  assign N10685 = N10461 & N1415;
  assign N10686 = N10461 & idx_w_i[8];
  assign N10687 = N10463 & N1415;
  assign N10688 = N10463 & idx_w_i[8];
  assign N10689 = N10465 & N1415;
  assign N10690 = N10465 & idx_w_i[8];
  assign N10691 = N10467 & N1415;
  assign N10692 = N10467 & idx_w_i[8];
  assign N10693 = N10469 & N1415;
  assign N10694 = N10469 & idx_w_i[8];
  assign N10695 = N10471 & N1415;
  assign N10696 = N10471 & idx_w_i[8];
  assign N10697 = N10473 & N1415;
  assign N10698 = N10473 & idx_w_i[8];
  assign N10699 = N10475 & N1415;
  assign N10700 = N10475 & idx_w_i[8];
  assign N10701 = N10477 & N1415;
  assign N10702 = N10477 & idx_w_i[8];
  assign N10703 = N10479 & N1415;
  assign N10704 = N10479 & idx_w_i[8];
  assign N10705 = N10481 & N1415;
  assign N10706 = N10481 & idx_w_i[8];
  assign N10707 = N10483 & N1415;
  assign N10708 = N10483 & idx_w_i[8];
  assign N10709 = N10485 & N1415;
  assign N10710 = N10485 & idx_w_i[8];
  assign N10711 = N10487 & N1415;
  assign N10712 = N10487 & idx_w_i[8];
  assign N10713 = N10489 & N1415;
  assign N10714 = N10489 & idx_w_i[8];
  assign N10715 = N10491 & N1415;
  assign N10716 = N10491 & idx_w_i[8];
  assign N10717 = N10493 & N1415;
  assign N10718 = N10493 & idx_w_i[8];
  assign N10719 = N10495 & N1415;
  assign N10720 = N10495 & idx_w_i[8];
  assign N10721 = N10497 & N1415;
  assign N10722 = N10497 & idx_w_i[8];
  assign N10723 = N10499 & N1415;
  assign N10724 = N10499 & idx_w_i[8];
  assign N10725 = N10501 & N1415;
  assign N10726 = N10501 & idx_w_i[8];
  assign N10727 = N10503 & N1415;
  assign N10728 = N10503 & idx_w_i[8];
  assign N10729 = N10505 & N1415;
  assign N10730 = N10505 & idx_w_i[8];
  assign N10731 = N10507 & N1415;
  assign N10732 = N10507 & idx_w_i[8];
  assign N10733 = N10509 & N1415;
  assign N10734 = N10509 & idx_w_i[8];
  assign N10735 = N10511 & N1415;
  assign N10736 = N10511 & idx_w_i[8];
  assign N10737 = N10513 & N1415;
  assign N10738 = N10513 & idx_w_i[8];
  assign N10739 = N10515 & N1415;
  assign N10740 = N10515 & idx_w_i[8];
  assign N10741 = N10517 & N1415;
  assign N10742 = N10517 & idx_w_i[8];
  assign N10743 = N10519 & N1415;
  assign N10744 = N10519 & idx_w_i[8];
  assign N10745 = N10521 & N1415;
  assign N10746 = N10521 & idx_w_i[8];
  assign N10747 = N10523 & N1415;
  assign N10748 = N10523 & idx_w_i[8];
  assign N10749 = N10525 & N1415;
  assign N10750 = N10525 & idx_w_i[8];
  assign N10751 = N10527 & N1415;
  assign N10752 = N10527 & idx_w_i[8];
  assign N10753 = N10529 & N1415;
  assign N10754 = N10529 & idx_w_i[8];
  assign N10755 = N10531 & N1415;
  assign N10756 = N10531 & idx_w_i[8];
  assign N10757 = N10533 & N1415;
  assign N10758 = N10533 & idx_w_i[8];
  assign N10759 = N10535 & N1415;
  assign N10760 = N10535 & idx_w_i[8];
  assign N10761 = N10537 & N1415;
  assign N10762 = N10537 & idx_w_i[8];
  assign N10763 = N10539 & N1415;
  assign N10764 = N10539 & idx_w_i[8];
  assign N10765 = N10541 & N1415;
  assign N10766 = N10541 & idx_w_i[8];
  assign N10767 = N10543 & N1415;
  assign N10768 = N10543 & idx_w_i[8];
  assign N10769 = N10545 & N1415;
  assign N10770 = N10545 & idx_w_i[8];
  assign N10771 = N10547 & N1415;
  assign N10772 = N10547 & idx_w_i[8];
  assign N10773 = N10549 & N1415;
  assign N10774 = N10549 & idx_w_i[8];
  assign N10775 = N10551 & N1415;
  assign N10776 = N10551 & idx_w_i[8];
  assign N10777 = N10553 & N1415;
  assign N10778 = N10553 & idx_w_i[8];
  assign N10779 = N10555 & N1415;
  assign N10780 = N10555 & idx_w_i[8];
  assign N10781 = N10557 & N1415;
  assign N10782 = N10557 & idx_w_i[8];
  assign N10783 = N10559 & N1415;
  assign N10784 = N10559 & idx_w_i[8];
  assign N10785 = N10561 & N1415;
  assign N10786 = N10561 & idx_w_i[8];
  assign N10787 = N10563 & N1415;
  assign N10788 = N10563 & idx_w_i[8];
  assign N10789 = N10565 & N1415;
  assign N10790 = N10565 & idx_w_i[8];
  assign N10791 = N10567 & N1415;
  assign N10792 = N10567 & idx_w_i[8];
  assign N10793 = N10569 & N1415;
  assign N10794 = N10569 & idx_w_i[8];
  assign N10795 = N10571 & N1415;
  assign N10796 = N10571 & idx_w_i[8];
  assign N10797 = N10573 & N1415;
  assign N10798 = N10573 & idx_w_i[8];
  assign N10799 = N10575 & N1415;
  assign N10800 = N10575 & idx_w_i[8];
  assign N10801 = N10576 & N1415;
  assign N10802 = N10576 & idx_w_i[8];
  assign N10803 = N10577 & N1415;
  assign N10804 = N10577 & idx_w_i[8];
  assign N10805 = N10578 & N1415;
  assign N10806 = N10578 & idx_w_i[8];
  assign N10807 = N10579 & N1415;
  assign N10808 = N10579 & idx_w_i[8];
  assign N10809 = N10580 & N1415;
  assign N10810 = N10580 & idx_w_i[8];
  assign N10811 = N10581 & N1415;
  assign N10812 = N10581 & idx_w_i[8];
  assign N10813 = N10582 & N1415;
  assign N10814 = N10582 & idx_w_i[8];
  assign N10815 = N10583 & N1415;
  assign N10816 = N10583 & idx_w_i[8];
  assign N10817 = N10584 & N1415;
  assign N10818 = N10584 & idx_w_i[8];
  assign N10819 = N10585 & N1415;
  assign N10820 = N10585 & idx_w_i[8];
  assign N10821 = N10586 & N1415;
  assign N10822 = N10586 & idx_w_i[8];
  assign N10823 = N10587 & N1415;
  assign N10824 = N10587 & idx_w_i[8];
  assign N10825 = N10588 & N1415;
  assign N10826 = N10588 & idx_w_i[8];
  assign N10827 = N10589 & N1415;
  assign N10828 = N10589 & idx_w_i[8];
  assign N10829 = N10590 & N1415;
  assign N10830 = N10590 & idx_w_i[8];
  assign N10831 = N10591 & N1415;
  assign N10832 = N10591 & idx_w_i[8];
  assign N10833 = N10592 & N1415;
  assign N10834 = N10592 & idx_w_i[8];
  assign N10835 = N10593 & N1415;
  assign N10836 = N10593 & idx_w_i[8];
  assign N10837 = N10594 & N1415;
  assign N10838 = N10594 & idx_w_i[8];
  assign N10839 = N10595 & N1415;
  assign N10840 = N10595 & idx_w_i[8];
  assign N10841 = N10596 & N1415;
  assign N10842 = N10596 & idx_w_i[8];
  assign N10843 = N10597 & N1415;
  assign N10844 = N10597 & idx_w_i[8];
  assign N10845 = N10598 & N1415;
  assign N10846 = N10598 & idx_w_i[8];
  assign N10847 = N10599 & N1415;
  assign N10848 = N10599 & idx_w_i[8];
  assign N10849 = N10600 & N1415;
  assign N10850 = N10600 & idx_w_i[8];
  assign N10851 = N10601 & N1415;
  assign N10852 = N10601 & idx_w_i[8];
  assign N10853 = N10602 & N1415;
  assign N10854 = N10602 & idx_w_i[8];
  assign N10855 = N10603 & N1415;
  assign N10856 = N10603 & idx_w_i[8];
  assign N10857 = N10604 & N1415;
  assign N10858 = N10604 & idx_w_i[8];
  assign N10859 = N10605 & N1415;
  assign N10860 = N10605 & idx_w_i[8];
  assign N10861 = N10606 & N1415;
  assign N10862 = N10606 & idx_w_i[8];
  assign N10863 = N10384 & N1415;
  assign N10864 = N10384 & idx_w_i[8];
  assign N10865 = N10386 & N1415;
  assign N10866 = N10386 & idx_w_i[8];
  assign N10867 = N10388 & N1415;
  assign N10868 = N10388 & idx_w_i[8];
  assign N10869 = N10390 & N1415;
  assign N10870 = N10390 & idx_w_i[8];
  assign N10871 = N10392 & N1415;
  assign N10872 = N10392 & idx_w_i[8];
  assign N10873 = N10394 & N1415;
  assign N10874 = N10394 & idx_w_i[8];
  assign N10875 = N10396 & N1415;
  assign N10876 = N10396 & idx_w_i[8];
  assign N10877 = N10398 & N1415;
  assign N10878 = N10398 & idx_w_i[8];
  assign N10879 = N10400 & N1415;
  assign N10880 = N10400 & idx_w_i[8];
  assign N10881 = N10402 & N1415;
  assign N10882 = N10402 & idx_w_i[8];
  assign N10883 = N10404 & N1415;
  assign N10884 = N10404 & idx_w_i[8];
  assign N10885 = N10406 & N1415;
  assign N10886 = N10406 & idx_w_i[8];
  assign N10887 = N10408 & N1415;
  assign N10888 = N10408 & idx_w_i[8];
  assign N10889 = N10410 & N1415;
  assign N10890 = N10410 & idx_w_i[8];
  assign N10891 = N10412 & N1415;
  assign N10892 = N10412 & idx_w_i[8];
  assign N10893 = N10414 & N1415;
  assign N10894 = N10414 & idx_w_i[8];
  assign N10895 = N10416 & N1415;
  assign N10896 = N10416 & idx_w_i[8];
  assign N10897 = N10418 & N1415;
  assign N10898 = N10418 & idx_w_i[8];
  assign N10899 = N10420 & N1415;
  assign N10900 = N10420 & idx_w_i[8];
  assign N10901 = N10422 & N1415;
  assign N10902 = N10422 & idx_w_i[8];
  assign N10903 = N10424 & N1415;
  assign N10904 = N10424 & idx_w_i[8];
  assign N10905 = N10426 & N1415;
  assign N10906 = N10426 & idx_w_i[8];
  assign N10907 = N10428 & N1415;
  assign N10908 = N10428 & idx_w_i[8];
  assign N10909 = N10430 & N1415;
  assign N10910 = N10430 & idx_w_i[8];
  assign N10911 = N10432 & N1415;
  assign N10912 = N10432 & idx_w_i[8];
  assign N10913 = N10434 & N1415;
  assign N10914 = N10434 & idx_w_i[8];
  assign N10915 = N10436 & N1415;
  assign N10916 = N10436 & idx_w_i[8];
  assign N10917 = N10438 & N1415;
  assign N10918 = N10438 & idx_w_i[8];
  assign N10919 = N10440 & N1415;
  assign N10920 = N10440 & idx_w_i[8];
  assign N10921 = N10442 & N1415;
  assign N10922 = N10442 & idx_w_i[8];
  assign N10923 = N10444 & N1415;
  assign N10924 = N10444 & idx_w_i[8];
  assign N10925 = N10446 & N1415;
  assign N10926 = N10446 & idx_w_i[8];
  assign N10927 = N10448 & N1415;
  assign N10928 = N10448 & idx_w_i[8];
  assign N10929 = N10450 & N1415;
  assign N10930 = N10450 & idx_w_i[8];
  assign N10931 = N10452 & N1415;
  assign N10932 = N10452 & idx_w_i[8];
  assign N10933 = N10454 & N1415;
  assign N10934 = N10454 & idx_w_i[8];
  assign N10935 = N10456 & N1415;
  assign N10936 = N10456 & idx_w_i[8];
  assign N10937 = N10458 & N1415;
  assign N10938 = N10458 & idx_w_i[8];
  assign N10939 = N10460 & N1415;
  assign N10940 = N10460 & idx_w_i[8];
  assign N10941 = N10462 & N1415;
  assign N10942 = N10462 & idx_w_i[8];
  assign N10943 = N10464 & N1415;
  assign N10944 = N10464 & idx_w_i[8];
  assign N10945 = N10466 & N1415;
  assign N10946 = N10466 & idx_w_i[8];
  assign N10947 = N10468 & N1415;
  assign N10948 = N10468 & idx_w_i[8];
  assign N10949 = N10470 & N1415;
  assign N10950 = N10470 & idx_w_i[8];
  assign N10951 = N10472 & N1415;
  assign N10952 = N10472 & idx_w_i[8];
  assign N10953 = N10474 & N1415;
  assign N10954 = N10474 & idx_w_i[8];
  assign N10955 = N10476 & N1415;
  assign N10956 = N10476 & idx_w_i[8];
  assign N10957 = N10478 & N1415;
  assign N10958 = N10478 & idx_w_i[8];
  assign N10959 = N10480 & N1415;
  assign N10960 = N10480 & idx_w_i[8];
  assign N10961 = N10482 & N1415;
  assign N10962 = N10482 & idx_w_i[8];
  assign N10963 = N10484 & N1415;
  assign N10964 = N10484 & idx_w_i[8];
  assign N10965 = N10486 & N1415;
  assign N10966 = N10486 & idx_w_i[8];
  assign N10967 = N10488 & N1415;
  assign N10968 = N10488 & idx_w_i[8];
  assign N10969 = N10490 & N1415;
  assign N10970 = N10490 & idx_w_i[8];
  assign N10971 = N10492 & N1415;
  assign N10972 = N10492 & idx_w_i[8];
  assign N10973 = N10494 & N1415;
  assign N10974 = N10494 & idx_w_i[8];
  assign N10975 = N10496 & N1415;
  assign N10976 = N10496 & idx_w_i[8];
  assign N10977 = N10498 & N1415;
  assign N10978 = N10498 & idx_w_i[8];
  assign N10979 = N10500 & N1415;
  assign N10980 = N10500 & idx_w_i[8];
  assign N10981 = N10502 & N1415;
  assign N10982 = N10502 & idx_w_i[8];
  assign N10983 = N10504 & N1415;
  assign N10984 = N10504 & idx_w_i[8];
  assign N10985 = N10506 & N1415;
  assign N10986 = N10506 & idx_w_i[8];
  assign N10987 = N10508 & N1415;
  assign N10988 = N10508 & idx_w_i[8];
  assign N10989 = N10510 & N1415;
  assign N10990 = N10510 & idx_w_i[8];
  assign N10991 = N10512 & N1415;
  assign N10992 = N10512 & idx_w_i[8];
  assign N10993 = N10514 & N1415;
  assign N10994 = N10514 & idx_w_i[8];
  assign N10995 = N10516 & N1415;
  assign N10996 = N10516 & idx_w_i[8];
  assign N10997 = N10518 & N1415;
  assign N10998 = N10518 & idx_w_i[8];
  assign N10999 = N10520 & N1415;
  assign N11000 = N10520 & idx_w_i[8];
  assign N11001 = N10522 & N1415;
  assign N11002 = N10522 & idx_w_i[8];
  assign N11003 = N10524 & N1415;
  assign N11004 = N10524 & idx_w_i[8];
  assign N11005 = N10526 & N1415;
  assign N11006 = N10526 & idx_w_i[8];
  assign N11007 = N10528 & N1415;
  assign N11008 = N10528 & idx_w_i[8];
  assign N11009 = N10530 & N1415;
  assign N11010 = N10530 & idx_w_i[8];
  assign N11011 = N10532 & N1415;
  assign N11012 = N10532 & idx_w_i[8];
  assign N11013 = N10534 & N1415;
  assign N11014 = N10534 & idx_w_i[8];
  assign N11015 = N10536 & N1415;
  assign N11016 = N10536 & idx_w_i[8];
  assign N11017 = N10538 & N1415;
  assign N11018 = N10538 & idx_w_i[8];
  assign N11019 = N10540 & N1415;
  assign N11020 = N10540 & idx_w_i[8];
  assign N11021 = N10542 & N1415;
  assign N11022 = N10542 & idx_w_i[8];
  assign N11023 = N10544 & N1415;
  assign N11024 = N10544 & idx_w_i[8];
  assign N11025 = N10546 & N1415;
  assign N11026 = N10546 & idx_w_i[8];
  assign N11027 = N10548 & N1415;
  assign N11028 = N10548 & idx_w_i[8];
  assign N11029 = N10550 & N1415;
  assign N11030 = N10550 & idx_w_i[8];
  assign N11031 = N10552 & N1415;
  assign N11032 = N10552 & idx_w_i[8];
  assign N11033 = N10554 & N1415;
  assign N11034 = N10554 & idx_w_i[8];
  assign N11035 = N10556 & N1415;
  assign N11036 = N10556 & idx_w_i[8];
  assign N11037 = N10558 & N1415;
  assign N11038 = N10558 & idx_w_i[8];
  assign N11039 = N10560 & N1415;
  assign N11040 = N10560 & idx_w_i[8];
  assign N11041 = N10562 & N1415;
  assign N11042 = N10562 & idx_w_i[8];
  assign N11043 = N10564 & N1415;
  assign N11044 = N10564 & idx_w_i[8];
  assign N11045 = N10566 & N1415;
  assign N11046 = N10566 & idx_w_i[8];
  assign N11047 = N10568 & N1415;
  assign N11048 = N10568 & idx_w_i[8];
  assign N11049 = N10570 & N1415;
  assign N11050 = N10570 & idx_w_i[8];
  assign N11051 = N10572 & N1415;
  assign N11052 = N10572 & idx_w_i[8];
  assign N11053 = N10574 & N1415;
  assign N11054 = N10574 & idx_w_i[8];
  assign N11055 = N11537 & N1415;
  assign N11056 = N11539 & N1415;
  assign N11057 = N11541 & N1415;
  assign N11058 = N11543 & N1415;
  assign N11059 = N11545 & N1415;
  assign N11060 = N11547 & N1415;
  assign N11061 = N11549 & N1415;
  assign N11062 = N11551 & N1415;
  assign N11063 = N11553 & N1415;
  assign N11064 = N11555 & N1415;
  assign N11065 = N11557 & N1415;
  assign N11066 = N11559 & N1415;
  assign N11067 = N11561 & N1415;
  assign N11068 = N11563 & N1415;
  assign N11069 = N11565 & N1415;
  assign N11070 = N11567 & N1415;
  assign N11071 = N11569 & N1415;
  assign N11072 = N11571 & N1415;
  assign N11073 = N11573 & N1415;
  assign N11074 = N11575 & N1415;
  assign N11075 = N11577 & N1415;
  assign N11076 = N11579 & N1415;
  assign N11077 = N11581 & N1415;
  assign N11078 = N11583 & N1415;
  assign N11079 = N11585 & N1415;
  assign N11080 = N11587 & N1415;
  assign N11081 = N11589 & N1415;
  assign N11082 = N11591 & N1415;
  assign N11083 = N11593 & N1415;
  assign N11084 = N11595 & N1415;
  assign N11085 = N11597 & N1415;
  assign N11086 = N11599 & N1415;
  assign N11089 = ~idx_w_i[0];
  assign N11090 = ~idx_w_i[1];
  assign N11091 = N11089 & N11090;
  assign N11092 = N11089 & idx_w_i[1];
  assign N11093 = idx_w_i[0] & N11090;
  assign N11094 = idx_w_i[0] & idx_w_i[1];
  assign N11095 = ~idx_w_i[2];
  assign N11096 = N11091 & N11095;
  assign N11097 = N11091 & idx_w_i[2];
  assign N11098 = N11093 & N11095;
  assign N11099 = N11093 & idx_w_i[2];
  assign N11100 = N11092 & N11095;
  assign N11101 = N11092 & idx_w_i[2];
  assign N11102 = N11094 & N11095;
  assign N11103 = N11094 & idx_w_i[2];
  assign N11104 = N11096 & N2689;
  assign N11105 = N11096 & idx_w_i[3];
  assign N11106 = N11098 & N2689;
  assign N11107 = N11098 & idx_w_i[3];
  assign N11108 = N11100 & N2689;
  assign N11109 = N11100 & idx_w_i[3];
  assign N11110 = N11102 & N2689;
  assign N11111 = N11102 & idx_w_i[3];
  assign N11112 = N11097 & N2689;
  assign N11113 = N11097 & idx_w_i[3];
  assign N11114 = N11099 & N2689;
  assign N11115 = N11099 & idx_w_i[3];
  assign N11116 = N11101 & N2689;
  assign N11117 = N11101 & idx_w_i[3];
  assign N11118 = N11103 & N2689;
  assign N11119 = N11103 & idx_w_i[3];
  assign N11120 = N11104 & N2698;
  assign N11121 = N11104 & idx_w_i[4];
  assign N11122 = N11106 & N2698;
  assign N11123 = N11106 & idx_w_i[4];
  assign N11124 = N11108 & N2698;
  assign N11125 = N11108 & idx_w_i[4];
  assign N11126 = N11110 & N2698;
  assign N11127 = N11110 & idx_w_i[4];
  assign N11128 = N11112 & N2698;
  assign N11129 = N11112 & idx_w_i[4];
  assign N11130 = N11114 & N2698;
  assign N11131 = N11114 & idx_w_i[4];
  assign N11132 = N11116 & N2698;
  assign N11133 = N11116 & idx_w_i[4];
  assign N11134 = N11118 & N2698;
  assign N11135 = N11118 & idx_w_i[4];
  assign N11136 = N11105 & N2698;
  assign N11137 = N11105 & idx_w_i[4];
  assign N11138 = N11107 & N2698;
  assign N11139 = N11107 & idx_w_i[4];
  assign N11140 = N11109 & N2698;
  assign N11141 = N11109 & idx_w_i[4];
  assign N11142 = N11111 & N2698;
  assign N11143 = N11111 & idx_w_i[4];
  assign N11144 = N11113 & N2698;
  assign N11145 = N11113 & idx_w_i[4];
  assign N11146 = N11115 & N2698;
  assign N11147 = N11115 & idx_w_i[4];
  assign N11148 = N11117 & N2698;
  assign N11149 = N11117 & idx_w_i[4];
  assign N11150 = N11119 & N2698;
  assign N11151 = N11119 & idx_w_i[4];
  assign N11152 = N11120 & N1060;
  assign N11153 = N11120 & idx_w_i[5];
  assign N11154 = N11122 & N1060;
  assign N11155 = N11122 & idx_w_i[5];
  assign N11156 = N11124 & N1060;
  assign N11157 = N11124 & idx_w_i[5];
  assign N11158 = N11126 & N1060;
  assign N11159 = N11126 & idx_w_i[5];
  assign N11160 = N11128 & N1060;
  assign N11161 = N11128 & idx_w_i[5];
  assign N11162 = N11130 & N1060;
  assign N11163 = N11130 & idx_w_i[5];
  assign N11164 = N11132 & N1060;
  assign N11165 = N11132 & idx_w_i[5];
  assign N11166 = N11134 & N1060;
  assign N11167 = N11134 & idx_w_i[5];
  assign N11168 = N11136 & N1060;
  assign N11169 = N11136 & idx_w_i[5];
  assign N11170 = N11138 & N1060;
  assign N11171 = N11138 & idx_w_i[5];
  assign N11172 = N11140 & N1060;
  assign N11173 = N11140 & idx_w_i[5];
  assign N11174 = N11142 & N1060;
  assign N11175 = N11142 & idx_w_i[5];
  assign N11176 = N11144 & N1060;
  assign N11177 = N11144 & idx_w_i[5];
  assign N11178 = N11146 & N1060;
  assign N11179 = N11146 & idx_w_i[5];
  assign N11180 = N11148 & N1060;
  assign N11181 = N11148 & idx_w_i[5];
  assign N11182 = N11150 & N1060;
  assign N11183 = N11150 & idx_w_i[5];
  assign N11184 = N11121 & N1060;
  assign N11185 = N11121 & idx_w_i[5];
  assign N11186 = N11123 & N1060;
  assign N11187 = N11123 & idx_w_i[5];
  assign N11188 = N11125 & N1060;
  assign N11189 = N11125 & idx_w_i[5];
  assign N11190 = N11127 & N1060;
  assign N11191 = N11127 & idx_w_i[5];
  assign N11192 = N11129 & N1060;
  assign N11193 = N11129 & idx_w_i[5];
  assign N11194 = N11131 & N1060;
  assign N11195 = N11131 & idx_w_i[5];
  assign N11196 = N11133 & N1060;
  assign N11197 = N11133 & idx_w_i[5];
  assign N11198 = N11135 & N1060;
  assign N11199 = N11135 & idx_w_i[5];
  assign N11200 = N11137 & N1060;
  assign N11201 = N11137 & idx_w_i[5];
  assign N11202 = N11139 & N1060;
  assign N11203 = N11139 & idx_w_i[5];
  assign N11204 = N11141 & N1060;
  assign N11205 = N11141 & idx_w_i[5];
  assign N11206 = N11143 & N1060;
  assign N11207 = N11143 & idx_w_i[5];
  assign N11208 = N11145 & N1060;
  assign N11209 = N11145 & idx_w_i[5];
  assign N11210 = N11147 & N1060;
  assign N11211 = N11147 & idx_w_i[5];
  assign N11212 = N11149 & N1060;
  assign N11213 = N11149 & idx_w_i[5];
  assign N11214 = N11151 & N1060;
  assign N11215 = N11151 & idx_w_i[5];
  assign N11216 = N11152 & N1093;
  assign N11217 = N11152 & idx_w_i[6];
  assign N11218 = N11154 & N1093;
  assign N11219 = N11154 & idx_w_i[6];
  assign N11220 = N11156 & N1093;
  assign N11221 = N11156 & idx_w_i[6];
  assign N11222 = N11158 & N1093;
  assign N11223 = N11158 & idx_w_i[6];
  assign N11224 = N11160 & N1093;
  assign N11225 = N11160 & idx_w_i[6];
  assign N11226 = N11162 & N1093;
  assign N11227 = N11162 & idx_w_i[6];
  assign N11228 = N11164 & N1093;
  assign N11229 = N11164 & idx_w_i[6];
  assign N11230 = N11166 & N1093;
  assign N11231 = N11166 & idx_w_i[6];
  assign N11232 = N11168 & N1093;
  assign N11233 = N11168 & idx_w_i[6];
  assign N11234 = N11170 & N1093;
  assign N11235 = N11170 & idx_w_i[6];
  assign N11236 = N11172 & N1093;
  assign N11237 = N11172 & idx_w_i[6];
  assign N11238 = N11174 & N1093;
  assign N11239 = N11174 & idx_w_i[6];
  assign N11240 = N11176 & N1093;
  assign N11241 = N11176 & idx_w_i[6];
  assign N11242 = N11178 & N1093;
  assign N11243 = N11178 & idx_w_i[6];
  assign N11244 = N11180 & N1093;
  assign N11245 = N11180 & idx_w_i[6];
  assign N11246 = N11182 & N1093;
  assign N11247 = N11182 & idx_w_i[6];
  assign N11248 = N11184 & N1093;
  assign N11249 = N11184 & idx_w_i[6];
  assign N11250 = N11186 & N1093;
  assign N11251 = N11186 & idx_w_i[6];
  assign N11252 = N11188 & N1093;
  assign N11253 = N11188 & idx_w_i[6];
  assign N11254 = N11190 & N1093;
  assign N11255 = N11190 & idx_w_i[6];
  assign N11256 = N11192 & N1093;
  assign N11257 = N11192 & idx_w_i[6];
  assign N11258 = N11194 & N1093;
  assign N11259 = N11194 & idx_w_i[6];
  assign N11260 = N11196 & N1093;
  assign N11261 = N11196 & idx_w_i[6];
  assign N11262 = N11198 & N1093;
  assign N11263 = N11198 & idx_w_i[6];
  assign N11264 = N11200 & N1093;
  assign N11265 = N11200 & idx_w_i[6];
  assign N11266 = N11202 & N1093;
  assign N11267 = N11202 & idx_w_i[6];
  assign N11268 = N11204 & N1093;
  assign N11269 = N11204 & idx_w_i[6];
  assign N11270 = N11206 & N1093;
  assign N11271 = N11206 & idx_w_i[6];
  assign N11272 = N11208 & N1093;
  assign N11273 = N11208 & idx_w_i[6];
  assign N11274 = N11210 & N1093;
  assign N11275 = N11210 & idx_w_i[6];
  assign N11276 = N11212 & N1093;
  assign N11277 = N11212 & idx_w_i[6];
  assign N11278 = N11214 & N1093;
  assign N11279 = N11214 & idx_w_i[6];
  assign N11280 = N11153 & N1093;
  assign N11281 = N11153 & idx_w_i[6];
  assign N11282 = N11155 & N1093;
  assign N11283 = N11155 & idx_w_i[6];
  assign N11284 = N11157 & N1093;
  assign N11285 = N11157 & idx_w_i[6];
  assign N11286 = N11159 & N1093;
  assign N11287 = N11159 & idx_w_i[6];
  assign N11288 = N11161 & N1093;
  assign N11289 = N11161 & idx_w_i[6];
  assign N11290 = N11163 & N1093;
  assign N11291 = N11163 & idx_w_i[6];
  assign N11292 = N11165 & N1093;
  assign N11293 = N11165 & idx_w_i[6];
  assign N11294 = N11167 & N1093;
  assign N11295 = N11167 & idx_w_i[6];
  assign N11296 = N11169 & N1093;
  assign N11297 = N11169 & idx_w_i[6];
  assign N11298 = N11171 & N1093;
  assign N11299 = N11171 & idx_w_i[6];
  assign N11300 = N11173 & N1093;
  assign N11301 = N11173 & idx_w_i[6];
  assign N11302 = N11175 & N1093;
  assign N11303 = N11175 & idx_w_i[6];
  assign N11304 = N11177 & N1093;
  assign N11305 = N11177 & idx_w_i[6];
  assign N11306 = N11179 & N1093;
  assign N11307 = N11179 & idx_w_i[6];
  assign N11308 = N11181 & N1093;
  assign N11309 = N11181 & idx_w_i[6];
  assign N11310 = N11183 & N1093;
  assign N11311 = N11183 & idx_w_i[6];
  assign N11312 = N11185 & N1093;
  assign N11313 = N11185 & idx_w_i[6];
  assign N11314 = N11187 & N1093;
  assign N11315 = N11187 & idx_w_i[6];
  assign N11316 = N11189 & N1093;
  assign N11317 = N11189 & idx_w_i[6];
  assign N11318 = N11191 & N1093;
  assign N11319 = N11191 & idx_w_i[6];
  assign N11320 = N11193 & N1093;
  assign N11321 = N11193 & idx_w_i[6];
  assign N11322 = N11195 & N1093;
  assign N11323 = N11195 & idx_w_i[6];
  assign N11324 = N11197 & N1093;
  assign N11325 = N11197 & idx_w_i[6];
  assign N11326 = N11199 & N1093;
  assign N11327 = N11199 & idx_w_i[6];
  assign N11328 = N11201 & N1093;
  assign N11329 = N11201 & idx_w_i[6];
  assign N11330 = N11203 & N1093;
  assign N11331 = N11203 & idx_w_i[6];
  assign N11332 = N11205 & N1093;
  assign N11333 = N11205 & idx_w_i[6];
  assign N11334 = N11207 & N1093;
  assign N11335 = N11207 & idx_w_i[6];
  assign N11336 = N11209 & N1093;
  assign N11337 = N11209 & idx_w_i[6];
  assign N11338 = N11211 & N1093;
  assign N11339 = N11211 & idx_w_i[6];
  assign N11340 = N11213 & N1093;
  assign N11341 = N11213 & idx_w_i[6];
  assign N11342 = N11215 & N1093;
  assign N11343 = N11215 & idx_w_i[6];
  assign N11344 = N11216 & N1190;
  assign N11345 = N11216 & idx_w_i[7];
  assign N11346 = N11218 & N1190;
  assign N11347 = N11218 & idx_w_i[7];
  assign N11348 = N11220 & N1190;
  assign N11349 = N11220 & idx_w_i[7];
  assign N11350 = N11222 & N1190;
  assign N11351 = N11222 & idx_w_i[7];
  assign N11352 = N11224 & N1190;
  assign N11353 = N11224 & idx_w_i[7];
  assign N11354 = N11226 & N1190;
  assign N11355 = N11226 & idx_w_i[7];
  assign N11356 = N11228 & N1190;
  assign N11357 = N11228 & idx_w_i[7];
  assign N11358 = N11230 & N1190;
  assign N11359 = N11230 & idx_w_i[7];
  assign N11360 = N11232 & N1190;
  assign N11361 = N11232 & idx_w_i[7];
  assign N11362 = N11234 & N1190;
  assign N11363 = N11234 & idx_w_i[7];
  assign N11364 = N11236 & N1190;
  assign N11365 = N11236 & idx_w_i[7];
  assign N11366 = N11238 & N1190;
  assign N11367 = N11238 & idx_w_i[7];
  assign N11368 = N11240 & N1190;
  assign N11369 = N11240 & idx_w_i[7];
  assign N11370 = N11242 & N1190;
  assign N11371 = N11242 & idx_w_i[7];
  assign N11372 = N11244 & N1190;
  assign N11373 = N11244 & idx_w_i[7];
  assign N11374 = N11246 & N1190;
  assign N11375 = N11246 & idx_w_i[7];
  assign N11376 = N11248 & N1190;
  assign N11377 = N11248 & idx_w_i[7];
  assign N11378 = N11250 & N1190;
  assign N11379 = N11250 & idx_w_i[7];
  assign N11380 = N11252 & N1190;
  assign N11381 = N11252 & idx_w_i[7];
  assign N11382 = N11254 & N1190;
  assign N11383 = N11254 & idx_w_i[7];
  assign N11384 = N11256 & N1190;
  assign N11385 = N11256 & idx_w_i[7];
  assign N11386 = N11258 & N1190;
  assign N11387 = N11258 & idx_w_i[7];
  assign N11388 = N11260 & N1190;
  assign N11389 = N11260 & idx_w_i[7];
  assign N11390 = N11262 & N1190;
  assign N11391 = N11262 & idx_w_i[7];
  assign N11392 = N11264 & N1190;
  assign N11393 = N11264 & idx_w_i[7];
  assign N11394 = N11266 & N1190;
  assign N11395 = N11266 & idx_w_i[7];
  assign N11396 = N11268 & N1190;
  assign N11397 = N11268 & idx_w_i[7];
  assign N11398 = N11270 & N1190;
  assign N11399 = N11270 & idx_w_i[7];
  assign N11400 = N11272 & N1190;
  assign N11401 = N11272 & idx_w_i[7];
  assign N11402 = N11274 & N1190;
  assign N11403 = N11274 & idx_w_i[7];
  assign N11404 = N11276 & N1190;
  assign N11405 = N11276 & idx_w_i[7];
  assign N11406 = N11278 & N1190;
  assign N11407 = N11278 & idx_w_i[7];
  assign N11408 = N11280 & N1190;
  assign N11409 = N11280 & idx_w_i[7];
  assign N11410 = N11282 & N1190;
  assign N11411 = N11282 & idx_w_i[7];
  assign N11412 = N11284 & N1190;
  assign N11413 = N11284 & idx_w_i[7];
  assign N11414 = N11286 & N1190;
  assign N11415 = N11286 & idx_w_i[7];
  assign N11416 = N11288 & N1190;
  assign N11417 = N11288 & idx_w_i[7];
  assign N11418 = N11290 & N1190;
  assign N11419 = N11290 & idx_w_i[7];
  assign N11420 = N11292 & N1190;
  assign N11421 = N11292 & idx_w_i[7];
  assign N11422 = N11294 & N1190;
  assign N11423 = N11294 & idx_w_i[7];
  assign N11424 = N11296 & N1190;
  assign N11425 = N11296 & idx_w_i[7];
  assign N11426 = N11298 & N1190;
  assign N11427 = N11298 & idx_w_i[7];
  assign N11428 = N11300 & N1190;
  assign N11429 = N11300 & idx_w_i[7];
  assign N11430 = N11302 & N1190;
  assign N11431 = N11302 & idx_w_i[7];
  assign N11432 = N11304 & N1190;
  assign N11433 = N11304 & idx_w_i[7];
  assign N11434 = N11306 & N1190;
  assign N11435 = N11306 & idx_w_i[7];
  assign N11436 = N11308 & N1190;
  assign N11437 = N11308 & idx_w_i[7];
  assign N11438 = N11310 & N1190;
  assign N11439 = N11310 & idx_w_i[7];
  assign N11440 = N11312 & N1190;
  assign N11441 = N11312 & idx_w_i[7];
  assign N11442 = N11314 & N1190;
  assign N11443 = N11314 & idx_w_i[7];
  assign N11444 = N11316 & N1190;
  assign N11445 = N11316 & idx_w_i[7];
  assign N11446 = N11318 & N1190;
  assign N11447 = N11318 & idx_w_i[7];
  assign N11448 = N11320 & N1190;
  assign N11449 = N11320 & idx_w_i[7];
  assign N11450 = N11322 & N1190;
  assign N11451 = N11322 & idx_w_i[7];
  assign N11452 = N11324 & N1190;
  assign N11453 = N11324 & idx_w_i[7];
  assign N11454 = N11326 & N1190;
  assign N11455 = N11326 & idx_w_i[7];
  assign N11456 = N11328 & N1190;
  assign N11457 = N11328 & idx_w_i[7];
  assign N11458 = N11330 & N1190;
  assign N11459 = N11330 & idx_w_i[7];
  assign N11460 = N11332 & N1190;
  assign N11461 = N11332 & idx_w_i[7];
  assign N11462 = N11334 & N1190;
  assign N11463 = N11334 & idx_w_i[7];
  assign N11464 = N11336 & N1190;
  assign N11465 = N11336 & idx_w_i[7];
  assign N11466 = N11338 & N1190;
  assign N11467 = N11338 & idx_w_i[7];
  assign N11468 = N11340 & N1190;
  assign N11469 = N11340 & idx_w_i[7];
  assign N11470 = N11342 & N1190;
  assign N11471 = N11342 & idx_w_i[7];
  assign N11472 = N11217 & N1190;
  assign N11473 = N11217 & idx_w_i[7];
  assign N11474 = N11219 & N1190;
  assign N11475 = N11219 & idx_w_i[7];
  assign N11476 = N11221 & N1190;
  assign N11477 = N11221 & idx_w_i[7];
  assign N11478 = N11223 & N1190;
  assign N11479 = N11223 & idx_w_i[7];
  assign N11480 = N11225 & N1190;
  assign N11481 = N11225 & idx_w_i[7];
  assign N11482 = N11227 & N1190;
  assign N11483 = N11227 & idx_w_i[7];
  assign N11484 = N11229 & N1190;
  assign N11485 = N11229 & idx_w_i[7];
  assign N11486 = N11231 & N1190;
  assign N11487 = N11231 & idx_w_i[7];
  assign N11488 = N11233 & N1190;
  assign N11489 = N11233 & idx_w_i[7];
  assign N11490 = N11235 & N1190;
  assign N11491 = N11235 & idx_w_i[7];
  assign N11492 = N11237 & N1190;
  assign N11493 = N11237 & idx_w_i[7];
  assign N11494 = N11239 & N1190;
  assign N11495 = N11239 & idx_w_i[7];
  assign N11496 = N11241 & N1190;
  assign N11497 = N11241 & idx_w_i[7];
  assign N11498 = N11243 & N1190;
  assign N11499 = N11243 & idx_w_i[7];
  assign N11500 = N11245 & N1190;
  assign N11501 = N11245 & idx_w_i[7];
  assign N11502 = N11247 & N1190;
  assign N11503 = N11247 & idx_w_i[7];
  assign N11504 = N11249 & N1190;
  assign N11505 = N11249 & idx_w_i[7];
  assign N11506 = N11251 & N1190;
  assign N11507 = N11251 & idx_w_i[7];
  assign N11508 = N11253 & N1190;
  assign N11509 = N11253 & idx_w_i[7];
  assign N11510 = N11255 & N1190;
  assign N11511 = N11255 & idx_w_i[7];
  assign N11512 = N11257 & N1190;
  assign N11513 = N11257 & idx_w_i[7];
  assign N11514 = N11259 & N1190;
  assign N11515 = N11259 & idx_w_i[7];
  assign N11516 = N11261 & N1190;
  assign N11517 = N11261 & idx_w_i[7];
  assign N11518 = N11263 & N1190;
  assign N11519 = N11263 & idx_w_i[7];
  assign N11520 = N11265 & N1190;
  assign N11521 = N11265 & idx_w_i[7];
  assign N11522 = N11267 & N1190;
  assign N11523 = N11267 & idx_w_i[7];
  assign N11524 = N11269 & N1190;
  assign N11525 = N11269 & idx_w_i[7];
  assign N11526 = N11271 & N1190;
  assign N11527 = N11271 & idx_w_i[7];
  assign N11528 = N11273 & N1190;
  assign N11529 = N11273 & idx_w_i[7];
  assign N11530 = N11275 & N1190;
  assign N11531 = N11275 & idx_w_i[7];
  assign N11532 = N11277 & N1190;
  assign N11533 = N11277 & idx_w_i[7];
  assign N11534 = N11279 & N1190;
  assign N11535 = N11279 & idx_w_i[7];
  assign N11536 = N11281 & N1190;
  assign N11537 = N11281 & idx_w_i[7];
  assign N11538 = N11283 & N1190;
  assign N11539 = N11283 & idx_w_i[7];
  assign N11540 = N11285 & N1190;
  assign N11541 = N11285 & idx_w_i[7];
  assign N11542 = N11287 & N1190;
  assign N11543 = N11287 & idx_w_i[7];
  assign N11544 = N11289 & N1190;
  assign N11545 = N11289 & idx_w_i[7];
  assign N11546 = N11291 & N1190;
  assign N11547 = N11291 & idx_w_i[7];
  assign N11548 = N11293 & N1190;
  assign N11549 = N11293 & idx_w_i[7];
  assign N11550 = N11295 & N1190;
  assign N11551 = N11295 & idx_w_i[7];
  assign N11552 = N11297 & N1190;
  assign N11553 = N11297 & idx_w_i[7];
  assign N11554 = N11299 & N1190;
  assign N11555 = N11299 & idx_w_i[7];
  assign N11556 = N11301 & N1190;
  assign N11557 = N11301 & idx_w_i[7];
  assign N11558 = N11303 & N1190;
  assign N11559 = N11303 & idx_w_i[7];
  assign N11560 = N11305 & N1190;
  assign N11561 = N11305 & idx_w_i[7];
  assign N11562 = N11307 & N1190;
  assign N11563 = N11307 & idx_w_i[7];
  assign N11564 = N11309 & N1190;
  assign N11565 = N11309 & idx_w_i[7];
  assign N11566 = N11311 & N1190;
  assign N11567 = N11311 & idx_w_i[7];
  assign N11568 = N11313 & N1190;
  assign N11569 = N11313 & idx_w_i[7];
  assign N11570 = N11315 & N1190;
  assign N11571 = N11315 & idx_w_i[7];
  assign N11572 = N11317 & N1190;
  assign N11573 = N11317 & idx_w_i[7];
  assign N11574 = N11319 & N1190;
  assign N11575 = N11319 & idx_w_i[7];
  assign N11576 = N11321 & N1190;
  assign N11577 = N11321 & idx_w_i[7];
  assign N11578 = N11323 & N1190;
  assign N11579 = N11323 & idx_w_i[7];
  assign N11580 = N11325 & N1190;
  assign N11581 = N11325 & idx_w_i[7];
  assign N11582 = N11327 & N1190;
  assign N11583 = N11327 & idx_w_i[7];
  assign N11584 = N11329 & N1190;
  assign N11585 = N11329 & idx_w_i[7];
  assign N11586 = N11331 & N1190;
  assign N11587 = N11331 & idx_w_i[7];
  assign N11588 = N11333 & N1190;
  assign N11589 = N11333 & idx_w_i[7];
  assign N11590 = N11335 & N1190;
  assign N11591 = N11335 & idx_w_i[7];
  assign N11592 = N11337 & N1190;
  assign N11593 = N11337 & idx_w_i[7];
  assign N11594 = N11339 & N1190;
  assign N11595 = N11339 & idx_w_i[7];
  assign N11596 = N11341 & N1190;
  assign N11597 = N11341 & idx_w_i[7];
  assign N11598 = N11343 & N1190;
  assign N11599 = N11343 & idx_w_i[7];
  assign N11600 = N11344 & N1415;
  assign N11601 = N11344 & idx_w_i[8];
  assign N11602 = N11346 & N1415;
  assign N11603 = N11346 & idx_w_i[8];
  assign N11604 = N11348 & N1415;
  assign N11605 = N11348 & idx_w_i[8];
  assign N11606 = N11350 & N1415;
  assign N11607 = N11350 & idx_w_i[8];
  assign N11608 = N11352 & N1415;
  assign N11609 = N11352 & idx_w_i[8];
  assign N11610 = N11354 & N1415;
  assign N11611 = N11354 & idx_w_i[8];
  assign N11612 = N11356 & N1415;
  assign N11613 = N11356 & idx_w_i[8];
  assign N11614 = N11358 & N1415;
  assign N11615 = N11358 & idx_w_i[8];
  assign N11616 = N11360 & N1415;
  assign N11617 = N11360 & idx_w_i[8];
  assign N11618 = N11362 & N1415;
  assign N11619 = N11362 & idx_w_i[8];
  assign N11620 = N11364 & N1415;
  assign N11621 = N11364 & idx_w_i[8];
  assign N11622 = N11366 & N1415;
  assign N11623 = N11366 & idx_w_i[8];
  assign N11624 = N11368 & N1415;
  assign N11625 = N11368 & idx_w_i[8];
  assign N11626 = N11370 & N1415;
  assign N11627 = N11370 & idx_w_i[8];
  assign N11628 = N11372 & N1415;
  assign N11629 = N11372 & idx_w_i[8];
  assign N11630 = N11374 & N1415;
  assign N11631 = N11374 & idx_w_i[8];
  assign N11632 = N11376 & N1415;
  assign N11633 = N11376 & idx_w_i[8];
  assign N11634 = N11378 & N1415;
  assign N11635 = N11378 & idx_w_i[8];
  assign N11636 = N11380 & N1415;
  assign N11637 = N11380 & idx_w_i[8];
  assign N11638 = N11382 & N1415;
  assign N11639 = N11382 & idx_w_i[8];
  assign N11640 = N11384 & N1415;
  assign N11641 = N11384 & idx_w_i[8];
  assign N11642 = N11386 & N1415;
  assign N11643 = N11386 & idx_w_i[8];
  assign N11644 = N11388 & N1415;
  assign N11645 = N11388 & idx_w_i[8];
  assign N11646 = N11390 & N1415;
  assign N11647 = N11390 & idx_w_i[8];
  assign N11648 = N11392 & N1415;
  assign N11649 = N11392 & idx_w_i[8];
  assign N11650 = N11394 & N1415;
  assign N11651 = N11394 & idx_w_i[8];
  assign N11652 = N11396 & N1415;
  assign N11653 = N11396 & idx_w_i[8];
  assign N11654 = N11398 & N1415;
  assign N11655 = N11398 & idx_w_i[8];
  assign N11656 = N11400 & N1415;
  assign N11657 = N11400 & idx_w_i[8];
  assign N11658 = N11402 & N1415;
  assign N11659 = N11402 & idx_w_i[8];
  assign N11660 = N11404 & N1415;
  assign N11661 = N11404 & idx_w_i[8];
  assign N11662 = N11406 & N1415;
  assign N11663 = N11406 & idx_w_i[8];
  assign N11664 = N11408 & N1415;
  assign N11665 = N11408 & idx_w_i[8];
  assign N11666 = N11410 & N1415;
  assign N11667 = N11410 & idx_w_i[8];
  assign N11668 = N11412 & N1415;
  assign N11669 = N11412 & idx_w_i[8];
  assign N11670 = N11414 & N1415;
  assign N11671 = N11414 & idx_w_i[8];
  assign N11672 = N11416 & N1415;
  assign N11673 = N11416 & idx_w_i[8];
  assign N11674 = N11418 & N1415;
  assign N11675 = N11418 & idx_w_i[8];
  assign N11676 = N11420 & N1415;
  assign N11677 = N11420 & idx_w_i[8];
  assign N11678 = N11422 & N1415;
  assign N11679 = N11422 & idx_w_i[8];
  assign N11680 = N11424 & N1415;
  assign N11681 = N11424 & idx_w_i[8];
  assign N11682 = N11426 & N1415;
  assign N11683 = N11426 & idx_w_i[8];
  assign N11684 = N11428 & N1415;
  assign N11685 = N11428 & idx_w_i[8];
  assign N11686 = N11430 & N1415;
  assign N11687 = N11430 & idx_w_i[8];
  assign N11688 = N11432 & N1415;
  assign N11689 = N11432 & idx_w_i[8];
  assign N11690 = N11434 & N1415;
  assign N11691 = N11434 & idx_w_i[8];
  assign N11692 = N11436 & N1415;
  assign N11693 = N11436 & idx_w_i[8];
  assign N11694 = N11438 & N1415;
  assign N11695 = N11438 & idx_w_i[8];
  assign N11696 = N11440 & N1415;
  assign N11697 = N11440 & idx_w_i[8];
  assign N11698 = N11442 & N1415;
  assign N11699 = N11442 & idx_w_i[8];
  assign N11700 = N11444 & N1415;
  assign N11701 = N11444 & idx_w_i[8];
  assign N11702 = N11446 & N1415;
  assign N11703 = N11446 & idx_w_i[8];
  assign N11704 = N11448 & N1415;
  assign N11705 = N11448 & idx_w_i[8];
  assign N11706 = N11450 & N1415;
  assign N11707 = N11450 & idx_w_i[8];
  assign N11708 = N11452 & N1415;
  assign N11709 = N11452 & idx_w_i[8];
  assign N11710 = N11454 & N1415;
  assign N11711 = N11454 & idx_w_i[8];
  assign N11712 = N11456 & N1415;
  assign N11713 = N11456 & idx_w_i[8];
  assign N11714 = N11458 & N1415;
  assign N11715 = N11458 & idx_w_i[8];
  assign N11716 = N11460 & N1415;
  assign N11717 = N11460 & idx_w_i[8];
  assign N11718 = N11462 & N1415;
  assign N11719 = N11462 & idx_w_i[8];
  assign N11720 = N11464 & N1415;
  assign N11721 = N11464 & idx_w_i[8];
  assign N11722 = N11466 & N1415;
  assign N11723 = N11466 & idx_w_i[8];
  assign N11724 = N11468 & N1415;
  assign N11725 = N11468 & idx_w_i[8];
  assign N11726 = N11470 & N1415;
  assign N11727 = N11470 & idx_w_i[8];
  assign N11728 = N11472 & N1415;
  assign N11729 = N11472 & idx_w_i[8];
  assign N11730 = N11474 & N1415;
  assign N11731 = N11474 & idx_w_i[8];
  assign N11732 = N11476 & N1415;
  assign N11733 = N11476 & idx_w_i[8];
  assign N11734 = N11478 & N1415;
  assign N11735 = N11478 & idx_w_i[8];
  assign N11736 = N11480 & N1415;
  assign N11737 = N11480 & idx_w_i[8];
  assign N11738 = N11482 & N1415;
  assign N11739 = N11482 & idx_w_i[8];
  assign N11740 = N11484 & N1415;
  assign N11741 = N11484 & idx_w_i[8];
  assign N11742 = N11486 & N1415;
  assign N11743 = N11486 & idx_w_i[8];
  assign N11744 = N11488 & N1415;
  assign N11745 = N11488 & idx_w_i[8];
  assign N11746 = N11490 & N1415;
  assign N11747 = N11490 & idx_w_i[8];
  assign N11748 = N11492 & N1415;
  assign N11749 = N11492 & idx_w_i[8];
  assign N11750 = N11494 & N1415;
  assign N11751 = N11494 & idx_w_i[8];
  assign N11752 = N11496 & N1415;
  assign N11753 = N11496 & idx_w_i[8];
  assign N11754 = N11498 & N1415;
  assign N11755 = N11498 & idx_w_i[8];
  assign N11756 = N11500 & N1415;
  assign N11757 = N11500 & idx_w_i[8];
  assign N11758 = N11502 & N1415;
  assign N11759 = N11502 & idx_w_i[8];
  assign N11760 = N11504 & N1415;
  assign N11761 = N11504 & idx_w_i[8];
  assign N11762 = N11506 & N1415;
  assign N11763 = N11506 & idx_w_i[8];
  assign N11764 = N11508 & N1415;
  assign N11765 = N11508 & idx_w_i[8];
  assign N11766 = N11510 & N1415;
  assign N11767 = N11510 & idx_w_i[8];
  assign N11768 = N11512 & N1415;
  assign N11769 = N11512 & idx_w_i[8];
  assign N11770 = N11514 & N1415;
  assign N11771 = N11514 & idx_w_i[8];
  assign N11772 = N11516 & N1415;
  assign N11773 = N11516 & idx_w_i[8];
  assign N11774 = N11518 & N1415;
  assign N11775 = N11518 & idx_w_i[8];
  assign N11776 = N11520 & N1415;
  assign N11777 = N11520 & idx_w_i[8];
  assign N11778 = N11522 & N1415;
  assign N11779 = N11522 & idx_w_i[8];
  assign N11780 = N11524 & N1415;
  assign N11781 = N11524 & idx_w_i[8];
  assign N11782 = N11526 & N1415;
  assign N11783 = N11526 & idx_w_i[8];
  assign N11784 = N11528 & N1415;
  assign N11785 = N11528 & idx_w_i[8];
  assign N11786 = N11530 & N1415;
  assign N11787 = N11530 & idx_w_i[8];
  assign N11788 = N11532 & N1415;
  assign N11789 = N11532 & idx_w_i[8];
  assign N11790 = N11534 & N1415;
  assign N11791 = N11534 & idx_w_i[8];
  assign N11792 = N11536 & N1415;
  assign N11793 = N11536 & idx_w_i[8];
  assign N11794 = N11538 & N1415;
  assign N11795 = N11538 & idx_w_i[8];
  assign N11796 = N11540 & N1415;
  assign N11797 = N11540 & idx_w_i[8];
  assign N11798 = N11542 & N1415;
  assign N11799 = N11542 & idx_w_i[8];
  assign N11800 = N11544 & N1415;
  assign N11801 = N11544 & idx_w_i[8];
  assign N11802 = N11546 & N1415;
  assign N11803 = N11546 & idx_w_i[8];
  assign N11804 = N11548 & N1415;
  assign N11805 = N11548 & idx_w_i[8];
  assign N11806 = N11550 & N1415;
  assign N11807 = N11550 & idx_w_i[8];
  assign N11808 = N11552 & N1415;
  assign N11809 = N11552 & idx_w_i[8];
  assign N11810 = N11554 & N1415;
  assign N11811 = N11554 & idx_w_i[8];
  assign N11812 = N11556 & N1415;
  assign N11813 = N11556 & idx_w_i[8];
  assign N11814 = N11558 & N1415;
  assign N11815 = N11558 & idx_w_i[8];
  assign N11816 = N11560 & N1415;
  assign N11817 = N11560 & idx_w_i[8];
  assign N11818 = N11562 & N1415;
  assign N11819 = N11562 & idx_w_i[8];
  assign N11820 = N11564 & N1415;
  assign N11821 = N11564 & idx_w_i[8];
  assign N11822 = N11566 & N1415;
  assign N11823 = N11566 & idx_w_i[8];
  assign N11824 = N11568 & N1415;
  assign N11825 = N11568 & idx_w_i[8];
  assign N11826 = N11570 & N1415;
  assign N11827 = N11570 & idx_w_i[8];
  assign N11828 = N11572 & N1415;
  assign N11829 = N11572 & idx_w_i[8];
  assign N11830 = N11574 & N1415;
  assign N11831 = N11574 & idx_w_i[8];
  assign N11832 = N11576 & N1415;
  assign N11833 = N11576 & idx_w_i[8];
  assign N11834 = N11578 & N1415;
  assign N11835 = N11578 & idx_w_i[8];
  assign N11836 = N11580 & N1415;
  assign N11837 = N11580 & idx_w_i[8];
  assign N11838 = N11582 & N1415;
  assign N11839 = N11582 & idx_w_i[8];
  assign N11840 = N11584 & N1415;
  assign N11841 = N11584 & idx_w_i[8];
  assign N11842 = N11586 & N1415;
  assign N11843 = N11586 & idx_w_i[8];
  assign N11844 = N11588 & N1415;
  assign N11845 = N11588 & idx_w_i[8];
  assign N11846 = N11590 & N1415;
  assign N11847 = N11590 & idx_w_i[8];
  assign N11848 = N11592 & N1415;
  assign N11849 = N11592 & idx_w_i[8];
  assign N11850 = N11594 & N1415;
  assign N11851 = N11594 & idx_w_i[8];
  assign N11852 = N11596 & N1415;
  assign N11853 = N11596 & idx_w_i[8];
  assign N11854 = N11598 & N1415;
  assign N11855 = N11598 & idx_w_i[8];
  assign N11856 = N11345 & N1415;
  assign N11857 = N11345 & idx_w_i[8];
  assign N11858 = N11347 & N1415;
  assign N11859 = N11347 & idx_w_i[8];
  assign N11860 = N11349 & N1415;
  assign N11861 = N11349 & idx_w_i[8];
  assign N11862 = N11351 & N1415;
  assign N11863 = N11351 & idx_w_i[8];
  assign N11864 = N11353 & N1415;
  assign N11865 = N11353 & idx_w_i[8];
  assign N11866 = N11355 & N1415;
  assign N11867 = N11355 & idx_w_i[8];
  assign N11868 = N11357 & N1415;
  assign N11869 = N11357 & idx_w_i[8];
  assign N11870 = N11359 & N1415;
  assign N11871 = N11359 & idx_w_i[8];
  assign N11872 = N11361 & N1415;
  assign N11873 = N11361 & idx_w_i[8];
  assign N11874 = N11363 & N1415;
  assign N11875 = N11363 & idx_w_i[8];
  assign N11876 = N11365 & N1415;
  assign N11877 = N11365 & idx_w_i[8];
  assign N11878 = N11367 & N1415;
  assign N11879 = N11367 & idx_w_i[8];
  assign N11880 = N11369 & N1415;
  assign N11881 = N11369 & idx_w_i[8];
  assign N11882 = N11371 & N1415;
  assign N11883 = N11371 & idx_w_i[8];
  assign N11884 = N11373 & N1415;
  assign N11885 = N11373 & idx_w_i[8];
  assign N11886 = N11375 & N1415;
  assign N11887 = N11375 & idx_w_i[8];
  assign N11888 = N11377 & N1415;
  assign N11889 = N11377 & idx_w_i[8];
  assign N11890 = N11379 & N1415;
  assign N11891 = N11379 & idx_w_i[8];
  assign N11892 = N11381 & N1415;
  assign N11893 = N11381 & idx_w_i[8];
  assign N11894 = N11383 & N1415;
  assign N11895 = N11383 & idx_w_i[8];
  assign N11896 = N11385 & N1415;
  assign N11897 = N11385 & idx_w_i[8];
  assign N11898 = N11387 & N1415;
  assign N11899 = N11387 & idx_w_i[8];
  assign N11900 = N11389 & N1415;
  assign N11901 = N11389 & idx_w_i[8];
  assign N11902 = N11391 & N1415;
  assign N11903 = N11391 & idx_w_i[8];
  assign N11904 = N11393 & N1415;
  assign N11905 = N11393 & idx_w_i[8];
  assign N11906 = N11395 & N1415;
  assign N11907 = N11395 & idx_w_i[8];
  assign N11908 = N11397 & N1415;
  assign N11909 = N11397 & idx_w_i[8];
  assign N11910 = N11399 & N1415;
  assign N11911 = N11399 & idx_w_i[8];
  assign N11912 = N11401 & N1415;
  assign N11913 = N11401 & idx_w_i[8];
  assign N11914 = N11403 & N1415;
  assign N11915 = N11403 & idx_w_i[8];
  assign N11916 = N11405 & N1415;
  assign N11917 = N11405 & idx_w_i[8];
  assign N11918 = N11407 & N1415;
  assign N11919 = N11407 & idx_w_i[8];
  assign N11920 = N11409 & N1415;
  assign N11921 = N11409 & idx_w_i[8];
  assign N11922 = N11411 & N1415;
  assign N11923 = N11411 & idx_w_i[8];
  assign N11924 = N11413 & N1415;
  assign N11925 = N11413 & idx_w_i[8];
  assign N11926 = N11415 & N1415;
  assign N11927 = N11415 & idx_w_i[8];
  assign N11928 = N11417 & N1415;
  assign N11929 = N11417 & idx_w_i[8];
  assign N11930 = N11419 & N1415;
  assign N11931 = N11419 & idx_w_i[8];
  assign N11932 = N11421 & N1415;
  assign N11933 = N11421 & idx_w_i[8];
  assign N11934 = N11423 & N1415;
  assign N11935 = N11423 & idx_w_i[8];
  assign N11936 = N11425 & N1415;
  assign N11937 = N11425 & idx_w_i[8];
  assign N11938 = N11427 & N1415;
  assign N11939 = N11427 & idx_w_i[8];
  assign N11940 = N11429 & N1415;
  assign N11941 = N11429 & idx_w_i[8];
  assign N11942 = N11431 & N1415;
  assign N11943 = N11431 & idx_w_i[8];
  assign N11944 = N11433 & N1415;
  assign N11945 = N11433 & idx_w_i[8];
  assign N11946 = N11435 & N1415;
  assign N11947 = N11435 & idx_w_i[8];
  assign N11948 = N11437 & N1415;
  assign N11949 = N11437 & idx_w_i[8];
  assign N11950 = N11439 & N1415;
  assign N11951 = N11439 & idx_w_i[8];
  assign N11952 = N11441 & N1415;
  assign N11953 = N11441 & idx_w_i[8];
  assign N11954 = N11443 & N1415;
  assign N11955 = N11443 & idx_w_i[8];
  assign N11956 = N11445 & N1415;
  assign N11957 = N11445 & idx_w_i[8];
  assign N11958 = N11447 & N1415;
  assign N11959 = N11447 & idx_w_i[8];
  assign N11960 = N11449 & N1415;
  assign N11961 = N11449 & idx_w_i[8];
  assign N11962 = N11451 & N1415;
  assign N11963 = N11451 & idx_w_i[8];
  assign N11964 = N11453 & N1415;
  assign N11965 = N11453 & idx_w_i[8];
  assign N11966 = N11455 & N1415;
  assign N11967 = N11455 & idx_w_i[8];
  assign N11968 = N11457 & N1415;
  assign N11969 = N11457 & idx_w_i[8];
  assign N11970 = N11459 & N1415;
  assign N11971 = N11459 & idx_w_i[8];
  assign N11972 = N11461 & N1415;
  assign N11973 = N11461 & idx_w_i[8];
  assign N11974 = N11463 & N1415;
  assign N11975 = N11463 & idx_w_i[8];
  assign N11976 = N11465 & N1415;
  assign N11977 = N11465 & idx_w_i[8];
  assign N11978 = N11467 & N1415;
  assign N11979 = N11467 & idx_w_i[8];
  assign N11980 = N11469 & N1415;
  assign N11981 = N11469 & idx_w_i[8];
  assign N11982 = N11471 & N1415;
  assign N11983 = N11471 & idx_w_i[8];
  assign N11984 = N11473 & N1415;
  assign N11985 = N11473 & idx_w_i[8];
  assign N11986 = N11475 & N1415;
  assign N11987 = N11475 & idx_w_i[8];
  assign N11988 = N11477 & N1415;
  assign N11989 = N11477 & idx_w_i[8];
  assign N11990 = N11479 & N1415;
  assign N11991 = N11479 & idx_w_i[8];
  assign N11992 = N11481 & N1415;
  assign N11993 = N11481 & idx_w_i[8];
  assign N11994 = N11483 & N1415;
  assign N11995 = N11483 & idx_w_i[8];
  assign N11996 = N11485 & N1415;
  assign N11997 = N11485 & idx_w_i[8];
  assign N11998 = N11487 & N1415;
  assign N11999 = N11487 & idx_w_i[8];
  assign N12000 = N11489 & N1415;
  assign N12001 = N11489 & idx_w_i[8];
  assign N12002 = N11491 & N1415;
  assign N12003 = N11491 & idx_w_i[8];
  assign N12004 = N11493 & N1415;
  assign N12005 = N11493 & idx_w_i[8];
  assign N12006 = N11495 & N1415;
  assign N12007 = N11495 & idx_w_i[8];
  assign N12008 = N11497 & N1415;
  assign N12009 = N11497 & idx_w_i[8];
  assign N12010 = N11499 & N1415;
  assign N12011 = N11499 & idx_w_i[8];
  assign N12012 = N11501 & N1415;
  assign N12013 = N11501 & idx_w_i[8];
  assign N12014 = N11503 & N1415;
  assign N12015 = N11503 & idx_w_i[8];
  assign N12016 = N11505 & N1415;
  assign N12017 = N11505 & idx_w_i[8];
  assign N12018 = N11507 & N1415;
  assign N12019 = N11507 & idx_w_i[8];
  assign N12020 = N11509 & N1415;
  assign N12021 = N11509 & idx_w_i[8];
  assign N12022 = N11511 & N1415;
  assign N12023 = N11511 & idx_w_i[8];
  assign N12024 = N11513 & N1415;
  assign N12025 = N11513 & idx_w_i[8];
  assign N12026 = N11515 & N1415;
  assign N12027 = N11515 & idx_w_i[8];
  assign N12028 = N11517 & N1415;
  assign N12029 = N11517 & idx_w_i[8];
  assign N12030 = N11519 & N1415;
  assign N12031 = N11519 & idx_w_i[8];
  assign N12032 = N11521 & N1415;
  assign N12033 = N11521 & idx_w_i[8];
  assign N12034 = N11523 & N1415;
  assign N12035 = N11523 & idx_w_i[8];
  assign N12036 = N11525 & N1415;
  assign N12037 = N11525 & idx_w_i[8];
  assign N12038 = N11527 & N1415;
  assign N12039 = N11527 & idx_w_i[8];
  assign N12040 = N11529 & N1415;
  assign N12041 = N11529 & idx_w_i[8];
  assign N12042 = N11531 & N1415;
  assign N12043 = N11531 & idx_w_i[8];
  assign N12044 = N11533 & N1415;
  assign N12045 = N11533 & idx_w_i[8];
  assign N12046 = N11535 & N1415;
  assign N12047 = N11535 & idx_w_i[8];
  assign N12048 = N11537 & N1415;
  assign N12049 = N11537 & idx_w_i[8];
  assign N12050 = N11539 & N1415;
  assign N12051 = N11539 & idx_w_i[8];
  assign N12052 = N11541 & N1415;
  assign N12053 = N11541 & idx_w_i[8];
  assign N12054 = N11543 & N1415;
  assign N12055 = N11543 & idx_w_i[8];
  assign N12056 = N11545 & N1415;
  assign N12057 = N11545 & idx_w_i[8];
  assign N12058 = N11547 & N1415;
  assign N12059 = N11547 & idx_w_i[8];
  assign N12060 = N11549 & N1415;
  assign N12061 = N11549 & idx_w_i[8];
  assign N12062 = N11551 & N1415;
  assign N12063 = N11551 & idx_w_i[8];
  assign N12064 = N11553 & N1415;
  assign N12065 = N11553 & idx_w_i[8];
  assign N12066 = N11555 & N1415;
  assign N12067 = N11555 & idx_w_i[8];
  assign N12068 = N11557 & N1415;
  assign N12069 = N11557 & idx_w_i[8];
  assign N12070 = N11559 & N1415;
  assign N12071 = N11559 & idx_w_i[8];
  assign N12072 = N11561 & N1415;
  assign N12073 = N11561 & idx_w_i[8];
  assign N12074 = N11563 & N1415;
  assign N12075 = N11563 & idx_w_i[8];
  assign N12076 = N11565 & N1415;
  assign N12077 = N11565 & idx_w_i[8];
  assign N12078 = N11567 & N1415;
  assign N12079 = N11567 & idx_w_i[8];
  assign N12080 = N11569 & N1415;
  assign N12081 = N11569 & idx_w_i[8];
  assign N12082 = N11571 & N1415;
  assign N12083 = N11571 & idx_w_i[8];
  assign N12084 = N11573 & N1415;
  assign N12085 = N11573 & idx_w_i[8];
  assign N12086 = N11575 & N1415;
  assign N12087 = N11575 & idx_w_i[8];
  assign N12088 = N11577 & N1415;
  assign N12089 = N11577 & idx_w_i[8];
  assign N12090 = N11579 & N1415;
  assign N12091 = N11579 & idx_w_i[8];
  assign N12092 = N11581 & N1415;
  assign N12093 = N11581 & idx_w_i[8];
  assign N12094 = N11583 & N1415;
  assign N12095 = N11583 & idx_w_i[8];
  assign N12096 = N11585 & N1415;
  assign N12097 = N11585 & idx_w_i[8];
  assign N12098 = N11587 & N1415;
  assign N12099 = N11587 & idx_w_i[8];
  assign N12100 = N11589 & N1415;
  assign N12101 = N11589 & idx_w_i[8];
  assign N12102 = N11591 & N1415;
  assign N12103 = N11591 & idx_w_i[8];
  assign N12104 = N11593 & N1415;
  assign N12105 = N11593 & idx_w_i[8];
  assign N12106 = N11595 & N1415;
  assign N12107 = N11595 & idx_w_i[8];
  assign N12108 = N11597 & N1415;
  assign N12109 = N11597 & idx_w_i[8];
  assign N12110 = N11599 & N1415;
  assign N12111 = N11599 & idx_w_i[8];
  assign N12113 = N10255 & N1093;
  assign N12114 = N10256 & N1093;
  assign N12115 = N10257 & N1093;
  assign N12116 = N10258 & N1093;
  assign N12117 = N10259 & N1093;
  assign N12118 = N10260 & N1093;
  assign N12119 = N10261 & N1093;
  assign N12120 = N10262 & N1093;
  assign N12121 = N10263 & N1093;
  assign N12122 = N10264 & N1093;
  assign N12123 = N10265 & N1093;
  assign N12124 = N10266 & N1093;
  assign N12125 = N10267 & N1093;
  assign N12126 = N10268 & N1093;
  assign N12127 = N10269 & N1093;
  assign N12128 = N10270 & N1093;
  assign N12129 = N10271 & N1093;
  assign N12130 = N10272 & N1093;
  assign N12131 = N10273 & N1093;
  assign N12132 = N10274 & N1093;
  assign N12133 = N10275 & N1093;
  assign N12134 = N10276 & N1093;
  assign N12135 = N10277 & N1093;
  assign N12136 = N10278 & N1093;
  assign N12137 = N10279 & N1093;
  assign N12138 = N10280 & N1093;
  assign N12139 = N10281 & N1093;
  assign N12140 = N10282 & N1093;
  assign N12141 = N10283 & N1093;
  assign N12142 = N10284 & N1093;
  assign N12143 = N10285 & N1093;
  assign N12144 = N10286 & N1093;
  assign N12145 = N11153 & N1093;
  assign N12146 = N11155 & N1093;
  assign N12147 = N11157 & N1093;
  assign N12148 = N11159 & N1093;
  assign N12149 = N11161 & N1093;
  assign N12150 = N11163 & N1093;
  assign N12151 = N11165 & N1093;
  assign N12152 = N11167 & N1093;
  assign N12153 = N11169 & N1093;
  assign N12154 = N11171 & N1093;
  assign N12155 = N11173 & N1093;
  assign N12156 = N11175 & N1093;
  assign N12157 = N11177 & N1093;
  assign N12158 = N11179 & N1093;
  assign N12159 = N11181 & N1093;
  assign N12160 = N11183 & N1093;
  assign N12161 = N11185 & N1093;
  assign N12162 = N11187 & N1093;
  assign N12163 = N11189 & N1093;
  assign N12164 = N11191 & N1093;
  assign N12165 = N11193 & N1093;
  assign N12166 = N11195 & N1093;
  assign N12167 = N11197 & N1093;
  assign N12168 = N11199 & N1093;
  assign N12169 = N11201 & N1093;
  assign N12170 = N11203 & N1093;
  assign N12171 = N11205 & N1093;
  assign N12172 = N11207 & N1093;
  assign N12173 = N11209 & N1093;
  assign N12174 = N11211 & N1093;
  assign N12175 = N11213 & N1093;
  assign N12176 = N11215 & N1093;
  assign N12177 = N12113 & N1190;
  assign N12178 = N12113 & idx_w_i[7];
  assign N12179 = N12114 & N1190;
  assign N12180 = N12114 & idx_w_i[7];
  assign N12181 = N12115 & N1190;
  assign N12182 = N12115 & idx_w_i[7];
  assign N12183 = N12116 & N1190;
  assign N12184 = N12116 & idx_w_i[7];
  assign N12185 = N12117 & N1190;
  assign N12186 = N12117 & idx_w_i[7];
  assign N12187 = N12118 & N1190;
  assign N12188 = N12118 & idx_w_i[7];
  assign N12189 = N12119 & N1190;
  assign N12190 = N12119 & idx_w_i[7];
  assign N12191 = N12120 & N1190;
  assign N12192 = N12120 & idx_w_i[7];
  assign N12193 = N12121 & N1190;
  assign N12194 = N12121 & idx_w_i[7];
  assign N12195 = N12122 & N1190;
  assign N12196 = N12122 & idx_w_i[7];
  assign N12197 = N12123 & N1190;
  assign N12198 = N12123 & idx_w_i[7];
  assign N12199 = N12124 & N1190;
  assign N12200 = N12124 & idx_w_i[7];
  assign N12201 = N12125 & N1190;
  assign N12202 = N12125 & idx_w_i[7];
  assign N12203 = N12126 & N1190;
  assign N12204 = N12126 & idx_w_i[7];
  assign N12205 = N12127 & N1190;
  assign N12206 = N12127 & idx_w_i[7];
  assign N12207 = N12128 & N1190;
  assign N12208 = N12128 & idx_w_i[7];
  assign N12209 = N12129 & N1190;
  assign N12210 = N12129 & idx_w_i[7];
  assign N12211 = N12130 & N1190;
  assign N12212 = N12130 & idx_w_i[7];
  assign N12213 = N12131 & N1190;
  assign N12214 = N12131 & idx_w_i[7];
  assign N12215 = N12132 & N1190;
  assign N12216 = N12132 & idx_w_i[7];
  assign N12217 = N12133 & N1190;
  assign N12218 = N12133 & idx_w_i[7];
  assign N12219 = N12134 & N1190;
  assign N12220 = N12134 & idx_w_i[7];
  assign N12221 = N12135 & N1190;
  assign N12222 = N12135 & idx_w_i[7];
  assign N12223 = N12136 & N1190;
  assign N12224 = N12136 & idx_w_i[7];
  assign N12225 = N12137 & N1190;
  assign N12226 = N12137 & idx_w_i[7];
  assign N12227 = N12138 & N1190;
  assign N12228 = N12138 & idx_w_i[7];
  assign N12229 = N12139 & N1190;
  assign N12230 = N12139 & idx_w_i[7];
  assign N12231 = N12140 & N1190;
  assign N12232 = N12140 & idx_w_i[7];
  assign N12233 = N12141 & N1190;
  assign N12234 = N12141 & idx_w_i[7];
  assign N12235 = N12142 & N1190;
  assign N12236 = N12142 & idx_w_i[7];
  assign N12237 = N12143 & N1190;
  assign N12238 = N12143 & idx_w_i[7];
  assign N12239 = N12144 & N1190;
  assign N12240 = N12144 & idx_w_i[7];
  assign N12241 = N12145 & N1190;
  assign N12242 = N12145 & idx_w_i[7];
  assign N12243 = N12146 & N1190;
  assign N12244 = N12146 & idx_w_i[7];
  assign N12245 = N12147 & N1190;
  assign N12246 = N12147 & idx_w_i[7];
  assign N12247 = N12148 & N1190;
  assign N12248 = N12148 & idx_w_i[7];
  assign N12249 = N12149 & N1190;
  assign N12250 = N12149 & idx_w_i[7];
  assign N12251 = N12150 & N1190;
  assign N12252 = N12150 & idx_w_i[7];
  assign N12253 = N12151 & N1190;
  assign N12254 = N12151 & idx_w_i[7];
  assign N12255 = N12152 & N1190;
  assign N12256 = N12152 & idx_w_i[7];
  assign N12257 = N12153 & N1190;
  assign N12258 = N12153 & idx_w_i[7];
  assign N12259 = N12154 & N1190;
  assign N12260 = N12154 & idx_w_i[7];
  assign N12261 = N12155 & N1190;
  assign N12262 = N12155 & idx_w_i[7];
  assign N12263 = N12156 & N1190;
  assign N12264 = N12156 & idx_w_i[7];
  assign N12265 = N12157 & N1190;
  assign N12266 = N12157 & idx_w_i[7];
  assign N12267 = N12158 & N1190;
  assign N12268 = N12158 & idx_w_i[7];
  assign N12269 = N12159 & N1190;
  assign N12270 = N12159 & idx_w_i[7];
  assign N12271 = N12160 & N1190;
  assign N12272 = N12160 & idx_w_i[7];
  assign N12273 = N12161 & N1190;
  assign N12274 = N12161 & idx_w_i[7];
  assign N12275 = N12162 & N1190;
  assign N12276 = N12162 & idx_w_i[7];
  assign N12277 = N12163 & N1190;
  assign N12278 = N12163 & idx_w_i[7];
  assign N12279 = N12164 & N1190;
  assign N12280 = N12164 & idx_w_i[7];
  assign N12281 = N12165 & N1190;
  assign N12282 = N12165 & idx_w_i[7];
  assign N12283 = N12166 & N1190;
  assign N12284 = N12166 & idx_w_i[7];
  assign N12285 = N12167 & N1190;
  assign N12286 = N12167 & idx_w_i[7];
  assign N12287 = N12168 & N1190;
  assign N12288 = N12168 & idx_w_i[7];
  assign N12289 = N12169 & N1190;
  assign N12290 = N12169 & idx_w_i[7];
  assign N12291 = N12170 & N1190;
  assign N12292 = N12170 & idx_w_i[7];
  assign N12293 = N12171 & N1190;
  assign N12294 = N12171 & idx_w_i[7];
  assign N12295 = N12172 & N1190;
  assign N12296 = N12172 & idx_w_i[7];
  assign N12297 = N12173 & N1190;
  assign N12298 = N12173 & idx_w_i[7];
  assign N12299 = N12174 & N1190;
  assign N12300 = N12174 & idx_w_i[7];
  assign N12301 = N12175 & N1190;
  assign N12302 = N12175 & idx_w_i[7];
  assign N12303 = N12176 & N1190;
  assign N12304 = N12176 & idx_w_i[7];
  assign N12305 = N10288 & N1190;
  assign N12306 = N10290 & N1190;
  assign N12307 = N10292 & N1190;
  assign N12308 = N10294 & N1190;
  assign N12309 = N10296 & N1190;
  assign N12310 = N10298 & N1190;
  assign N12311 = N10300 & N1190;
  assign N12312 = N10302 & N1190;
  assign N12313 = N10304 & N1190;
  assign N12314 = N10306 & N1190;
  assign N12315 = N10308 & N1190;
  assign N12316 = N10310 & N1190;
  assign N12317 = N10312 & N1190;
  assign N12318 = N10314 & N1190;
  assign N12319 = N10316 & N1190;
  assign N12320 = N10318 & N1190;
  assign N12321 = N10320 & N1190;
  assign N12322 = N10322 & N1190;
  assign N12323 = N10324 & N1190;
  assign N12324 = N10326 & N1190;
  assign N12325 = N10328 & N1190;
  assign N12326 = N10330 & N1190;
  assign N12327 = N10332 & N1190;
  assign N12328 = N10334 & N1190;
  assign N12329 = N10336 & N1190;
  assign N12330 = N10338 & N1190;
  assign N12331 = N10340 & N1190;
  assign N12332 = N10342 & N1190;
  assign N12333 = N10344 & N1190;
  assign N12334 = N10346 & N1190;
  assign N12335 = N10348 & N1190;
  assign N12336 = N10350 & N1190;
  assign N12337 = N11281 & N1190;
  assign N12338 = N11283 & N1190;
  assign N12339 = N11285 & N1190;
  assign N12340 = N11287 & N1190;
  assign N12341 = N11289 & N1190;
  assign N12342 = N11291 & N1190;
  assign N12343 = N11293 & N1190;
  assign N12344 = N11295 & N1190;
  assign N12345 = N11297 & N1190;
  assign N12346 = N11299 & N1190;
  assign N12347 = N11301 & N1190;
  assign N12348 = N11303 & N1190;
  assign N12349 = N11305 & N1190;
  assign N12350 = N11307 & N1190;
  assign N12351 = N11309 & N1190;
  assign N12352 = N11311 & N1190;
  assign N12353 = N11313 & N1190;
  assign N12354 = N11315 & N1190;
  assign N12355 = N11317 & N1190;
  assign N12356 = N11319 & N1190;
  assign N12357 = N11321 & N1190;
  assign N12358 = N11323 & N1190;
  assign N12359 = N11325 & N1190;
  assign N12360 = N11327 & N1190;
  assign N12361 = N11329 & N1190;
  assign N12362 = N11331 & N1190;
  assign N12363 = N11333 & N1190;
  assign N12364 = N11335 & N1190;
  assign N12365 = N11337 & N1190;
  assign N12366 = N11339 & N1190;
  assign N12367 = N11341 & N1190;
  assign N12368 = N11343 & N1190;
  assign N12369 = N12177 & N1415;
  assign N12370 = N12177 & idx_w_i[8];
  assign N12371 = N12179 & N1415;
  assign N12372 = N12179 & idx_w_i[8];
  assign N12373 = N12181 & N1415;
  assign N12374 = N12181 & idx_w_i[8];
  assign N12375 = N12183 & N1415;
  assign N12376 = N12183 & idx_w_i[8];
  assign N12377 = N12185 & N1415;
  assign N12378 = N12185 & idx_w_i[8];
  assign N12379 = N12187 & N1415;
  assign N12380 = N12187 & idx_w_i[8];
  assign N12381 = N12189 & N1415;
  assign N12382 = N12189 & idx_w_i[8];
  assign N12383 = N12191 & N1415;
  assign N12384 = N12191 & idx_w_i[8];
  assign N12385 = N12193 & N1415;
  assign N12386 = N12193 & idx_w_i[8];
  assign N12387 = N12195 & N1415;
  assign N12388 = N12195 & idx_w_i[8];
  assign N12389 = N12197 & N1415;
  assign N12390 = N12197 & idx_w_i[8];
  assign N12391 = N12199 & N1415;
  assign N12392 = N12199 & idx_w_i[8];
  assign N12393 = N12201 & N1415;
  assign N12394 = N12201 & idx_w_i[8];
  assign N12395 = N12203 & N1415;
  assign N12396 = N12203 & idx_w_i[8];
  assign N12397 = N12205 & N1415;
  assign N12398 = N12205 & idx_w_i[8];
  assign N12399 = N12207 & N1415;
  assign N12400 = N12207 & idx_w_i[8];
  assign N12401 = N12209 & N1415;
  assign N12402 = N12209 & idx_w_i[8];
  assign N12403 = N12211 & N1415;
  assign N12404 = N12211 & idx_w_i[8];
  assign N12405 = N12213 & N1415;
  assign N12406 = N12213 & idx_w_i[8];
  assign N12407 = N12215 & N1415;
  assign N12408 = N12215 & idx_w_i[8];
  assign N12409 = N12217 & N1415;
  assign N12410 = N12217 & idx_w_i[8];
  assign N12411 = N12219 & N1415;
  assign N12412 = N12219 & idx_w_i[8];
  assign N12413 = N12221 & N1415;
  assign N12414 = N12221 & idx_w_i[8];
  assign N12415 = N12223 & N1415;
  assign N12416 = N12223 & idx_w_i[8];
  assign N12417 = N12225 & N1415;
  assign N12418 = N12225 & idx_w_i[8];
  assign N12419 = N12227 & N1415;
  assign N12420 = N12227 & idx_w_i[8];
  assign N12421 = N12229 & N1415;
  assign N12422 = N12229 & idx_w_i[8];
  assign N12423 = N12231 & N1415;
  assign N12424 = N12231 & idx_w_i[8];
  assign N12425 = N12233 & N1415;
  assign N12426 = N12233 & idx_w_i[8];
  assign N12427 = N12235 & N1415;
  assign N12428 = N12235 & idx_w_i[8];
  assign N12429 = N12237 & N1415;
  assign N12430 = N12237 & idx_w_i[8];
  assign N12431 = N12239 & N1415;
  assign N12432 = N12239 & idx_w_i[8];
  assign N12433 = N12241 & N1415;
  assign N12434 = N12241 & idx_w_i[8];
  assign N12435 = N12243 & N1415;
  assign N12436 = N12243 & idx_w_i[8];
  assign N12437 = N12245 & N1415;
  assign N12438 = N12245 & idx_w_i[8];
  assign N12439 = N12247 & N1415;
  assign N12440 = N12247 & idx_w_i[8];
  assign N12441 = N12249 & N1415;
  assign N12442 = N12249 & idx_w_i[8];
  assign N12443 = N12251 & N1415;
  assign N12444 = N12251 & idx_w_i[8];
  assign N12445 = N12253 & N1415;
  assign N12446 = N12253 & idx_w_i[8];
  assign N12447 = N12255 & N1415;
  assign N12448 = N12255 & idx_w_i[8];
  assign N12449 = N12257 & N1415;
  assign N12450 = N12257 & idx_w_i[8];
  assign N12451 = N12259 & N1415;
  assign N12452 = N12259 & idx_w_i[8];
  assign N12453 = N12261 & N1415;
  assign N12454 = N12261 & idx_w_i[8];
  assign N12455 = N12263 & N1415;
  assign N12456 = N12263 & idx_w_i[8];
  assign N12457 = N12265 & N1415;
  assign N12458 = N12265 & idx_w_i[8];
  assign N12459 = N12267 & N1415;
  assign N12460 = N12267 & idx_w_i[8];
  assign N12461 = N12269 & N1415;
  assign N12462 = N12269 & idx_w_i[8];
  assign N12463 = N12271 & N1415;
  assign N12464 = N12271 & idx_w_i[8];
  assign N12465 = N12273 & N1415;
  assign N12466 = N12273 & idx_w_i[8];
  assign N12467 = N12275 & N1415;
  assign N12468 = N12275 & idx_w_i[8];
  assign N12469 = N12277 & N1415;
  assign N12470 = N12277 & idx_w_i[8];
  assign N12471 = N12279 & N1415;
  assign N12472 = N12279 & idx_w_i[8];
  assign N12473 = N12281 & N1415;
  assign N12474 = N12281 & idx_w_i[8];
  assign N12475 = N12283 & N1415;
  assign N12476 = N12283 & idx_w_i[8];
  assign N12477 = N12285 & N1415;
  assign N12478 = N12285 & idx_w_i[8];
  assign N12479 = N12287 & N1415;
  assign N12480 = N12287 & idx_w_i[8];
  assign N12481 = N12289 & N1415;
  assign N12482 = N12289 & idx_w_i[8];
  assign N12483 = N12291 & N1415;
  assign N12484 = N12291 & idx_w_i[8];
  assign N12485 = N12293 & N1415;
  assign N12486 = N12293 & idx_w_i[8];
  assign N12487 = N12295 & N1415;
  assign N12488 = N12295 & idx_w_i[8];
  assign N12489 = N12297 & N1415;
  assign N12490 = N12297 & idx_w_i[8];
  assign N12491 = N12299 & N1415;
  assign N12492 = N12299 & idx_w_i[8];
  assign N12493 = N12301 & N1415;
  assign N12494 = N12301 & idx_w_i[8];
  assign N12495 = N12303 & N1415;
  assign N12496 = N12303 & idx_w_i[8];
  assign N12497 = N12305 & N1415;
  assign N12498 = N12305 & idx_w_i[8];
  assign N12499 = N12306 & N1415;
  assign N12500 = N12306 & idx_w_i[8];
  assign N12501 = N12307 & N1415;
  assign N12502 = N12307 & idx_w_i[8];
  assign N12503 = N12308 & N1415;
  assign N12504 = N12308 & idx_w_i[8];
  assign N12505 = N12309 & N1415;
  assign N12506 = N12309 & idx_w_i[8];
  assign N12507 = N12310 & N1415;
  assign N12508 = N12310 & idx_w_i[8];
  assign N12509 = N12311 & N1415;
  assign N12510 = N12311 & idx_w_i[8];
  assign N12511 = N12312 & N1415;
  assign N12512 = N12312 & idx_w_i[8];
  assign N12513 = N12313 & N1415;
  assign N12514 = N12313 & idx_w_i[8];
  assign N12515 = N12314 & N1415;
  assign N12516 = N12314 & idx_w_i[8];
  assign N12517 = N12315 & N1415;
  assign N12518 = N12315 & idx_w_i[8];
  assign N12519 = N12316 & N1415;
  assign N12520 = N12316 & idx_w_i[8];
  assign N12521 = N12317 & N1415;
  assign N12522 = N12317 & idx_w_i[8];
  assign N12523 = N12318 & N1415;
  assign N12524 = N12318 & idx_w_i[8];
  assign N12525 = N12319 & N1415;
  assign N12526 = N12319 & idx_w_i[8];
  assign N12527 = N12320 & N1415;
  assign N12528 = N12320 & idx_w_i[8];
  assign N12529 = N12321 & N1415;
  assign N12530 = N12321 & idx_w_i[8];
  assign N12531 = N12322 & N1415;
  assign N12532 = N12322 & idx_w_i[8];
  assign N12533 = N12323 & N1415;
  assign N12534 = N12323 & idx_w_i[8];
  assign N12535 = N12324 & N1415;
  assign N12536 = N12324 & idx_w_i[8];
  assign N12537 = N12325 & N1415;
  assign N12538 = N12325 & idx_w_i[8];
  assign N12539 = N12326 & N1415;
  assign N12540 = N12326 & idx_w_i[8];
  assign N12541 = N12327 & N1415;
  assign N12542 = N12327 & idx_w_i[8];
  assign N12543 = N12328 & N1415;
  assign N12544 = N12328 & idx_w_i[8];
  assign N12545 = N12329 & N1415;
  assign N12546 = N12329 & idx_w_i[8];
  assign N12547 = N12330 & N1415;
  assign N12548 = N12330 & idx_w_i[8];
  assign N12549 = N12331 & N1415;
  assign N12550 = N12331 & idx_w_i[8];
  assign N12551 = N12332 & N1415;
  assign N12552 = N12332 & idx_w_i[8];
  assign N12553 = N12333 & N1415;
  assign N12554 = N12333 & idx_w_i[8];
  assign N12555 = N12334 & N1415;
  assign N12556 = N12334 & idx_w_i[8];
  assign N12557 = N12335 & N1415;
  assign N12558 = N12335 & idx_w_i[8];
  assign N12559 = N12336 & N1415;
  assign N12560 = N12336 & idx_w_i[8];
  assign N12561 = N12337 & N1415;
  assign N12562 = N12337 & idx_w_i[8];
  assign N12563 = N12338 & N1415;
  assign N12564 = N12338 & idx_w_i[8];
  assign N12565 = N12339 & N1415;
  assign N12566 = N12339 & idx_w_i[8];
  assign N12567 = N12340 & N1415;
  assign N12568 = N12340 & idx_w_i[8];
  assign N12569 = N12341 & N1415;
  assign N12570 = N12341 & idx_w_i[8];
  assign N12571 = N12342 & N1415;
  assign N12572 = N12342 & idx_w_i[8];
  assign N12573 = N12343 & N1415;
  assign N12574 = N12343 & idx_w_i[8];
  assign N12575 = N12344 & N1415;
  assign N12576 = N12344 & idx_w_i[8];
  assign N12577 = N12345 & N1415;
  assign N12578 = N12345 & idx_w_i[8];
  assign N12579 = N12346 & N1415;
  assign N12580 = N12346 & idx_w_i[8];
  assign N12581 = N12347 & N1415;
  assign N12582 = N12347 & idx_w_i[8];
  assign N12583 = N12348 & N1415;
  assign N12584 = N12348 & idx_w_i[8];
  assign N12585 = N12349 & N1415;
  assign N12586 = N12349 & idx_w_i[8];
  assign N12587 = N12350 & N1415;
  assign N12588 = N12350 & idx_w_i[8];
  assign N12589 = N12351 & N1415;
  assign N12590 = N12351 & idx_w_i[8];
  assign N12591 = N12352 & N1415;
  assign N12592 = N12352 & idx_w_i[8];
  assign N12593 = N12353 & N1415;
  assign N12594 = N12353 & idx_w_i[8];
  assign N12595 = N12354 & N1415;
  assign N12596 = N12354 & idx_w_i[8];
  assign N12597 = N12355 & N1415;
  assign N12598 = N12355 & idx_w_i[8];
  assign N12599 = N12356 & N1415;
  assign N12600 = N12356 & idx_w_i[8];
  assign N12601 = N12357 & N1415;
  assign N12602 = N12357 & idx_w_i[8];
  assign N12603 = N12358 & N1415;
  assign N12604 = N12358 & idx_w_i[8];
  assign N12605 = N12359 & N1415;
  assign N12606 = N12359 & idx_w_i[8];
  assign N12607 = N12360 & N1415;
  assign N12608 = N12360 & idx_w_i[8];
  assign N12609 = N12361 & N1415;
  assign N12610 = N12361 & idx_w_i[8];
  assign N12611 = N12362 & N1415;
  assign N12612 = N12362 & idx_w_i[8];
  assign N12613 = N12363 & N1415;
  assign N12614 = N12363 & idx_w_i[8];
  assign N12615 = N12364 & N1415;
  assign N12616 = N12364 & idx_w_i[8];
  assign N12617 = N12365 & N1415;
  assign N12618 = N12365 & idx_w_i[8];
  assign N12619 = N12366 & N1415;
  assign N12620 = N12366 & idx_w_i[8];
  assign N12621 = N12367 & N1415;
  assign N12622 = N12367 & idx_w_i[8];
  assign N12623 = N12368 & N1415;
  assign N12624 = N12368 & idx_w_i[8];
  assign N12625 = N12178 & N1415;
  assign N12626 = N12178 & idx_w_i[8];
  assign N12627 = N12180 & N1415;
  assign N12628 = N12180 & idx_w_i[8];
  assign N12629 = N12182 & N1415;
  assign N12630 = N12182 & idx_w_i[8];
  assign N12631 = N12184 & N1415;
  assign N12632 = N12184 & idx_w_i[8];
  assign N12633 = N12186 & N1415;
  assign N12634 = N12186 & idx_w_i[8];
  assign N12635 = N12188 & N1415;
  assign N12636 = N12188 & idx_w_i[8];
  assign N12637 = N12190 & N1415;
  assign N12638 = N12190 & idx_w_i[8];
  assign N12639 = N12192 & N1415;
  assign N12640 = N12192 & idx_w_i[8];
  assign N12641 = N12194 & N1415;
  assign N12642 = N12194 & idx_w_i[8];
  assign N12643 = N12196 & N1415;
  assign N12644 = N12196 & idx_w_i[8];
  assign N12645 = N12198 & N1415;
  assign N12646 = N12198 & idx_w_i[8];
  assign N12647 = N12200 & N1415;
  assign N12648 = N12200 & idx_w_i[8];
  assign N12649 = N12202 & N1415;
  assign N12650 = N12202 & idx_w_i[8];
  assign N12651 = N12204 & N1415;
  assign N12652 = N12204 & idx_w_i[8];
  assign N12653 = N12206 & N1415;
  assign N12654 = N12206 & idx_w_i[8];
  assign N12655 = N12208 & N1415;
  assign N12656 = N12208 & idx_w_i[8];
  assign N12657 = N12210 & N1415;
  assign N12658 = N12210 & idx_w_i[8];
  assign N12659 = N12212 & N1415;
  assign N12660 = N12212 & idx_w_i[8];
  assign N12661 = N12214 & N1415;
  assign N12662 = N12214 & idx_w_i[8];
  assign N12663 = N12216 & N1415;
  assign N12664 = N12216 & idx_w_i[8];
  assign N12665 = N12218 & N1415;
  assign N12666 = N12218 & idx_w_i[8];
  assign N12667 = N12220 & N1415;
  assign N12668 = N12220 & idx_w_i[8];
  assign N12669 = N12222 & N1415;
  assign N12670 = N12222 & idx_w_i[8];
  assign N12671 = N12224 & N1415;
  assign N12672 = N12224 & idx_w_i[8];
  assign N12673 = N12226 & N1415;
  assign N12674 = N12226 & idx_w_i[8];
  assign N12675 = N12228 & N1415;
  assign N12676 = N12228 & idx_w_i[8];
  assign N12677 = N12230 & N1415;
  assign N12678 = N12230 & idx_w_i[8];
  assign N12679 = N12232 & N1415;
  assign N12680 = N12232 & idx_w_i[8];
  assign N12681 = N12234 & N1415;
  assign N12682 = N12234 & idx_w_i[8];
  assign N12683 = N12236 & N1415;
  assign N12684 = N12236 & idx_w_i[8];
  assign N12685 = N12238 & N1415;
  assign N12686 = N12238 & idx_w_i[8];
  assign N12687 = N12240 & N1415;
  assign N12688 = N12240 & idx_w_i[8];
  assign N12689 = N12242 & N1415;
  assign N12690 = N12242 & idx_w_i[8];
  assign N12691 = N12244 & N1415;
  assign N12692 = N12244 & idx_w_i[8];
  assign N12693 = N12246 & N1415;
  assign N12694 = N12246 & idx_w_i[8];
  assign N12695 = N12248 & N1415;
  assign N12696 = N12248 & idx_w_i[8];
  assign N12697 = N12250 & N1415;
  assign N12698 = N12250 & idx_w_i[8];
  assign N12699 = N12252 & N1415;
  assign N12700 = N12252 & idx_w_i[8];
  assign N12701 = N12254 & N1415;
  assign N12702 = N12254 & idx_w_i[8];
  assign N12703 = N12256 & N1415;
  assign N12704 = N12256 & idx_w_i[8];
  assign N12705 = N12258 & N1415;
  assign N12706 = N12258 & idx_w_i[8];
  assign N12707 = N12260 & N1415;
  assign N12708 = N12260 & idx_w_i[8];
  assign N12709 = N12262 & N1415;
  assign N12710 = N12262 & idx_w_i[8];
  assign N12711 = N12264 & N1415;
  assign N12712 = N12264 & idx_w_i[8];
  assign N12713 = N12266 & N1415;
  assign N12714 = N12266 & idx_w_i[8];
  assign N12715 = N12268 & N1415;
  assign N12716 = N12268 & idx_w_i[8];
  assign N12717 = N12270 & N1415;
  assign N12718 = N12270 & idx_w_i[8];
  assign N12719 = N12272 & N1415;
  assign N12720 = N12272 & idx_w_i[8];
  assign N12721 = N12274 & N1415;
  assign N12722 = N12274 & idx_w_i[8];
  assign N12723 = N12276 & N1415;
  assign N12724 = N12276 & idx_w_i[8];
  assign N12725 = N12278 & N1415;
  assign N12726 = N12278 & idx_w_i[8];
  assign N12727 = N12280 & N1415;
  assign N12728 = N12280 & idx_w_i[8];
  assign N12729 = N12282 & N1415;
  assign N12730 = N12282 & idx_w_i[8];
  assign N12731 = N12284 & N1415;
  assign N12732 = N12284 & idx_w_i[8];
  assign N12733 = N12286 & N1415;
  assign N12734 = N12286 & idx_w_i[8];
  assign N12735 = N12288 & N1415;
  assign N12736 = N12288 & idx_w_i[8];
  assign N12737 = N12290 & N1415;
  assign N12738 = N12290 & idx_w_i[8];
  assign N12739 = N12292 & N1415;
  assign N12740 = N12292 & idx_w_i[8];
  assign N12741 = N12294 & N1415;
  assign N12742 = N12294 & idx_w_i[8];
  assign N12743 = N12296 & N1415;
  assign N12744 = N12296 & idx_w_i[8];
  assign N12745 = N12298 & N1415;
  assign N12746 = N12298 & idx_w_i[8];
  assign N12747 = N12300 & N1415;
  assign N12748 = N12300 & idx_w_i[8];
  assign N12749 = N12302 & N1415;
  assign N12750 = N12302 & idx_w_i[8];
  assign N12751 = N12304 & N1415;
  assign N12752 = N12304 & idx_w_i[8];
  assign N12753 = N10512 & N1415;
  assign N12754 = N10514 & N1415;
  assign N12755 = N10516 & N1415;
  assign N12756 = N10518 & N1415;
  assign N12757 = N10520 & N1415;
  assign N12758 = N10522 & N1415;
  assign N12759 = N10524 & N1415;
  assign N12760 = N10526 & N1415;
  assign N12761 = N10528 & N1415;
  assign N12762 = N10530 & N1415;
  assign N12763 = N10532 & N1415;
  assign N12764 = N10534 & N1415;
  assign N12765 = N10536 & N1415;
  assign N12766 = N10538 & N1415;
  assign N12767 = N10540 & N1415;
  assign N12768 = N10542 & N1415;
  assign N12769 = N10544 & N1415;
  assign N12770 = N10546 & N1415;
  assign N12771 = N10548 & N1415;
  assign N12772 = N10550 & N1415;
  assign N12773 = N10552 & N1415;
  assign N12774 = N10554 & N1415;
  assign N12775 = N10556 & N1415;
  assign N12776 = N10558 & N1415;
  assign N12777 = N10560 & N1415;
  assign N12778 = N10562 & N1415;
  assign N12779 = N10564 & N1415;
  assign N12780 = N10566 & N1415;
  assign N12781 = N10568 & N1415;
  assign N12782 = N10570 & N1415;
  assign N12783 = N10572 & N1415;
  assign N12784 = N10574 & N1415;
  assign N12785 = N11537 & N1415;
  assign N12786 = N11539 & N1415;
  assign N12787 = N11541 & N1415;
  assign N12788 = N11543 & N1415;
  assign N12789 = N11545 & N1415;
  assign N12790 = N11547 & N1415;
  assign N12791 = N11549 & N1415;
  assign N12792 = N11551 & N1415;
  assign N12793 = N11553 & N1415;
  assign N12794 = N11555 & N1415;
  assign N12795 = N11557 & N1415;
  assign N12796 = N11559 & N1415;
  assign N12797 = N11561 & N1415;
  assign N12798 = N11563 & N1415;
  assign N12799 = N11565 & N1415;
  assign N12800 = N11567 & N1415;
  assign N12801 = N11569 & N1415;
  assign N12802 = N11571 & N1415;
  assign N12803 = N11573 & N1415;
  assign N12804 = N11575 & N1415;
  assign N12805 = N11577 & N1415;
  assign N12806 = N11579 & N1415;
  assign N12807 = N11581 & N1415;
  assign N12808 = N11583 & N1415;
  assign N12809 = N11585 & N1415;
  assign N12810 = N11587 & N1415;
  assign N12811 = N11589 & N1415;
  assign N12812 = N11591 & N1415;
  assign N12813 = N11593 & N1415;
  assign N12814 = N11595 & N1415;
  assign N12815 = N11597 & N1415;
  assign N12816 = N11599 & N1415;
  assign N12818 = ~N12817;
  assign N12819 = N10255 & N1093;
  assign N12820 = N10256 & N1093;
  assign N12821 = N10257 & N1093;
  assign N12822 = N10258 & N1093;
  assign N12823 = N10259 & N1093;
  assign N12824 = N10260 & N1093;
  assign N12825 = N10261 & N1093;
  assign N12826 = N10262 & N1093;
  assign N12827 = N10263 & N1093;
  assign N12828 = N10264 & N1093;
  assign N12829 = N10265 & N1093;
  assign N12830 = N10266 & N1093;
  assign N12831 = N10267 & N1093;
  assign N12832 = N10268 & N1093;
  assign N12833 = N10269 & N1093;
  assign N12834 = N10270 & N1093;
  assign N12835 = N10271 & N1093;
  assign N12836 = N10272 & N1093;
  assign N12837 = N10273 & N1093;
  assign N12838 = N10274 & N1093;
  assign N12839 = N10275 & N1093;
  assign N12840 = N10276 & N1093;
  assign N12841 = N10277 & N1093;
  assign N12842 = N10278 & N1093;
  assign N12843 = N10279 & N1093;
  assign N12844 = N10280 & N1093;
  assign N12845 = N10281 & N1093;
  assign N12846 = N10282 & N1093;
  assign N12847 = N10283 & N1093;
  assign N12848 = N10284 & N1093;
  assign N12849 = N10285 & N1093;
  assign N12850 = N10286 & N1093;
  assign N12851 = N11153 & N1093;
  assign N12852 = N11155 & N1093;
  assign N12853 = N11157 & N1093;
  assign N12854 = N11159 & N1093;
  assign N12855 = N11161 & N1093;
  assign N12856 = N11163 & N1093;
  assign N12857 = N11165 & N1093;
  assign N12858 = N11167 & N1093;
  assign N12859 = N11169 & N1093;
  assign N12860 = N11171 & N1093;
  assign N12861 = N11173 & N1093;
  assign N12862 = N11175 & N1093;
  assign N12863 = N11177 & N1093;
  assign N12864 = N11179 & N1093;
  assign N12865 = N11181 & N1093;
  assign N12866 = N11183 & N1093;
  assign N12867 = N11185 & N1093;
  assign N12868 = N11187 & N1093;
  assign N12869 = N11189 & N1093;
  assign N12870 = N11191 & N1093;
  assign N12871 = N11193 & N1093;
  assign N12872 = N11195 & N1093;
  assign N12873 = N11197 & N1093;
  assign N12874 = N11199 & N1093;
  assign N12875 = N11201 & N1093;
  assign N12876 = N11203 & N1093;
  assign N12877 = N11205 & N1093;
  assign N12878 = N11207 & N1093;
  assign N12879 = N11209 & N1093;
  assign N12880 = N11211 & N1093;
  assign N12881 = N11213 & N1093;
  assign N12882 = N11215 & N1093;
  assign N12883 = N12819 & N1190;
  assign N12884 = N12819 & idx_w_i[7];
  assign N12885 = N12820 & N1190;
  assign N12886 = N12820 & idx_w_i[7];
  assign N12887 = N12821 & N1190;
  assign N12888 = N12821 & idx_w_i[7];
  assign N12889 = N12822 & N1190;
  assign N12890 = N12822 & idx_w_i[7];
  assign N12891 = N12823 & N1190;
  assign N12892 = N12823 & idx_w_i[7];
  assign N12893 = N12824 & N1190;
  assign N12894 = N12824 & idx_w_i[7];
  assign N12895 = N12825 & N1190;
  assign N12896 = N12825 & idx_w_i[7];
  assign N12897 = N12826 & N1190;
  assign N12898 = N12826 & idx_w_i[7];
  assign N12899 = N12827 & N1190;
  assign N12900 = N12827 & idx_w_i[7];
  assign N12901 = N12828 & N1190;
  assign N12902 = N12828 & idx_w_i[7];
  assign N12903 = N12829 & N1190;
  assign N12904 = N12829 & idx_w_i[7];
  assign N12905 = N12830 & N1190;
  assign N12906 = N12830 & idx_w_i[7];
  assign N12907 = N12831 & N1190;
  assign N12908 = N12831 & idx_w_i[7];
  assign N12909 = N12832 & N1190;
  assign N12910 = N12832 & idx_w_i[7];
  assign N12911 = N12833 & N1190;
  assign N12912 = N12833 & idx_w_i[7];
  assign N12913 = N12834 & N1190;
  assign N12914 = N12834 & idx_w_i[7];
  assign N12915 = N12835 & N1190;
  assign N12916 = N12835 & idx_w_i[7];
  assign N12917 = N12836 & N1190;
  assign N12918 = N12836 & idx_w_i[7];
  assign N12919 = N12837 & N1190;
  assign N12920 = N12837 & idx_w_i[7];
  assign N12921 = N12838 & N1190;
  assign N12922 = N12838 & idx_w_i[7];
  assign N12923 = N12839 & N1190;
  assign N12924 = N12839 & idx_w_i[7];
  assign N12925 = N12840 & N1190;
  assign N12926 = N12840 & idx_w_i[7];
  assign N12927 = N12841 & N1190;
  assign N12928 = N12841 & idx_w_i[7];
  assign N12929 = N12842 & N1190;
  assign N12930 = N12842 & idx_w_i[7];
  assign N12931 = N12843 & N1190;
  assign N12932 = N12843 & idx_w_i[7];
  assign N12933 = N12844 & N1190;
  assign N12934 = N12844 & idx_w_i[7];
  assign N12935 = N12845 & N1190;
  assign N12936 = N12845 & idx_w_i[7];
  assign N12937 = N12846 & N1190;
  assign N12938 = N12846 & idx_w_i[7];
  assign N12939 = N12847 & N1190;
  assign N12940 = N12847 & idx_w_i[7];
  assign N12941 = N12848 & N1190;
  assign N12942 = N12848 & idx_w_i[7];
  assign N12943 = N12849 & N1190;
  assign N12944 = N12849 & idx_w_i[7];
  assign N12945 = N12850 & N1190;
  assign N12946 = N12850 & idx_w_i[7];
  assign N12947 = N12851 & N1190;
  assign N12948 = N12851 & idx_w_i[7];
  assign N12949 = N12852 & N1190;
  assign N12950 = N12852 & idx_w_i[7];
  assign N12951 = N12853 & N1190;
  assign N12952 = N12853 & idx_w_i[7];
  assign N12953 = N12854 & N1190;
  assign N12954 = N12854 & idx_w_i[7];
  assign N12955 = N12855 & N1190;
  assign N12956 = N12855 & idx_w_i[7];
  assign N12957 = N12856 & N1190;
  assign N12958 = N12856 & idx_w_i[7];
  assign N12959 = N12857 & N1190;
  assign N12960 = N12857 & idx_w_i[7];
  assign N12961 = N12858 & N1190;
  assign N12962 = N12858 & idx_w_i[7];
  assign N12963 = N12859 & N1190;
  assign N12964 = N12859 & idx_w_i[7];
  assign N12965 = N12860 & N1190;
  assign N12966 = N12860 & idx_w_i[7];
  assign N12967 = N12861 & N1190;
  assign N12968 = N12861 & idx_w_i[7];
  assign N12969 = N12862 & N1190;
  assign N12970 = N12862 & idx_w_i[7];
  assign N12971 = N12863 & N1190;
  assign N12972 = N12863 & idx_w_i[7];
  assign N12973 = N12864 & N1190;
  assign N12974 = N12864 & idx_w_i[7];
  assign N12975 = N12865 & N1190;
  assign N12976 = N12865 & idx_w_i[7];
  assign N12977 = N12866 & N1190;
  assign N12978 = N12866 & idx_w_i[7];
  assign N12979 = N12867 & N1190;
  assign N12980 = N12867 & idx_w_i[7];
  assign N12981 = N12868 & N1190;
  assign N12982 = N12868 & idx_w_i[7];
  assign N12983 = N12869 & N1190;
  assign N12984 = N12869 & idx_w_i[7];
  assign N12985 = N12870 & N1190;
  assign N12986 = N12870 & idx_w_i[7];
  assign N12987 = N12871 & N1190;
  assign N12988 = N12871 & idx_w_i[7];
  assign N12989 = N12872 & N1190;
  assign N12990 = N12872 & idx_w_i[7];
  assign N12991 = N12873 & N1190;
  assign N12992 = N12873 & idx_w_i[7];
  assign N12993 = N12874 & N1190;
  assign N12994 = N12874 & idx_w_i[7];
  assign N12995 = N12875 & N1190;
  assign N12996 = N12875 & idx_w_i[7];
  assign N12997 = N12876 & N1190;
  assign N12998 = N12876 & idx_w_i[7];
  assign N12999 = N12877 & N1190;
  assign N13000 = N12877 & idx_w_i[7];
  assign N13001 = N12878 & N1190;
  assign N13002 = N12878 & idx_w_i[7];
  assign N13003 = N12879 & N1190;
  assign N13004 = N12879 & idx_w_i[7];
  assign N13005 = N12880 & N1190;
  assign N13006 = N12880 & idx_w_i[7];
  assign N13007 = N12881 & N1190;
  assign N13008 = N12881 & idx_w_i[7];
  assign N13009 = N12882 & N1190;
  assign N13010 = N12882 & idx_w_i[7];
  assign N13011 = N10288 & N1190;
  assign N13012 = N10290 & N1190;
  assign N13013 = N10292 & N1190;
  assign N13014 = N10294 & N1190;
  assign N13015 = N10296 & N1190;
  assign N13016 = N10298 & N1190;
  assign N13017 = N10300 & N1190;
  assign N13018 = N10302 & N1190;
  assign N13019 = N10304 & N1190;
  assign N13020 = N10306 & N1190;
  assign N13021 = N10308 & N1190;
  assign N13022 = N10310 & N1190;
  assign N13023 = N10312 & N1190;
  assign N13024 = N10314 & N1190;
  assign N13025 = N10316 & N1190;
  assign N13026 = N10318 & N1190;
  assign N13027 = N10320 & N1190;
  assign N13028 = N10322 & N1190;
  assign N13029 = N10324 & N1190;
  assign N13030 = N10326 & N1190;
  assign N13031 = N10328 & N1190;
  assign N13032 = N10330 & N1190;
  assign N13033 = N10332 & N1190;
  assign N13034 = N10334 & N1190;
  assign N13035 = N10336 & N1190;
  assign N13036 = N10338 & N1190;
  assign N13037 = N10340 & N1190;
  assign N13038 = N10342 & N1190;
  assign N13039 = N10344 & N1190;
  assign N13040 = N10346 & N1190;
  assign N13041 = N10348 & N1190;
  assign N13042 = N10350 & N1190;
  assign N13043 = N11281 & N1190;
  assign N13044 = N11283 & N1190;
  assign N13045 = N11285 & N1190;
  assign N13046 = N11287 & N1190;
  assign N13047 = N11289 & N1190;
  assign N13048 = N11291 & N1190;
  assign N13049 = N11293 & N1190;
  assign N13050 = N11295 & N1190;
  assign N13051 = N11297 & N1190;
  assign N13052 = N11299 & N1190;
  assign N13053 = N11301 & N1190;
  assign N13054 = N11303 & N1190;
  assign N13055 = N11305 & N1190;
  assign N13056 = N11307 & N1190;
  assign N13057 = N11309 & N1190;
  assign N13058 = N11311 & N1190;
  assign N13059 = N11313 & N1190;
  assign N13060 = N11315 & N1190;
  assign N13061 = N11317 & N1190;
  assign N13062 = N11319 & N1190;
  assign N13063 = N11321 & N1190;
  assign N13064 = N11323 & N1190;
  assign N13065 = N11325 & N1190;
  assign N13066 = N11327 & N1190;
  assign N13067 = N11329 & N1190;
  assign N13068 = N11331 & N1190;
  assign N13069 = N11333 & N1190;
  assign N13070 = N11335 & N1190;
  assign N13071 = N11337 & N1190;
  assign N13072 = N11339 & N1190;
  assign N13073 = N11341 & N1190;
  assign N13074 = N11343 & N1190;
  assign N13075 = N12883 & N1415;
  assign N13076 = N12883 & idx_w_i[8];
  assign N13077 = N12885 & N1415;
  assign N13078 = N12885 & idx_w_i[8];
  assign N13079 = N12887 & N1415;
  assign N13080 = N12887 & idx_w_i[8];
  assign N13081 = N12889 & N1415;
  assign N13082 = N12889 & idx_w_i[8];
  assign N13083 = N12891 & N1415;
  assign N13084 = N12891 & idx_w_i[8];
  assign N13085 = N12893 & N1415;
  assign N13086 = N12893 & idx_w_i[8];
  assign N13087 = N12895 & N1415;
  assign N13088 = N12895 & idx_w_i[8];
  assign N13089 = N12897 & N1415;
  assign N13090 = N12897 & idx_w_i[8];
  assign N13091 = N12899 & N1415;
  assign N13092 = N12899 & idx_w_i[8];
  assign N13093 = N12901 & N1415;
  assign N13094 = N12901 & idx_w_i[8];
  assign N13095 = N12903 & N1415;
  assign N13096 = N12903 & idx_w_i[8];
  assign N13097 = N12905 & N1415;
  assign N13098 = N12905 & idx_w_i[8];
  assign N13099 = N12907 & N1415;
  assign N13100 = N12907 & idx_w_i[8];
  assign N13101 = N12909 & N1415;
  assign N13102 = N12909 & idx_w_i[8];
  assign N13103 = N12911 & N1415;
  assign N13104 = N12911 & idx_w_i[8];
  assign N13105 = N12913 & N1415;
  assign N13106 = N12913 & idx_w_i[8];
  assign N13107 = N12915 & N1415;
  assign N13108 = N12915 & idx_w_i[8];
  assign N13109 = N12917 & N1415;
  assign N13110 = N12917 & idx_w_i[8];
  assign N13111 = N12919 & N1415;
  assign N13112 = N12919 & idx_w_i[8];
  assign N13113 = N12921 & N1415;
  assign N13114 = N12921 & idx_w_i[8];
  assign N13115 = N12923 & N1415;
  assign N13116 = N12923 & idx_w_i[8];
  assign N13117 = N12925 & N1415;
  assign N13118 = N12925 & idx_w_i[8];
  assign N13119 = N12927 & N1415;
  assign N13120 = N12927 & idx_w_i[8];
  assign N13121 = N12929 & N1415;
  assign N13122 = N12929 & idx_w_i[8];
  assign N13123 = N12931 & N1415;
  assign N13124 = N12931 & idx_w_i[8];
  assign N13125 = N12933 & N1415;
  assign N13126 = N12933 & idx_w_i[8];
  assign N13127 = N12935 & N1415;
  assign N13128 = N12935 & idx_w_i[8];
  assign N13129 = N12937 & N1415;
  assign N13130 = N12937 & idx_w_i[8];
  assign N13131 = N12939 & N1415;
  assign N13132 = N12939 & idx_w_i[8];
  assign N13133 = N12941 & N1415;
  assign N13134 = N12941 & idx_w_i[8];
  assign N13135 = N12943 & N1415;
  assign N13136 = N12943 & idx_w_i[8];
  assign N13137 = N12945 & N1415;
  assign N13138 = N12945 & idx_w_i[8];
  assign N13139 = N12947 & N1415;
  assign N13140 = N12947 & idx_w_i[8];
  assign N13141 = N12949 & N1415;
  assign N13142 = N12949 & idx_w_i[8];
  assign N13143 = N12951 & N1415;
  assign N13144 = N12951 & idx_w_i[8];
  assign N13145 = N12953 & N1415;
  assign N13146 = N12953 & idx_w_i[8];
  assign N13147 = N12955 & N1415;
  assign N13148 = N12955 & idx_w_i[8];
  assign N13149 = N12957 & N1415;
  assign N13150 = N12957 & idx_w_i[8];
  assign N13151 = N12959 & N1415;
  assign N13152 = N12959 & idx_w_i[8];
  assign N13153 = N12961 & N1415;
  assign N13154 = N12961 & idx_w_i[8];
  assign N13155 = N12963 & N1415;
  assign N13156 = N12963 & idx_w_i[8];
  assign N13157 = N12965 & N1415;
  assign N13158 = N12965 & idx_w_i[8];
  assign N13159 = N12967 & N1415;
  assign N13160 = N12967 & idx_w_i[8];
  assign N13161 = N12969 & N1415;
  assign N13162 = N12969 & idx_w_i[8];
  assign N13163 = N12971 & N1415;
  assign N13164 = N12971 & idx_w_i[8];
  assign N13165 = N12973 & N1415;
  assign N13166 = N12973 & idx_w_i[8];
  assign N13167 = N12975 & N1415;
  assign N13168 = N12975 & idx_w_i[8];
  assign N13169 = N12977 & N1415;
  assign N13170 = N12977 & idx_w_i[8];
  assign N13171 = N12979 & N1415;
  assign N13172 = N12979 & idx_w_i[8];
  assign N13173 = N12981 & N1415;
  assign N13174 = N12981 & idx_w_i[8];
  assign N13175 = N12983 & N1415;
  assign N13176 = N12983 & idx_w_i[8];
  assign N13177 = N12985 & N1415;
  assign N13178 = N12985 & idx_w_i[8];
  assign N13179 = N12987 & N1415;
  assign N13180 = N12987 & idx_w_i[8];
  assign N13181 = N12989 & N1415;
  assign N13182 = N12989 & idx_w_i[8];
  assign N13183 = N12991 & N1415;
  assign N13184 = N12991 & idx_w_i[8];
  assign N13185 = N12993 & N1415;
  assign N13186 = N12993 & idx_w_i[8];
  assign N13187 = N12995 & N1415;
  assign N13188 = N12995 & idx_w_i[8];
  assign N13189 = N12997 & N1415;
  assign N13190 = N12997 & idx_w_i[8];
  assign N13191 = N12999 & N1415;
  assign N13192 = N12999 & idx_w_i[8];
  assign N13193 = N13001 & N1415;
  assign N13194 = N13001 & idx_w_i[8];
  assign N13195 = N13003 & N1415;
  assign N13196 = N13003 & idx_w_i[8];
  assign N13197 = N13005 & N1415;
  assign N13198 = N13005 & idx_w_i[8];
  assign N13199 = N13007 & N1415;
  assign N13200 = N13007 & idx_w_i[8];
  assign N13201 = N13009 & N1415;
  assign N13202 = N13009 & idx_w_i[8];
  assign N13203 = N13011 & N1415;
  assign N13204 = N13011 & idx_w_i[8];
  assign N13205 = N13012 & N1415;
  assign N13206 = N13012 & idx_w_i[8];
  assign N13207 = N13013 & N1415;
  assign N13208 = N13013 & idx_w_i[8];
  assign N13209 = N13014 & N1415;
  assign N13210 = N13014 & idx_w_i[8];
  assign N13211 = N13015 & N1415;
  assign N13212 = N13015 & idx_w_i[8];
  assign N13213 = N13016 & N1415;
  assign N13214 = N13016 & idx_w_i[8];
  assign N13215 = N13017 & N1415;
  assign N13216 = N13017 & idx_w_i[8];
  assign N13217 = N13018 & N1415;
  assign N13218 = N13018 & idx_w_i[8];
  assign N13219 = N13019 & N1415;
  assign N13220 = N13019 & idx_w_i[8];
  assign N13221 = N13020 & N1415;
  assign N13222 = N13020 & idx_w_i[8];
  assign N13223 = N13021 & N1415;
  assign N13224 = N13021 & idx_w_i[8];
  assign N13225 = N13022 & N1415;
  assign N13226 = N13022 & idx_w_i[8];
  assign N13227 = N13023 & N1415;
  assign N13228 = N13023 & idx_w_i[8];
  assign N13229 = N13024 & N1415;
  assign N13230 = N13024 & idx_w_i[8];
  assign N13231 = N13025 & N1415;
  assign N13232 = N13025 & idx_w_i[8];
  assign N13233 = N13026 & N1415;
  assign N13234 = N13026 & idx_w_i[8];
  assign N13235 = N13027 & N1415;
  assign N13236 = N13027 & idx_w_i[8];
  assign N13237 = N13028 & N1415;
  assign N13238 = N13028 & idx_w_i[8];
  assign N13239 = N13029 & N1415;
  assign N13240 = N13029 & idx_w_i[8];
  assign N13241 = N13030 & N1415;
  assign N13242 = N13030 & idx_w_i[8];
  assign N13243 = N13031 & N1415;
  assign N13244 = N13031 & idx_w_i[8];
  assign N13245 = N13032 & N1415;
  assign N13246 = N13032 & idx_w_i[8];
  assign N13247 = N13033 & N1415;
  assign N13248 = N13033 & idx_w_i[8];
  assign N13249 = N13034 & N1415;
  assign N13250 = N13034 & idx_w_i[8];
  assign N13251 = N13035 & N1415;
  assign N13252 = N13035 & idx_w_i[8];
  assign N13253 = N13036 & N1415;
  assign N13254 = N13036 & idx_w_i[8];
  assign N13255 = N13037 & N1415;
  assign N13256 = N13037 & idx_w_i[8];
  assign N13257 = N13038 & N1415;
  assign N13258 = N13038 & idx_w_i[8];
  assign N13259 = N13039 & N1415;
  assign N13260 = N13039 & idx_w_i[8];
  assign N13261 = N13040 & N1415;
  assign N13262 = N13040 & idx_w_i[8];
  assign N13263 = N13041 & N1415;
  assign N13264 = N13041 & idx_w_i[8];
  assign N13265 = N13042 & N1415;
  assign N13266 = N13042 & idx_w_i[8];
  assign N13267 = N13043 & N1415;
  assign N13268 = N13043 & idx_w_i[8];
  assign N13269 = N13044 & N1415;
  assign N13270 = N13044 & idx_w_i[8];
  assign N13271 = N13045 & N1415;
  assign N13272 = N13045 & idx_w_i[8];
  assign N13273 = N13046 & N1415;
  assign N13274 = N13046 & idx_w_i[8];
  assign N13275 = N13047 & N1415;
  assign N13276 = N13047 & idx_w_i[8];
  assign N13277 = N13048 & N1415;
  assign N13278 = N13048 & idx_w_i[8];
  assign N13279 = N13049 & N1415;
  assign N13280 = N13049 & idx_w_i[8];
  assign N13281 = N13050 & N1415;
  assign N13282 = N13050 & idx_w_i[8];
  assign N13283 = N13051 & N1415;
  assign N13284 = N13051 & idx_w_i[8];
  assign N13285 = N13052 & N1415;
  assign N13286 = N13052 & idx_w_i[8];
  assign N13287 = N13053 & N1415;
  assign N13288 = N13053 & idx_w_i[8];
  assign N13289 = N13054 & N1415;
  assign N13290 = N13054 & idx_w_i[8];
  assign N13291 = N13055 & N1415;
  assign N13292 = N13055 & idx_w_i[8];
  assign N13293 = N13056 & N1415;
  assign N13294 = N13056 & idx_w_i[8];
  assign N13295 = N13057 & N1415;
  assign N13296 = N13057 & idx_w_i[8];
  assign N13297 = N13058 & N1415;
  assign N13298 = N13058 & idx_w_i[8];
  assign N13299 = N13059 & N1415;
  assign N13300 = N13059 & idx_w_i[8];
  assign N13301 = N13060 & N1415;
  assign N13302 = N13060 & idx_w_i[8];
  assign N13303 = N13061 & N1415;
  assign N13304 = N13061 & idx_w_i[8];
  assign N13305 = N13062 & N1415;
  assign N13306 = N13062 & idx_w_i[8];
  assign N13307 = N13063 & N1415;
  assign N13308 = N13063 & idx_w_i[8];
  assign N13309 = N13064 & N1415;
  assign N13310 = N13064 & idx_w_i[8];
  assign N13311 = N13065 & N1415;
  assign N13312 = N13065 & idx_w_i[8];
  assign N13313 = N13066 & N1415;
  assign N13314 = N13066 & idx_w_i[8];
  assign N13315 = N13067 & N1415;
  assign N13316 = N13067 & idx_w_i[8];
  assign N13317 = N13068 & N1415;
  assign N13318 = N13068 & idx_w_i[8];
  assign N13319 = N13069 & N1415;
  assign N13320 = N13069 & idx_w_i[8];
  assign N13321 = N13070 & N1415;
  assign N13322 = N13070 & idx_w_i[8];
  assign N13323 = N13071 & N1415;
  assign N13324 = N13071 & idx_w_i[8];
  assign N13325 = N13072 & N1415;
  assign N13326 = N13072 & idx_w_i[8];
  assign N13327 = N13073 & N1415;
  assign N13328 = N13073 & idx_w_i[8];
  assign N13329 = N13074 & N1415;
  assign N13330 = N13074 & idx_w_i[8];
  assign N13331 = N12884 & N1415;
  assign N13332 = N12884 & idx_w_i[8];
  assign N13333 = N12886 & N1415;
  assign N13334 = N12886 & idx_w_i[8];
  assign N13335 = N12888 & N1415;
  assign N13336 = N12888 & idx_w_i[8];
  assign N13337 = N12890 & N1415;
  assign N13338 = N12890 & idx_w_i[8];
  assign N13339 = N12892 & N1415;
  assign N13340 = N12892 & idx_w_i[8];
  assign N13341 = N12894 & N1415;
  assign N13342 = N12894 & idx_w_i[8];
  assign N13343 = N12896 & N1415;
  assign N13344 = N12896 & idx_w_i[8];
  assign N13345 = N12898 & N1415;
  assign N13346 = N12898 & idx_w_i[8];
  assign N13347 = N12900 & N1415;
  assign N13348 = N12900 & idx_w_i[8];
  assign N13349 = N12902 & N1415;
  assign N13350 = N12902 & idx_w_i[8];
  assign N13351 = N12904 & N1415;
  assign N13352 = N12904 & idx_w_i[8];
  assign N13353 = N12906 & N1415;
  assign N13354 = N12906 & idx_w_i[8];
  assign N13355 = N12908 & N1415;
  assign N13356 = N12908 & idx_w_i[8];
  assign N13357 = N12910 & N1415;
  assign N13358 = N12910 & idx_w_i[8];
  assign N13359 = N12912 & N1415;
  assign N13360 = N12912 & idx_w_i[8];
  assign N13361 = N12914 & N1415;
  assign N13362 = N12914 & idx_w_i[8];
  assign N13363 = N12916 & N1415;
  assign N13364 = N12916 & idx_w_i[8];
  assign N13365 = N12918 & N1415;
  assign N13366 = N12918 & idx_w_i[8];
  assign N13367 = N12920 & N1415;
  assign N13368 = N12920 & idx_w_i[8];
  assign N13369 = N12922 & N1415;
  assign N13370 = N12922 & idx_w_i[8];
  assign N13371 = N12924 & N1415;
  assign N13372 = N12924 & idx_w_i[8];
  assign N13373 = N12926 & N1415;
  assign N13374 = N12926 & idx_w_i[8];
  assign N13375 = N12928 & N1415;
  assign N13376 = N12928 & idx_w_i[8];
  assign N13377 = N12930 & N1415;
  assign N13378 = N12930 & idx_w_i[8];
  assign N13379 = N12932 & N1415;
  assign N13380 = N12932 & idx_w_i[8];
  assign N13381 = N12934 & N1415;
  assign N13382 = N12934 & idx_w_i[8];
  assign N13383 = N12936 & N1415;
  assign N13384 = N12936 & idx_w_i[8];
  assign N13385 = N12938 & N1415;
  assign N13386 = N12938 & idx_w_i[8];
  assign N13387 = N12940 & N1415;
  assign N13388 = N12940 & idx_w_i[8];
  assign N13389 = N12942 & N1415;
  assign N13390 = N12942 & idx_w_i[8];
  assign N13391 = N12944 & N1415;
  assign N13392 = N12944 & idx_w_i[8];
  assign N13393 = N12946 & N1415;
  assign N13394 = N12946 & idx_w_i[8];
  assign N13395 = N12948 & N1415;
  assign N13396 = N12948 & idx_w_i[8];
  assign N13397 = N12950 & N1415;
  assign N13398 = N12950 & idx_w_i[8];
  assign N13399 = N12952 & N1415;
  assign N13400 = N12952 & idx_w_i[8];
  assign N13401 = N12954 & N1415;
  assign N13402 = N12954 & idx_w_i[8];
  assign N13403 = N12956 & N1415;
  assign N13404 = N12956 & idx_w_i[8];
  assign N13405 = N12958 & N1415;
  assign N13406 = N12958 & idx_w_i[8];
  assign N13407 = N12960 & N1415;
  assign N13408 = N12960 & idx_w_i[8];
  assign N13409 = N12962 & N1415;
  assign N13410 = N12962 & idx_w_i[8];
  assign N13411 = N12964 & N1415;
  assign N13412 = N12964 & idx_w_i[8];
  assign N13413 = N12966 & N1415;
  assign N13414 = N12966 & idx_w_i[8];
  assign N13415 = N12968 & N1415;
  assign N13416 = N12968 & idx_w_i[8];
  assign N13417 = N12970 & N1415;
  assign N13418 = N12970 & idx_w_i[8];
  assign N13419 = N12972 & N1415;
  assign N13420 = N12972 & idx_w_i[8];
  assign N13421 = N12974 & N1415;
  assign N13422 = N12974 & idx_w_i[8];
  assign N13423 = N12976 & N1415;
  assign N13424 = N12976 & idx_w_i[8];
  assign N13425 = N12978 & N1415;
  assign N13426 = N12978 & idx_w_i[8];
  assign N13427 = N12980 & N1415;
  assign N13428 = N12980 & idx_w_i[8];
  assign N13429 = N12982 & N1415;
  assign N13430 = N12982 & idx_w_i[8];
  assign N13431 = N12984 & N1415;
  assign N13432 = N12984 & idx_w_i[8];
  assign N13433 = N12986 & N1415;
  assign N13434 = N12986 & idx_w_i[8];
  assign N13435 = N12988 & N1415;
  assign N13436 = N12988 & idx_w_i[8];
  assign N13437 = N12990 & N1415;
  assign N13438 = N12990 & idx_w_i[8];
  assign N13439 = N12992 & N1415;
  assign N13440 = N12992 & idx_w_i[8];
  assign N13441 = N12994 & N1415;
  assign N13442 = N12994 & idx_w_i[8];
  assign N13443 = N12996 & N1415;
  assign N13444 = N12996 & idx_w_i[8];
  assign N13445 = N12998 & N1415;
  assign N13446 = N12998 & idx_w_i[8];
  assign N13447 = N13000 & N1415;
  assign N13448 = N13000 & idx_w_i[8];
  assign N13449 = N13002 & N1415;
  assign N13450 = N13002 & idx_w_i[8];
  assign N13451 = N13004 & N1415;
  assign N13452 = N13004 & idx_w_i[8];
  assign N13453 = N13006 & N1415;
  assign N13454 = N13006 & idx_w_i[8];
  assign N13455 = N13008 & N1415;
  assign N13456 = N13008 & idx_w_i[8];
  assign N13457 = N13010 & N1415;
  assign N13458 = N13010 & idx_w_i[8];
  assign N13459 = N10512 & N1415;
  assign N13460 = N10514 & N1415;
  assign N13461 = N10516 & N1415;
  assign N13462 = N10518 & N1415;
  assign N13463 = N10520 & N1415;
  assign N13464 = N10522 & N1415;
  assign N13465 = N10524 & N1415;
  assign N13466 = N10526 & N1415;
  assign N13467 = N10528 & N1415;
  assign N13468 = N10530 & N1415;
  assign N13469 = N10532 & N1415;
  assign N13470 = N10534 & N1415;
  assign N13471 = N10536 & N1415;
  assign N13472 = N10538 & N1415;
  assign N13473 = N10540 & N1415;
  assign N13474 = N10542 & N1415;
  assign N13475 = N10544 & N1415;
  assign N13476 = N10546 & N1415;
  assign N13477 = N10548 & N1415;
  assign N13478 = N10550 & N1415;
  assign N13479 = N10552 & N1415;
  assign N13480 = N10554 & N1415;
  assign N13481 = N10556 & N1415;
  assign N13482 = N10558 & N1415;
  assign N13483 = N10560 & N1415;
  assign N13484 = N10562 & N1415;
  assign N13485 = N10564 & N1415;
  assign N13486 = N10566 & N1415;
  assign N13487 = N10568 & N1415;
  assign N13488 = N10570 & N1415;
  assign N13489 = N10572 & N1415;
  assign N13490 = N10574 & N1415;
  assign N13491 = N11537 & N1415;
  assign N13492 = N11539 & N1415;
  assign N13493 = N11541 & N1415;
  assign N13494 = N11543 & N1415;
  assign N13495 = N11545 & N1415;
  assign N13496 = N11547 & N1415;
  assign N13497 = N11549 & N1415;
  assign N13498 = N11551 & N1415;
  assign N13499 = N11553 & N1415;
  assign N13500 = N11555 & N1415;
  assign N13501 = N11557 & N1415;
  assign N13502 = N11559 & N1415;
  assign N13503 = N11561 & N1415;
  assign N13504 = N11563 & N1415;
  assign N13505 = N11565 & N1415;
  assign N13506 = N11567 & N1415;
  assign N13507 = N11569 & N1415;
  assign N13508 = N11571 & N1415;
  assign N13509 = N11573 & N1415;
  assign N13510 = N11575 & N1415;
  assign N13511 = N11577 & N1415;
  assign N13512 = N11579 & N1415;
  assign N13513 = N11581 & N1415;
  assign N13514 = N11583 & N1415;
  assign N13515 = N11585 & N1415;
  assign N13516 = N11587 & N1415;
  assign N13517 = N11589 & N1415;
  assign N13518 = N11591 & N1415;
  assign N13519 = N11593 & N1415;
  assign N13520 = N11595 & N1415;
  assign N13521 = N11597 & N1415;
  assign N13522 = N11599 & N1415;
  assign N14037 = N11152 & N1093;
  assign N14038 = N11154 & N1093;
  assign N14039 = N11156 & N1093;
  assign N14040 = N11158 & N1093;
  assign N14041 = N11160 & N1093;
  assign N14042 = N11162 & N1093;
  assign N14043 = N11164 & N1093;
  assign N14044 = N11166 & N1093;
  assign N14045 = N11168 & N1093;
  assign N14046 = N11170 & N1093;
  assign N14047 = N11172 & N1093;
  assign N14048 = N11174 & N1093;
  assign N14049 = N11176 & N1093;
  assign N14050 = N11178 & N1093;
  assign N14051 = N11180 & N1093;
  assign N14052 = N11182 & N1093;
  assign N14053 = N11184 & N1093;
  assign N14054 = N11186 & N1093;
  assign N14055 = N11188 & N1093;
  assign N14056 = N11190 & N1093;
  assign N14057 = N11192 & N1093;
  assign N14058 = N11194 & N1093;
  assign N14059 = N11196 & N1093;
  assign N14060 = N11198 & N1093;
  assign N14061 = N11200 & N1093;
  assign N14062 = N11202 & N1093;
  assign N14063 = N11204 & N1093;
  assign N14064 = N11206 & N1093;
  assign N14065 = N11208 & N1093;
  assign N14066 = N11210 & N1093;
  assign N14067 = N11212 & N1093;
  assign N14068 = N11214 & N1093;
  assign N14069 = N11153 & N1093;
  assign N14070 = N11155 & N1093;
  assign N14071 = N11157 & N1093;
  assign N14072 = N11159 & N1093;
  assign N14073 = N11161 & N1093;
  assign N14074 = N11163 & N1093;
  assign N14075 = N11165 & N1093;
  assign N14076 = N11167 & N1093;
  assign N14077 = N11169 & N1093;
  assign N14078 = N11171 & N1093;
  assign N14079 = N11173 & N1093;
  assign N14080 = N11175 & N1093;
  assign N14081 = N11177 & N1093;
  assign N14082 = N11179 & N1093;
  assign N14083 = N11181 & N1093;
  assign N14084 = N11183 & N1093;
  assign N14085 = N11185 & N1093;
  assign N14086 = N11187 & N1093;
  assign N14087 = N11189 & N1093;
  assign N14088 = N11191 & N1093;
  assign N14089 = N11193 & N1093;
  assign N14090 = N11195 & N1093;
  assign N14091 = N11197 & N1093;
  assign N14092 = N11199 & N1093;
  assign N14093 = N11201 & N1093;
  assign N14094 = N11203 & N1093;
  assign N14095 = N11205 & N1093;
  assign N14096 = N11207 & N1093;
  assign N14097 = N11209 & N1093;
  assign N14098 = N11211 & N1093;
  assign N14099 = N11213 & N1093;
  assign N14100 = N11215 & N1093;
  assign N14101 = N14037 & N1190;
  assign N14102 = N14037 & idx_w_i[7];
  assign N14103 = N14038 & N1190;
  assign N14104 = N14038 & idx_w_i[7];
  assign N14105 = N14039 & N1190;
  assign N14106 = N14039 & idx_w_i[7];
  assign N14107 = N14040 & N1190;
  assign N14108 = N14040 & idx_w_i[7];
  assign N14109 = N14041 & N1190;
  assign N14110 = N14041 & idx_w_i[7];
  assign N14111 = N14042 & N1190;
  assign N14112 = N14042 & idx_w_i[7];
  assign N14113 = N14043 & N1190;
  assign N14114 = N14043 & idx_w_i[7];
  assign N14115 = N14044 & N1190;
  assign N14116 = N14044 & idx_w_i[7];
  assign N14117 = N14045 & N1190;
  assign N14118 = N14045 & idx_w_i[7];
  assign N14119 = N14046 & N1190;
  assign N14120 = N14046 & idx_w_i[7];
  assign N14121 = N14047 & N1190;
  assign N14122 = N14047 & idx_w_i[7];
  assign N14123 = N14048 & N1190;
  assign N14124 = N14048 & idx_w_i[7];
  assign N14125 = N14049 & N1190;
  assign N14126 = N14049 & idx_w_i[7];
  assign N14127 = N14050 & N1190;
  assign N14128 = N14050 & idx_w_i[7];
  assign N14129 = N14051 & N1190;
  assign N14130 = N14051 & idx_w_i[7];
  assign N14131 = N14052 & N1190;
  assign N14132 = N14052 & idx_w_i[7];
  assign N14133 = N14053 & N1190;
  assign N14134 = N14053 & idx_w_i[7];
  assign N14135 = N14054 & N1190;
  assign N14136 = N14054 & idx_w_i[7];
  assign N14137 = N14055 & N1190;
  assign N14138 = N14055 & idx_w_i[7];
  assign N14139 = N14056 & N1190;
  assign N14140 = N14056 & idx_w_i[7];
  assign N14141 = N14057 & N1190;
  assign N14142 = N14057 & idx_w_i[7];
  assign N14143 = N14058 & N1190;
  assign N14144 = N14058 & idx_w_i[7];
  assign N14145 = N14059 & N1190;
  assign N14146 = N14059 & idx_w_i[7];
  assign N14147 = N14060 & N1190;
  assign N14148 = N14060 & idx_w_i[7];
  assign N14149 = N14061 & N1190;
  assign N14150 = N14061 & idx_w_i[7];
  assign N14151 = N14062 & N1190;
  assign N14152 = N14062 & idx_w_i[7];
  assign N14153 = N14063 & N1190;
  assign N14154 = N14063 & idx_w_i[7];
  assign N14155 = N14064 & N1190;
  assign N14156 = N14064 & idx_w_i[7];
  assign N14157 = N14065 & N1190;
  assign N14158 = N14065 & idx_w_i[7];
  assign N14159 = N14066 & N1190;
  assign N14160 = N14066 & idx_w_i[7];
  assign N14161 = N14067 & N1190;
  assign N14162 = N14067 & idx_w_i[7];
  assign N14163 = N14068 & N1190;
  assign N14164 = N14068 & idx_w_i[7];
  assign N14165 = N14069 & N1190;
  assign N14166 = N14069 & idx_w_i[7];
  assign N14167 = N14070 & N1190;
  assign N14168 = N14070 & idx_w_i[7];
  assign N14169 = N14071 & N1190;
  assign N14170 = N14071 & idx_w_i[7];
  assign N14171 = N14072 & N1190;
  assign N14172 = N14072 & idx_w_i[7];
  assign N14173 = N14073 & N1190;
  assign N14174 = N14073 & idx_w_i[7];
  assign N14175 = N14074 & N1190;
  assign N14176 = N14074 & idx_w_i[7];
  assign N14177 = N14075 & N1190;
  assign N14178 = N14075 & idx_w_i[7];
  assign N14179 = N14076 & N1190;
  assign N14180 = N14076 & idx_w_i[7];
  assign N14181 = N14077 & N1190;
  assign N14182 = N14077 & idx_w_i[7];
  assign N14183 = N14078 & N1190;
  assign N14184 = N14078 & idx_w_i[7];
  assign N14185 = N14079 & N1190;
  assign N14186 = N14079 & idx_w_i[7];
  assign N14187 = N14080 & N1190;
  assign N14188 = N14080 & idx_w_i[7];
  assign N14189 = N14081 & N1190;
  assign N14190 = N14081 & idx_w_i[7];
  assign N14191 = N14082 & N1190;
  assign N14192 = N14082 & idx_w_i[7];
  assign N14193 = N14083 & N1190;
  assign N14194 = N14083 & idx_w_i[7];
  assign N14195 = N14084 & N1190;
  assign N14196 = N14084 & idx_w_i[7];
  assign N14197 = N14085 & N1190;
  assign N14198 = N14085 & idx_w_i[7];
  assign N14199 = N14086 & N1190;
  assign N14200 = N14086 & idx_w_i[7];
  assign N14201 = N14087 & N1190;
  assign N14202 = N14087 & idx_w_i[7];
  assign N14203 = N14088 & N1190;
  assign N14204 = N14088 & idx_w_i[7];
  assign N14205 = N14089 & N1190;
  assign N14206 = N14089 & idx_w_i[7];
  assign N14207 = N14090 & N1190;
  assign N14208 = N14090 & idx_w_i[7];
  assign N14209 = N14091 & N1190;
  assign N14210 = N14091 & idx_w_i[7];
  assign N14211 = N14092 & N1190;
  assign N14212 = N14092 & idx_w_i[7];
  assign N14213 = N14093 & N1190;
  assign N14214 = N14093 & idx_w_i[7];
  assign N14215 = N14094 & N1190;
  assign N14216 = N14094 & idx_w_i[7];
  assign N14217 = N14095 & N1190;
  assign N14218 = N14095 & idx_w_i[7];
  assign N14219 = N14096 & N1190;
  assign N14220 = N14096 & idx_w_i[7];
  assign N14221 = N14097 & N1190;
  assign N14222 = N14097 & idx_w_i[7];
  assign N14223 = N14098 & N1190;
  assign N14224 = N14098 & idx_w_i[7];
  assign N14225 = N14099 & N1190;
  assign N14226 = N14099 & idx_w_i[7];
  assign N14227 = N14100 & N1190;
  assign N14228 = N14100 & idx_w_i[7];
  assign N14229 = N11217 & N1190;
  assign N14230 = N11219 & N1190;
  assign N14231 = N11221 & N1190;
  assign N14232 = N11223 & N1190;
  assign N14233 = N11225 & N1190;
  assign N14234 = N11227 & N1190;
  assign N14235 = N11229 & N1190;
  assign N14236 = N11231 & N1190;
  assign N14237 = N11233 & N1190;
  assign N14238 = N11235 & N1190;
  assign N14239 = N11237 & N1190;
  assign N14240 = N11239 & N1190;
  assign N14241 = N11241 & N1190;
  assign N14242 = N11243 & N1190;
  assign N14243 = N11245 & N1190;
  assign N14244 = N11247 & N1190;
  assign N14245 = N11249 & N1190;
  assign N14246 = N11251 & N1190;
  assign N14247 = N11253 & N1190;
  assign N14248 = N11255 & N1190;
  assign N14249 = N11257 & N1190;
  assign N14250 = N11259 & N1190;
  assign N14251 = N11261 & N1190;
  assign N14252 = N11263 & N1190;
  assign N14253 = N11265 & N1190;
  assign N14254 = N11267 & N1190;
  assign N14255 = N11269 & N1190;
  assign N14256 = N11271 & N1190;
  assign N14257 = N11273 & N1190;
  assign N14258 = N11275 & N1190;
  assign N14259 = N11277 & N1190;
  assign N14260 = N11279 & N1190;
  assign N14261 = N11281 & N1190;
  assign N14262 = N11283 & N1190;
  assign N14263 = N11285 & N1190;
  assign N14264 = N11287 & N1190;
  assign N14265 = N11289 & N1190;
  assign N14266 = N11291 & N1190;
  assign N14267 = N11293 & N1190;
  assign N14268 = N11295 & N1190;
  assign N14269 = N11297 & N1190;
  assign N14270 = N11299 & N1190;
  assign N14271 = N11301 & N1190;
  assign N14272 = N11303 & N1190;
  assign N14273 = N11305 & N1190;
  assign N14274 = N11307 & N1190;
  assign N14275 = N11309 & N1190;
  assign N14276 = N11311 & N1190;
  assign N14277 = N11313 & N1190;
  assign N14278 = N11315 & N1190;
  assign N14279 = N11317 & N1190;
  assign N14280 = N11319 & N1190;
  assign N14281 = N11321 & N1190;
  assign N14282 = N11323 & N1190;
  assign N14283 = N11325 & N1190;
  assign N14284 = N11327 & N1190;
  assign N14285 = N11329 & N1190;
  assign N14286 = N11331 & N1190;
  assign N14287 = N11333 & N1190;
  assign N14288 = N11335 & N1190;
  assign N14289 = N11337 & N1190;
  assign N14290 = N11339 & N1190;
  assign N14291 = N11341 & N1190;
  assign N14292 = N11343 & N1190;
  assign N14293 = N14101 & N1415;
  assign N14294 = N14101 & idx_w_i[8];
  assign N14295 = N14103 & N1415;
  assign N14296 = N14103 & idx_w_i[8];
  assign N14297 = N14105 & N1415;
  assign N14298 = N14105 & idx_w_i[8];
  assign N14299 = N14107 & N1415;
  assign N14300 = N14107 & idx_w_i[8];
  assign N14301 = N14109 & N1415;
  assign N14302 = N14109 & idx_w_i[8];
  assign N14303 = N14111 & N1415;
  assign N14304 = N14111 & idx_w_i[8];
  assign N14305 = N14113 & N1415;
  assign N14306 = N14113 & idx_w_i[8];
  assign N14307 = N14115 & N1415;
  assign N14308 = N14115 & idx_w_i[8];
  assign N14309 = N14117 & N1415;
  assign N14310 = N14117 & idx_w_i[8];
  assign N14311 = N14119 & N1415;
  assign N14312 = N14119 & idx_w_i[8];
  assign N14313 = N14121 & N1415;
  assign N14314 = N14121 & idx_w_i[8];
  assign N14315 = N14123 & N1415;
  assign N14316 = N14123 & idx_w_i[8];
  assign N14317 = N14125 & N1415;
  assign N14318 = N14125 & idx_w_i[8];
  assign N14319 = N14127 & N1415;
  assign N14320 = N14127 & idx_w_i[8];
  assign N14321 = N14129 & N1415;
  assign N14322 = N14129 & idx_w_i[8];
  assign N14323 = N14131 & N1415;
  assign N14324 = N14131 & idx_w_i[8];
  assign N14325 = N14133 & N1415;
  assign N14326 = N14133 & idx_w_i[8];
  assign N14327 = N14135 & N1415;
  assign N14328 = N14135 & idx_w_i[8];
  assign N14329 = N14137 & N1415;
  assign N14330 = N14137 & idx_w_i[8];
  assign N14331 = N14139 & N1415;
  assign N14332 = N14139 & idx_w_i[8];
  assign N14333 = N14141 & N1415;
  assign N14334 = N14141 & idx_w_i[8];
  assign N14335 = N14143 & N1415;
  assign N14336 = N14143 & idx_w_i[8];
  assign N14337 = N14145 & N1415;
  assign N14338 = N14145 & idx_w_i[8];
  assign N14339 = N14147 & N1415;
  assign N14340 = N14147 & idx_w_i[8];
  assign N14341 = N14149 & N1415;
  assign N14342 = N14149 & idx_w_i[8];
  assign N14343 = N14151 & N1415;
  assign N14344 = N14151 & idx_w_i[8];
  assign N14345 = N14153 & N1415;
  assign N14346 = N14153 & idx_w_i[8];
  assign N14347 = N14155 & N1415;
  assign N14348 = N14155 & idx_w_i[8];
  assign N14349 = N14157 & N1415;
  assign N14350 = N14157 & idx_w_i[8];
  assign N14351 = N14159 & N1415;
  assign N14352 = N14159 & idx_w_i[8];
  assign N14353 = N14161 & N1415;
  assign N14354 = N14161 & idx_w_i[8];
  assign N14355 = N14163 & N1415;
  assign N14356 = N14163 & idx_w_i[8];
  assign N14357 = N14165 & N1415;
  assign N14358 = N14165 & idx_w_i[8];
  assign N14359 = N14167 & N1415;
  assign N14360 = N14167 & idx_w_i[8];
  assign N14361 = N14169 & N1415;
  assign N14362 = N14169 & idx_w_i[8];
  assign N14363 = N14171 & N1415;
  assign N14364 = N14171 & idx_w_i[8];
  assign N14365 = N14173 & N1415;
  assign N14366 = N14173 & idx_w_i[8];
  assign N14367 = N14175 & N1415;
  assign N14368 = N14175 & idx_w_i[8];
  assign N14369 = N14177 & N1415;
  assign N14370 = N14177 & idx_w_i[8];
  assign N14371 = N14179 & N1415;
  assign N14372 = N14179 & idx_w_i[8];
  assign N14373 = N14181 & N1415;
  assign N14374 = N14181 & idx_w_i[8];
  assign N14375 = N14183 & N1415;
  assign N14376 = N14183 & idx_w_i[8];
  assign N14377 = N14185 & N1415;
  assign N14378 = N14185 & idx_w_i[8];
  assign N14379 = N14187 & N1415;
  assign N14380 = N14187 & idx_w_i[8];
  assign N14381 = N14189 & N1415;
  assign N14382 = N14189 & idx_w_i[8];
  assign N14383 = N14191 & N1415;
  assign N14384 = N14191 & idx_w_i[8];
  assign N14385 = N14193 & N1415;
  assign N14386 = N14193 & idx_w_i[8];
  assign N14387 = N14195 & N1415;
  assign N14388 = N14195 & idx_w_i[8];
  assign N14389 = N14197 & N1415;
  assign N14390 = N14197 & idx_w_i[8];
  assign N14391 = N14199 & N1415;
  assign N14392 = N14199 & idx_w_i[8];
  assign N14393 = N14201 & N1415;
  assign N14394 = N14201 & idx_w_i[8];
  assign N14395 = N14203 & N1415;
  assign N14396 = N14203 & idx_w_i[8];
  assign N14397 = N14205 & N1415;
  assign N14398 = N14205 & idx_w_i[8];
  assign N14399 = N14207 & N1415;
  assign N14400 = N14207 & idx_w_i[8];
  assign N14401 = N14209 & N1415;
  assign N14402 = N14209 & idx_w_i[8];
  assign N14403 = N14211 & N1415;
  assign N14404 = N14211 & idx_w_i[8];
  assign N14405 = N14213 & N1415;
  assign N14406 = N14213 & idx_w_i[8];
  assign N14407 = N14215 & N1415;
  assign N14408 = N14215 & idx_w_i[8];
  assign N14409 = N14217 & N1415;
  assign N14410 = N14217 & idx_w_i[8];
  assign N14411 = N14219 & N1415;
  assign N14412 = N14219 & idx_w_i[8];
  assign N14413 = N14221 & N1415;
  assign N14414 = N14221 & idx_w_i[8];
  assign N14415 = N14223 & N1415;
  assign N14416 = N14223 & idx_w_i[8];
  assign N14417 = N14225 & N1415;
  assign N14418 = N14225 & idx_w_i[8];
  assign N14419 = N14227 & N1415;
  assign N14420 = N14227 & idx_w_i[8];
  assign N14421 = N14229 & N1415;
  assign N14422 = N14229 & idx_w_i[8];
  assign N14423 = N14230 & N1415;
  assign N14424 = N14230 & idx_w_i[8];
  assign N14425 = N14231 & N1415;
  assign N14426 = N14231 & idx_w_i[8];
  assign N14427 = N14232 & N1415;
  assign N14428 = N14232 & idx_w_i[8];
  assign N14429 = N14233 & N1415;
  assign N14430 = N14233 & idx_w_i[8];
  assign N14431 = N14234 & N1415;
  assign N14432 = N14234 & idx_w_i[8];
  assign N14433 = N14235 & N1415;
  assign N14434 = N14235 & idx_w_i[8];
  assign N14435 = N14236 & N1415;
  assign N14436 = N14236 & idx_w_i[8];
  assign N14437 = N14237 & N1415;
  assign N14438 = N14237 & idx_w_i[8];
  assign N14439 = N14238 & N1415;
  assign N14440 = N14238 & idx_w_i[8];
  assign N14441 = N14239 & N1415;
  assign N14442 = N14239 & idx_w_i[8];
  assign N14443 = N14240 & N1415;
  assign N14444 = N14240 & idx_w_i[8];
  assign N14445 = N14241 & N1415;
  assign N14446 = N14241 & idx_w_i[8];
  assign N14447 = N14242 & N1415;
  assign N14448 = N14242 & idx_w_i[8];
  assign N14449 = N14243 & N1415;
  assign N14450 = N14243 & idx_w_i[8];
  assign N14451 = N14244 & N1415;
  assign N14452 = N14244 & idx_w_i[8];
  assign N14453 = N14245 & N1415;
  assign N14454 = N14245 & idx_w_i[8];
  assign N14455 = N14246 & N1415;
  assign N14456 = N14246 & idx_w_i[8];
  assign N14457 = N14247 & N1415;
  assign N14458 = N14247 & idx_w_i[8];
  assign N14459 = N14248 & N1415;
  assign N14460 = N14248 & idx_w_i[8];
  assign N14461 = N14249 & N1415;
  assign N14462 = N14249 & idx_w_i[8];
  assign N14463 = N14250 & N1415;
  assign N14464 = N14250 & idx_w_i[8];
  assign N14465 = N14251 & N1415;
  assign N14466 = N14251 & idx_w_i[8];
  assign N14467 = N14252 & N1415;
  assign N14468 = N14252 & idx_w_i[8];
  assign N14469 = N14253 & N1415;
  assign N14470 = N14253 & idx_w_i[8];
  assign N14471 = N14254 & N1415;
  assign N14472 = N14254 & idx_w_i[8];
  assign N14473 = N14255 & N1415;
  assign N14474 = N14255 & idx_w_i[8];
  assign N14475 = N14256 & N1415;
  assign N14476 = N14256 & idx_w_i[8];
  assign N14477 = N14257 & N1415;
  assign N14478 = N14257 & idx_w_i[8];
  assign N14479 = N14258 & N1415;
  assign N14480 = N14258 & idx_w_i[8];
  assign N14481 = N14259 & N1415;
  assign N14482 = N14259 & idx_w_i[8];
  assign N14483 = N14260 & N1415;
  assign N14484 = N14260 & idx_w_i[8];
  assign N14485 = N14261 & N1415;
  assign N14486 = N14261 & idx_w_i[8];
  assign N14487 = N14262 & N1415;
  assign N14488 = N14262 & idx_w_i[8];
  assign N14489 = N14263 & N1415;
  assign N14490 = N14263 & idx_w_i[8];
  assign N14491 = N14264 & N1415;
  assign N14492 = N14264 & idx_w_i[8];
  assign N14493 = N14265 & N1415;
  assign N14494 = N14265 & idx_w_i[8];
  assign N14495 = N14266 & N1415;
  assign N14496 = N14266 & idx_w_i[8];
  assign N14497 = N14267 & N1415;
  assign N14498 = N14267 & idx_w_i[8];
  assign N14499 = N14268 & N1415;
  assign N14500 = N14268 & idx_w_i[8];
  assign N14501 = N14269 & N1415;
  assign N14502 = N14269 & idx_w_i[8];
  assign N14503 = N14270 & N1415;
  assign N14504 = N14270 & idx_w_i[8];
  assign N14505 = N14271 & N1415;
  assign N14506 = N14271 & idx_w_i[8];
  assign N14507 = N14272 & N1415;
  assign N14508 = N14272 & idx_w_i[8];
  assign N14509 = N14273 & N1415;
  assign N14510 = N14273 & idx_w_i[8];
  assign N14511 = N14274 & N1415;
  assign N14512 = N14274 & idx_w_i[8];
  assign N14513 = N14275 & N1415;
  assign N14514 = N14275 & idx_w_i[8];
  assign N14515 = N14276 & N1415;
  assign N14516 = N14276 & idx_w_i[8];
  assign N14517 = N14277 & N1415;
  assign N14518 = N14277 & idx_w_i[8];
  assign N14519 = N14278 & N1415;
  assign N14520 = N14278 & idx_w_i[8];
  assign N14521 = N14279 & N1415;
  assign N14522 = N14279 & idx_w_i[8];
  assign N14523 = N14280 & N1415;
  assign N14524 = N14280 & idx_w_i[8];
  assign N14525 = N14281 & N1415;
  assign N14526 = N14281 & idx_w_i[8];
  assign N14527 = N14282 & N1415;
  assign N14528 = N14282 & idx_w_i[8];
  assign N14529 = N14283 & N1415;
  assign N14530 = N14283 & idx_w_i[8];
  assign N14531 = N14284 & N1415;
  assign N14532 = N14284 & idx_w_i[8];
  assign N14533 = N14285 & N1415;
  assign N14534 = N14285 & idx_w_i[8];
  assign N14535 = N14286 & N1415;
  assign N14536 = N14286 & idx_w_i[8];
  assign N14537 = N14287 & N1415;
  assign N14538 = N14287 & idx_w_i[8];
  assign N14539 = N14288 & N1415;
  assign N14540 = N14288 & idx_w_i[8];
  assign N14541 = N14289 & N1415;
  assign N14542 = N14289 & idx_w_i[8];
  assign N14543 = N14290 & N1415;
  assign N14544 = N14290 & idx_w_i[8];
  assign N14545 = N14291 & N1415;
  assign N14546 = N14291 & idx_w_i[8];
  assign N14547 = N14292 & N1415;
  assign N14548 = N14292 & idx_w_i[8];
  assign N14549 = N14102 & N1415;
  assign N14550 = N14102 & idx_w_i[8];
  assign N14551 = N14104 & N1415;
  assign N14552 = N14104 & idx_w_i[8];
  assign N14553 = N14106 & N1415;
  assign N14554 = N14106 & idx_w_i[8];
  assign N14555 = N14108 & N1415;
  assign N14556 = N14108 & idx_w_i[8];
  assign N14557 = N14110 & N1415;
  assign N14558 = N14110 & idx_w_i[8];
  assign N14559 = N14112 & N1415;
  assign N14560 = N14112 & idx_w_i[8];
  assign N14561 = N14114 & N1415;
  assign N14562 = N14114 & idx_w_i[8];
  assign N14563 = N14116 & N1415;
  assign N14564 = N14116 & idx_w_i[8];
  assign N14565 = N14118 & N1415;
  assign N14566 = N14118 & idx_w_i[8];
  assign N14567 = N14120 & N1415;
  assign N14568 = N14120 & idx_w_i[8];
  assign N14569 = N14122 & N1415;
  assign N14570 = N14122 & idx_w_i[8];
  assign N14571 = N14124 & N1415;
  assign N14572 = N14124 & idx_w_i[8];
  assign N14573 = N14126 & N1415;
  assign N14574 = N14126 & idx_w_i[8];
  assign N14575 = N14128 & N1415;
  assign N14576 = N14128 & idx_w_i[8];
  assign N14577 = N14130 & N1415;
  assign N14578 = N14130 & idx_w_i[8];
  assign N14579 = N14132 & N1415;
  assign N14580 = N14132 & idx_w_i[8];
  assign N14581 = N14134 & N1415;
  assign N14582 = N14134 & idx_w_i[8];
  assign N14583 = N14136 & N1415;
  assign N14584 = N14136 & idx_w_i[8];
  assign N14585 = N14138 & N1415;
  assign N14586 = N14138 & idx_w_i[8];
  assign N14587 = N14140 & N1415;
  assign N14588 = N14140 & idx_w_i[8];
  assign N14589 = N14142 & N1415;
  assign N14590 = N14142 & idx_w_i[8];
  assign N14591 = N14144 & N1415;
  assign N14592 = N14144 & idx_w_i[8];
  assign N14593 = N14146 & N1415;
  assign N14594 = N14146 & idx_w_i[8];
  assign N14595 = N14148 & N1415;
  assign N14596 = N14148 & idx_w_i[8];
  assign N14597 = N14150 & N1415;
  assign N14598 = N14150 & idx_w_i[8];
  assign N14599 = N14152 & N1415;
  assign N14600 = N14152 & idx_w_i[8];
  assign N14601 = N14154 & N1415;
  assign N14602 = N14154 & idx_w_i[8];
  assign N14603 = N14156 & N1415;
  assign N14604 = N14156 & idx_w_i[8];
  assign N14605 = N14158 & N1415;
  assign N14606 = N14158 & idx_w_i[8];
  assign N14607 = N14160 & N1415;
  assign N14608 = N14160 & idx_w_i[8];
  assign N14609 = N14162 & N1415;
  assign N14610 = N14162 & idx_w_i[8];
  assign N14611 = N14164 & N1415;
  assign N14612 = N14164 & idx_w_i[8];
  assign N14613 = N14166 & N1415;
  assign N14614 = N14166 & idx_w_i[8];
  assign N14615 = N14168 & N1415;
  assign N14616 = N14168 & idx_w_i[8];
  assign N14617 = N14170 & N1415;
  assign N14618 = N14170 & idx_w_i[8];
  assign N14619 = N14172 & N1415;
  assign N14620 = N14172 & idx_w_i[8];
  assign N14621 = N14174 & N1415;
  assign N14622 = N14174 & idx_w_i[8];
  assign N14623 = N14176 & N1415;
  assign N14624 = N14176 & idx_w_i[8];
  assign N14625 = N14178 & N1415;
  assign N14626 = N14178 & idx_w_i[8];
  assign N14627 = N14180 & N1415;
  assign N14628 = N14180 & idx_w_i[8];
  assign N14629 = N14182 & N1415;
  assign N14630 = N14182 & idx_w_i[8];
  assign N14631 = N14184 & N1415;
  assign N14632 = N14184 & idx_w_i[8];
  assign N14633 = N14186 & N1415;
  assign N14634 = N14186 & idx_w_i[8];
  assign N14635 = N14188 & N1415;
  assign N14636 = N14188 & idx_w_i[8];
  assign N14637 = N14190 & N1415;
  assign N14638 = N14190 & idx_w_i[8];
  assign N14639 = N14192 & N1415;
  assign N14640 = N14192 & idx_w_i[8];
  assign N14641 = N14194 & N1415;
  assign N14642 = N14194 & idx_w_i[8];
  assign N14643 = N14196 & N1415;
  assign N14644 = N14196 & idx_w_i[8];
  assign N14645 = N14198 & N1415;
  assign N14646 = N14198 & idx_w_i[8];
  assign N14647 = N14200 & N1415;
  assign N14648 = N14200 & idx_w_i[8];
  assign N14649 = N14202 & N1415;
  assign N14650 = N14202 & idx_w_i[8];
  assign N14651 = N14204 & N1415;
  assign N14652 = N14204 & idx_w_i[8];
  assign N14653 = N14206 & N1415;
  assign N14654 = N14206 & idx_w_i[8];
  assign N14655 = N14208 & N1415;
  assign N14656 = N14208 & idx_w_i[8];
  assign N14657 = N14210 & N1415;
  assign N14658 = N14210 & idx_w_i[8];
  assign N14659 = N14212 & N1415;
  assign N14660 = N14212 & idx_w_i[8];
  assign N14661 = N14214 & N1415;
  assign N14662 = N14214 & idx_w_i[8];
  assign N14663 = N14216 & N1415;
  assign N14664 = N14216 & idx_w_i[8];
  assign N14665 = N14218 & N1415;
  assign N14666 = N14218 & idx_w_i[8];
  assign N14667 = N14220 & N1415;
  assign N14668 = N14220 & idx_w_i[8];
  assign N14669 = N14222 & N1415;
  assign N14670 = N14222 & idx_w_i[8];
  assign N14671 = N14224 & N1415;
  assign N14672 = N14224 & idx_w_i[8];
  assign N14673 = N14226 & N1415;
  assign N14674 = N14226 & idx_w_i[8];
  assign N14675 = N14228 & N1415;
  assign N14676 = N14228 & idx_w_i[8];
  assign N14677 = N11473 & N1415;
  assign N14678 = N11475 & N1415;
  assign N14679 = N11477 & N1415;
  assign N14680 = N11479 & N1415;
  assign N14681 = N11481 & N1415;
  assign N14682 = N11483 & N1415;
  assign N14683 = N11485 & N1415;
  assign N14684 = N11487 & N1415;
  assign N14685 = N11489 & N1415;
  assign N14686 = N11491 & N1415;
  assign N14687 = N11493 & N1415;
  assign N14688 = N11495 & N1415;
  assign N14689 = N11497 & N1415;
  assign N14690 = N11499 & N1415;
  assign N14691 = N11501 & N1415;
  assign N14692 = N11503 & N1415;
  assign N14693 = N11505 & N1415;
  assign N14694 = N11507 & N1415;
  assign N14695 = N11509 & N1415;
  assign N14696 = N11511 & N1415;
  assign N14697 = N11513 & N1415;
  assign N14698 = N11515 & N1415;
  assign N14699 = N11517 & N1415;
  assign N14700 = N11519 & N1415;
  assign N14701 = N11521 & N1415;
  assign N14702 = N11523 & N1415;
  assign N14703 = N11525 & N1415;
  assign N14704 = N11527 & N1415;
  assign N14705 = N11529 & N1415;
  assign N14706 = N11531 & N1415;
  assign N14707 = N11533 & N1415;
  assign N14708 = N11535 & N1415;
  assign N14709 = N11537 & N1415;
  assign N14710 = N11539 & N1415;
  assign N14711 = N11541 & N1415;
  assign N14712 = N11543 & N1415;
  assign N14713 = N11545 & N1415;
  assign N14714 = N11547 & N1415;
  assign N14715 = N11549 & N1415;
  assign N14716 = N11551 & N1415;
  assign N14717 = N11553 & N1415;
  assign N14718 = N11555 & N1415;
  assign N14719 = N11557 & N1415;
  assign N14720 = N11559 & N1415;
  assign N14721 = N11561 & N1415;
  assign N14722 = N11563 & N1415;
  assign N14723 = N11565 & N1415;
  assign N14724 = N11567 & N1415;
  assign N14725 = N11569 & N1415;
  assign N14726 = N11571 & N1415;
  assign N14727 = N11573 & N1415;
  assign N14728 = N11575 & N1415;
  assign N14729 = N11577 & N1415;
  assign N14730 = N11579 & N1415;
  assign N14731 = N11581 & N1415;
  assign N14732 = N11583 & N1415;
  assign N14733 = N11585 & N1415;
  assign N14734 = N11587 & N1415;
  assign N14735 = N11589 & N1415;
  assign N14736 = N11591 & N1415;
  assign N14737 = N11593 & N1415;
  assign N14738 = N11595 & N1415;
  assign N14739 = N11597 & N1415;
  assign N14740 = N11599 & N1415;
  assign N14742 = N11152 & N1093;
  assign N14743 = N11154 & N1093;
  assign N14744 = N11156 & N1093;
  assign N14745 = N11158 & N1093;
  assign N14746 = N11160 & N1093;
  assign N14747 = N11162 & N1093;
  assign N14748 = N11164 & N1093;
  assign N14749 = N11166 & N1093;
  assign N14750 = N11168 & N1093;
  assign N14751 = N11170 & N1093;
  assign N14752 = N11172 & N1093;
  assign N14753 = N11174 & N1093;
  assign N14754 = N11176 & N1093;
  assign N14755 = N11178 & N1093;
  assign N14756 = N11180 & N1093;
  assign N14757 = N11182 & N1093;
  assign N14758 = N11184 & N1093;
  assign N14759 = N11186 & N1093;
  assign N14760 = N11188 & N1093;
  assign N14761 = N11190 & N1093;
  assign N14762 = N11192 & N1093;
  assign N14763 = N11194 & N1093;
  assign N14764 = N11196 & N1093;
  assign N14765 = N11198 & N1093;
  assign N14766 = N11200 & N1093;
  assign N14767 = N11202 & N1093;
  assign N14768 = N11204 & N1093;
  assign N14769 = N11206 & N1093;
  assign N14770 = N11208 & N1093;
  assign N14771 = N11210 & N1093;
  assign N14772 = N11212 & N1093;
  assign N14773 = N11214 & N1093;
  assign N14774 = N11153 & N1093;
  assign N14775 = N11155 & N1093;
  assign N14776 = N11157 & N1093;
  assign N14777 = N11159 & N1093;
  assign N14778 = N11161 & N1093;
  assign N14779 = N11163 & N1093;
  assign N14780 = N11165 & N1093;
  assign N14781 = N11167 & N1093;
  assign N14782 = N11169 & N1093;
  assign N14783 = N11171 & N1093;
  assign N14784 = N11173 & N1093;
  assign N14785 = N11175 & N1093;
  assign N14786 = N11177 & N1093;
  assign N14787 = N11179 & N1093;
  assign N14788 = N11181 & N1093;
  assign N14789 = N11183 & N1093;
  assign N14790 = N11185 & N1093;
  assign N14791 = N11187 & N1093;
  assign N14792 = N11189 & N1093;
  assign N14793 = N11191 & N1093;
  assign N14794 = N11193 & N1093;
  assign N14795 = N11195 & N1093;
  assign N14796 = N11197 & N1093;
  assign N14797 = N11199 & N1093;
  assign N14798 = N11201 & N1093;
  assign N14799 = N11203 & N1093;
  assign N14800 = N11205 & N1093;
  assign N14801 = N11207 & N1093;
  assign N14802 = N11209 & N1093;
  assign N14803 = N11211 & N1093;
  assign N14804 = N11213 & N1093;
  assign N14805 = N11215 & N1093;
  assign N14806 = N14742 & N1190;
  assign N14807 = N14742 & idx_w_i[7];
  assign N14808 = N14743 & N1190;
  assign N14809 = N14743 & idx_w_i[7];
  assign N14810 = N14744 & N1190;
  assign N14811 = N14744 & idx_w_i[7];
  assign N14812 = N14745 & N1190;
  assign N14813 = N14745 & idx_w_i[7];
  assign N14814 = N14746 & N1190;
  assign N14815 = N14746 & idx_w_i[7];
  assign N14816 = N14747 & N1190;
  assign N14817 = N14747 & idx_w_i[7];
  assign N14818 = N14748 & N1190;
  assign N14819 = N14748 & idx_w_i[7];
  assign N14820 = N14749 & N1190;
  assign N14821 = N14749 & idx_w_i[7];
  assign N14822 = N14750 & N1190;
  assign N14823 = N14750 & idx_w_i[7];
  assign N14824 = N14751 & N1190;
  assign N14825 = N14751 & idx_w_i[7];
  assign N14826 = N14752 & N1190;
  assign N14827 = N14752 & idx_w_i[7];
  assign N14828 = N14753 & N1190;
  assign N14829 = N14753 & idx_w_i[7];
  assign N14830 = N14754 & N1190;
  assign N14831 = N14754 & idx_w_i[7];
  assign N14832 = N14755 & N1190;
  assign N14833 = N14755 & idx_w_i[7];
  assign N14834 = N14756 & N1190;
  assign N14835 = N14756 & idx_w_i[7];
  assign N14836 = N14757 & N1190;
  assign N14837 = N14757 & idx_w_i[7];
  assign N14838 = N14758 & N1190;
  assign N14839 = N14758 & idx_w_i[7];
  assign N14840 = N14759 & N1190;
  assign N14841 = N14759 & idx_w_i[7];
  assign N14842 = N14760 & N1190;
  assign N14843 = N14760 & idx_w_i[7];
  assign N14844 = N14761 & N1190;
  assign N14845 = N14761 & idx_w_i[7];
  assign N14846 = N14762 & N1190;
  assign N14847 = N14762 & idx_w_i[7];
  assign N14848 = N14763 & N1190;
  assign N14849 = N14763 & idx_w_i[7];
  assign N14850 = N14764 & N1190;
  assign N14851 = N14764 & idx_w_i[7];
  assign N14852 = N14765 & N1190;
  assign N14853 = N14765 & idx_w_i[7];
  assign N14854 = N14766 & N1190;
  assign N14855 = N14766 & idx_w_i[7];
  assign N14856 = N14767 & N1190;
  assign N14857 = N14767 & idx_w_i[7];
  assign N14858 = N14768 & N1190;
  assign N14859 = N14768 & idx_w_i[7];
  assign N14860 = N14769 & N1190;
  assign N14861 = N14769 & idx_w_i[7];
  assign N14862 = N14770 & N1190;
  assign N14863 = N14770 & idx_w_i[7];
  assign N14864 = N14771 & N1190;
  assign N14865 = N14771 & idx_w_i[7];
  assign N14866 = N14772 & N1190;
  assign N14867 = N14772 & idx_w_i[7];
  assign N14868 = N14773 & N1190;
  assign N14869 = N14773 & idx_w_i[7];
  assign N14870 = N14774 & N1190;
  assign N14871 = N14774 & idx_w_i[7];
  assign N14872 = N14775 & N1190;
  assign N14873 = N14775 & idx_w_i[7];
  assign N14874 = N14776 & N1190;
  assign N14875 = N14776 & idx_w_i[7];
  assign N14876 = N14777 & N1190;
  assign N14877 = N14777 & idx_w_i[7];
  assign N14878 = N14778 & N1190;
  assign N14879 = N14778 & idx_w_i[7];
  assign N14880 = N14779 & N1190;
  assign N14881 = N14779 & idx_w_i[7];
  assign N14882 = N14780 & N1190;
  assign N14883 = N14780 & idx_w_i[7];
  assign N14884 = N14781 & N1190;
  assign N14885 = N14781 & idx_w_i[7];
  assign N14886 = N14782 & N1190;
  assign N14887 = N14782 & idx_w_i[7];
  assign N14888 = N14783 & N1190;
  assign N14889 = N14783 & idx_w_i[7];
  assign N14890 = N14784 & N1190;
  assign N14891 = N14784 & idx_w_i[7];
  assign N14892 = N14785 & N1190;
  assign N14893 = N14785 & idx_w_i[7];
  assign N14894 = N14786 & N1190;
  assign N14895 = N14786 & idx_w_i[7];
  assign N14896 = N14787 & N1190;
  assign N14897 = N14787 & idx_w_i[7];
  assign N14898 = N14788 & N1190;
  assign N14899 = N14788 & idx_w_i[7];
  assign N14900 = N14789 & N1190;
  assign N14901 = N14789 & idx_w_i[7];
  assign N14902 = N14790 & N1190;
  assign N14903 = N14790 & idx_w_i[7];
  assign N14904 = N14791 & N1190;
  assign N14905 = N14791 & idx_w_i[7];
  assign N14906 = N14792 & N1190;
  assign N14907 = N14792 & idx_w_i[7];
  assign N14908 = N14793 & N1190;
  assign N14909 = N14793 & idx_w_i[7];
  assign N14910 = N14794 & N1190;
  assign N14911 = N14794 & idx_w_i[7];
  assign N14912 = N14795 & N1190;
  assign N14913 = N14795 & idx_w_i[7];
  assign N14914 = N14796 & N1190;
  assign N14915 = N14796 & idx_w_i[7];
  assign N14916 = N14797 & N1190;
  assign N14917 = N14797 & idx_w_i[7];
  assign N14918 = N14798 & N1190;
  assign N14919 = N14798 & idx_w_i[7];
  assign N14920 = N14799 & N1190;
  assign N14921 = N14799 & idx_w_i[7];
  assign N14922 = N14800 & N1190;
  assign N14923 = N14800 & idx_w_i[7];
  assign N14924 = N14801 & N1190;
  assign N14925 = N14801 & idx_w_i[7];
  assign N14926 = N14802 & N1190;
  assign N14927 = N14802 & idx_w_i[7];
  assign N14928 = N14803 & N1190;
  assign N14929 = N14803 & idx_w_i[7];
  assign N14930 = N14804 & N1190;
  assign N14931 = N14804 & idx_w_i[7];
  assign N14932 = N14805 & N1190;
  assign N14933 = N14805 & idx_w_i[7];
  assign N14934 = N11217 & N1190;
  assign N14935 = N11219 & N1190;
  assign N14936 = N11221 & N1190;
  assign N14937 = N11223 & N1190;
  assign N14938 = N11225 & N1190;
  assign N14939 = N11227 & N1190;
  assign N14940 = N11229 & N1190;
  assign N14941 = N11231 & N1190;
  assign N14942 = N11233 & N1190;
  assign N14943 = N11235 & N1190;
  assign N14944 = N11237 & N1190;
  assign N14945 = N11239 & N1190;
  assign N14946 = N11241 & N1190;
  assign N14947 = N11243 & N1190;
  assign N14948 = N11245 & N1190;
  assign N14949 = N11247 & N1190;
  assign N14950 = N11249 & N1190;
  assign N14951 = N11251 & N1190;
  assign N14952 = N11253 & N1190;
  assign N14953 = N11255 & N1190;
  assign N14954 = N11257 & N1190;
  assign N14955 = N11259 & N1190;
  assign N14956 = N11261 & N1190;
  assign N14957 = N11263 & N1190;
  assign N14958 = N11265 & N1190;
  assign N14959 = N11267 & N1190;
  assign N14960 = N11269 & N1190;
  assign N14961 = N11271 & N1190;
  assign N14962 = N11273 & N1190;
  assign N14963 = N11275 & N1190;
  assign N14964 = N11277 & N1190;
  assign N14965 = N11279 & N1190;
  assign N14966 = N11281 & N1190;
  assign N14967 = N11283 & N1190;
  assign N14968 = N11285 & N1190;
  assign N14969 = N11287 & N1190;
  assign N14970 = N11289 & N1190;
  assign N14971 = N11291 & N1190;
  assign N14972 = N11293 & N1190;
  assign N14973 = N11295 & N1190;
  assign N14974 = N11297 & N1190;
  assign N14975 = N11299 & N1190;
  assign N14976 = N11301 & N1190;
  assign N14977 = N11303 & N1190;
  assign N14978 = N11305 & N1190;
  assign N14979 = N11307 & N1190;
  assign N14980 = N11309 & N1190;
  assign N14981 = N11311 & N1190;
  assign N14982 = N11313 & N1190;
  assign N14983 = N11315 & N1190;
  assign N14984 = N11317 & N1190;
  assign N14985 = N11319 & N1190;
  assign N14986 = N11321 & N1190;
  assign N14987 = N11323 & N1190;
  assign N14988 = N11325 & N1190;
  assign N14989 = N11327 & N1190;
  assign N14990 = N11329 & N1190;
  assign N14991 = N11331 & N1190;
  assign N14992 = N11333 & N1190;
  assign N14993 = N11335 & N1190;
  assign N14994 = N11337 & N1190;
  assign N14995 = N11339 & N1190;
  assign N14996 = N11341 & N1190;
  assign N14997 = N11343 & N1190;
  assign N14998 = N14806 & N1415;
  assign N14999 = N14806 & idx_w_i[8];
  assign N15000 = N14808 & N1415;
  assign N15001 = N14808 & idx_w_i[8];
  assign N15002 = N14810 & N1415;
  assign N15003 = N14810 & idx_w_i[8];
  assign N15004 = N14812 & N1415;
  assign N15005 = N14812 & idx_w_i[8];
  assign N15006 = N14814 & N1415;
  assign N15007 = N14814 & idx_w_i[8];
  assign N15008 = N14816 & N1415;
  assign N15009 = N14816 & idx_w_i[8];
  assign N15010 = N14818 & N1415;
  assign N15011 = N14818 & idx_w_i[8];
  assign N15012 = N14820 & N1415;
  assign N15013 = N14820 & idx_w_i[8];
  assign N15014 = N14822 & N1415;
  assign N15015 = N14822 & idx_w_i[8];
  assign N15016 = N14824 & N1415;
  assign N15017 = N14824 & idx_w_i[8];
  assign N15018 = N14826 & N1415;
  assign N15019 = N14826 & idx_w_i[8];
  assign N15020 = N14828 & N1415;
  assign N15021 = N14828 & idx_w_i[8];
  assign N15022 = N14830 & N1415;
  assign N15023 = N14830 & idx_w_i[8];
  assign N15024 = N14832 & N1415;
  assign N15025 = N14832 & idx_w_i[8];
  assign N15026 = N14834 & N1415;
  assign N15027 = N14834 & idx_w_i[8];
  assign N15028 = N14836 & N1415;
  assign N15029 = N14836 & idx_w_i[8];
  assign N15030 = N14838 & N1415;
  assign N15031 = N14838 & idx_w_i[8];
  assign N15032 = N14840 & N1415;
  assign N15033 = N14840 & idx_w_i[8];
  assign N15034 = N14842 & N1415;
  assign N15035 = N14842 & idx_w_i[8];
  assign N15036 = N14844 & N1415;
  assign N15037 = N14844 & idx_w_i[8];
  assign N15038 = N14846 & N1415;
  assign N15039 = N14846 & idx_w_i[8];
  assign N15040 = N14848 & N1415;
  assign N15041 = N14848 & idx_w_i[8];
  assign N15042 = N14850 & N1415;
  assign N15043 = N14850 & idx_w_i[8];
  assign N15044 = N14852 & N1415;
  assign N15045 = N14852 & idx_w_i[8];
  assign N15046 = N14854 & N1415;
  assign N15047 = N14854 & idx_w_i[8];
  assign N15048 = N14856 & N1415;
  assign N15049 = N14856 & idx_w_i[8];
  assign N15050 = N14858 & N1415;
  assign N15051 = N14858 & idx_w_i[8];
  assign N15052 = N14860 & N1415;
  assign N15053 = N14860 & idx_w_i[8];
  assign N15054 = N14862 & N1415;
  assign N15055 = N14862 & idx_w_i[8];
  assign N15056 = N14864 & N1415;
  assign N15057 = N14864 & idx_w_i[8];
  assign N15058 = N14866 & N1415;
  assign N15059 = N14866 & idx_w_i[8];
  assign N15060 = N14868 & N1415;
  assign N15061 = N14868 & idx_w_i[8];
  assign N15062 = N14870 & N1415;
  assign N15063 = N14870 & idx_w_i[8];
  assign N15064 = N14872 & N1415;
  assign N15065 = N14872 & idx_w_i[8];
  assign N15066 = N14874 & N1415;
  assign N15067 = N14874 & idx_w_i[8];
  assign N15068 = N14876 & N1415;
  assign N15069 = N14876 & idx_w_i[8];
  assign N15070 = N14878 & N1415;
  assign N15071 = N14878 & idx_w_i[8];
  assign N15072 = N14880 & N1415;
  assign N15073 = N14880 & idx_w_i[8];
  assign N15074 = N14882 & N1415;
  assign N15075 = N14882 & idx_w_i[8];
  assign N15076 = N14884 & N1415;
  assign N15077 = N14884 & idx_w_i[8];
  assign N15078 = N14886 & N1415;
  assign N15079 = N14886 & idx_w_i[8];
  assign N15080 = N14888 & N1415;
  assign N15081 = N14888 & idx_w_i[8];
  assign N15082 = N14890 & N1415;
  assign N15083 = N14890 & idx_w_i[8];
  assign N15084 = N14892 & N1415;
  assign N15085 = N14892 & idx_w_i[8];
  assign N15086 = N14894 & N1415;
  assign N15087 = N14894 & idx_w_i[8];
  assign N15088 = N14896 & N1415;
  assign N15089 = N14896 & idx_w_i[8];
  assign N15090 = N14898 & N1415;
  assign N15091 = N14898 & idx_w_i[8];
  assign N15092 = N14900 & N1415;
  assign N15093 = N14900 & idx_w_i[8];
  assign N15094 = N14902 & N1415;
  assign N15095 = N14902 & idx_w_i[8];
  assign N15096 = N14904 & N1415;
  assign N15097 = N14904 & idx_w_i[8];
  assign N15098 = N14906 & N1415;
  assign N15099 = N14906 & idx_w_i[8];
  assign N15100 = N14908 & N1415;
  assign N15101 = N14908 & idx_w_i[8];
  assign N15102 = N14910 & N1415;
  assign N15103 = N14910 & idx_w_i[8];
  assign N15104 = N14912 & N1415;
  assign N15105 = N14912 & idx_w_i[8];
  assign N15106 = N14914 & N1415;
  assign N15107 = N14914 & idx_w_i[8];
  assign N15108 = N14916 & N1415;
  assign N15109 = N14916 & idx_w_i[8];
  assign N15110 = N14918 & N1415;
  assign N15111 = N14918 & idx_w_i[8];
  assign N15112 = N14920 & N1415;
  assign N15113 = N14920 & idx_w_i[8];
  assign N15114 = N14922 & N1415;
  assign N15115 = N14922 & idx_w_i[8];
  assign N15116 = N14924 & N1415;
  assign N15117 = N14924 & idx_w_i[8];
  assign N15118 = N14926 & N1415;
  assign N15119 = N14926 & idx_w_i[8];
  assign N15120 = N14928 & N1415;
  assign N15121 = N14928 & idx_w_i[8];
  assign N15122 = N14930 & N1415;
  assign N15123 = N14930 & idx_w_i[8];
  assign N15124 = N14932 & N1415;
  assign N15125 = N14932 & idx_w_i[8];
  assign N15126 = N14934 & N1415;
  assign N15127 = N14934 & idx_w_i[8];
  assign N15128 = N14935 & N1415;
  assign N15129 = N14935 & idx_w_i[8];
  assign N15130 = N14936 & N1415;
  assign N15131 = N14936 & idx_w_i[8];
  assign N15132 = N14937 & N1415;
  assign N15133 = N14937 & idx_w_i[8];
  assign N15134 = N14938 & N1415;
  assign N15135 = N14938 & idx_w_i[8];
  assign N15136 = N14939 & N1415;
  assign N15137 = N14939 & idx_w_i[8];
  assign N15138 = N14940 & N1415;
  assign N15139 = N14940 & idx_w_i[8];
  assign N15140 = N14941 & N1415;
  assign N15141 = N14941 & idx_w_i[8];
  assign N15142 = N14942 & N1415;
  assign N15143 = N14942 & idx_w_i[8];
  assign N15144 = N14943 & N1415;
  assign N15145 = N14943 & idx_w_i[8];
  assign N15146 = N14944 & N1415;
  assign N15147 = N14944 & idx_w_i[8];
  assign N15148 = N14945 & N1415;
  assign N15149 = N14945 & idx_w_i[8];
  assign N15150 = N14946 & N1415;
  assign N15151 = N14946 & idx_w_i[8];
  assign N15152 = N14947 & N1415;
  assign N15153 = N14947 & idx_w_i[8];
  assign N15154 = N14948 & N1415;
  assign N15155 = N14948 & idx_w_i[8];
  assign N15156 = N14949 & N1415;
  assign N15157 = N14949 & idx_w_i[8];
  assign N15158 = N14950 & N1415;
  assign N15159 = N14950 & idx_w_i[8];
  assign N15160 = N14951 & N1415;
  assign N15161 = N14951 & idx_w_i[8];
  assign N15162 = N14952 & N1415;
  assign N15163 = N14952 & idx_w_i[8];
  assign N15164 = N14953 & N1415;
  assign N15165 = N14953 & idx_w_i[8];
  assign N15166 = N14954 & N1415;
  assign N15167 = N14954 & idx_w_i[8];
  assign N15168 = N14955 & N1415;
  assign N15169 = N14955 & idx_w_i[8];
  assign N15170 = N14956 & N1415;
  assign N15171 = N14956 & idx_w_i[8];
  assign N15172 = N14957 & N1415;
  assign N15173 = N14957 & idx_w_i[8];
  assign N15174 = N14958 & N1415;
  assign N15175 = N14958 & idx_w_i[8];
  assign N15176 = N14959 & N1415;
  assign N15177 = N14959 & idx_w_i[8];
  assign N15178 = N14960 & N1415;
  assign N15179 = N14960 & idx_w_i[8];
  assign N15180 = N14961 & N1415;
  assign N15181 = N14961 & idx_w_i[8];
  assign N15182 = N14962 & N1415;
  assign N15183 = N14962 & idx_w_i[8];
  assign N15184 = N14963 & N1415;
  assign N15185 = N14963 & idx_w_i[8];
  assign N15186 = N14964 & N1415;
  assign N15187 = N14964 & idx_w_i[8];
  assign N15188 = N14965 & N1415;
  assign N15189 = N14965 & idx_w_i[8];
  assign N15190 = N14966 & N1415;
  assign N15191 = N14966 & idx_w_i[8];
  assign N15192 = N14967 & N1415;
  assign N15193 = N14967 & idx_w_i[8];
  assign N15194 = N14968 & N1415;
  assign N15195 = N14968 & idx_w_i[8];
  assign N15196 = N14969 & N1415;
  assign N15197 = N14969 & idx_w_i[8];
  assign N15198 = N14970 & N1415;
  assign N15199 = N14970 & idx_w_i[8];
  assign N15200 = N14971 & N1415;
  assign N15201 = N14971 & idx_w_i[8];
  assign N15202 = N14972 & N1415;
  assign N15203 = N14972 & idx_w_i[8];
  assign N15204 = N14973 & N1415;
  assign N15205 = N14973 & idx_w_i[8];
  assign N15206 = N14974 & N1415;
  assign N15207 = N14974 & idx_w_i[8];
  assign N15208 = N14975 & N1415;
  assign N15209 = N14975 & idx_w_i[8];
  assign N15210 = N14976 & N1415;
  assign N15211 = N14976 & idx_w_i[8];
  assign N15212 = N14977 & N1415;
  assign N15213 = N14977 & idx_w_i[8];
  assign N15214 = N14978 & N1415;
  assign N15215 = N14978 & idx_w_i[8];
  assign N15216 = N14979 & N1415;
  assign N15217 = N14979 & idx_w_i[8];
  assign N15218 = N14980 & N1415;
  assign N15219 = N14980 & idx_w_i[8];
  assign N15220 = N14981 & N1415;
  assign N15221 = N14981 & idx_w_i[8];
  assign N15222 = N14982 & N1415;
  assign N15223 = N14982 & idx_w_i[8];
  assign N15224 = N14983 & N1415;
  assign N15225 = N14983 & idx_w_i[8];
  assign N15226 = N14984 & N1415;
  assign N15227 = N14984 & idx_w_i[8];
  assign N15228 = N14985 & N1415;
  assign N15229 = N14985 & idx_w_i[8];
  assign N15230 = N14986 & N1415;
  assign N15231 = N14986 & idx_w_i[8];
  assign N15232 = N14987 & N1415;
  assign N15233 = N14987 & idx_w_i[8];
  assign N15234 = N14988 & N1415;
  assign N15235 = N14988 & idx_w_i[8];
  assign N15236 = N14989 & N1415;
  assign N15237 = N14989 & idx_w_i[8];
  assign N15238 = N14990 & N1415;
  assign N15239 = N14990 & idx_w_i[8];
  assign N15240 = N14991 & N1415;
  assign N15241 = N14991 & idx_w_i[8];
  assign N15242 = N14992 & N1415;
  assign N15243 = N14992 & idx_w_i[8];
  assign N15244 = N14993 & N1415;
  assign N15245 = N14993 & idx_w_i[8];
  assign N15246 = N14994 & N1415;
  assign N15247 = N14994 & idx_w_i[8];
  assign N15248 = N14995 & N1415;
  assign N15249 = N14995 & idx_w_i[8];
  assign N15250 = N14996 & N1415;
  assign N15251 = N14996 & idx_w_i[8];
  assign N15252 = N14997 & N1415;
  assign N15253 = N14997 & idx_w_i[8];
  assign N15254 = N14807 & N1415;
  assign N15255 = N14807 & idx_w_i[8];
  assign N15256 = N14809 & N1415;
  assign N15257 = N14809 & idx_w_i[8];
  assign N15258 = N14811 & N1415;
  assign N15259 = N14811 & idx_w_i[8];
  assign N15260 = N14813 & N1415;
  assign N15261 = N14813 & idx_w_i[8];
  assign N15262 = N14815 & N1415;
  assign N15263 = N14815 & idx_w_i[8];
  assign N15264 = N14817 & N1415;
  assign N15265 = N14817 & idx_w_i[8];
  assign N15266 = N14819 & N1415;
  assign N15267 = N14819 & idx_w_i[8];
  assign N15268 = N14821 & N1415;
  assign N15269 = N14821 & idx_w_i[8];
  assign N15270 = N14823 & N1415;
  assign N15271 = N14823 & idx_w_i[8];
  assign N15272 = N14825 & N1415;
  assign N15273 = N14825 & idx_w_i[8];
  assign N15274 = N14827 & N1415;
  assign N15275 = N14827 & idx_w_i[8];
  assign N15276 = N14829 & N1415;
  assign N15277 = N14829 & idx_w_i[8];
  assign N15278 = N14831 & N1415;
  assign N15279 = N14831 & idx_w_i[8];
  assign N15280 = N14833 & N1415;
  assign N15281 = N14833 & idx_w_i[8];
  assign N15282 = N14835 & N1415;
  assign N15283 = N14835 & idx_w_i[8];
  assign N15284 = N14837 & N1415;
  assign N15285 = N14837 & idx_w_i[8];
  assign N15286 = N14839 & N1415;
  assign N15287 = N14839 & idx_w_i[8];
  assign N15288 = N14841 & N1415;
  assign N15289 = N14841 & idx_w_i[8];
  assign N15290 = N14843 & N1415;
  assign N15291 = N14843 & idx_w_i[8];
  assign N15292 = N14845 & N1415;
  assign N15293 = N14845 & idx_w_i[8];
  assign N15294 = N14847 & N1415;
  assign N15295 = N14847 & idx_w_i[8];
  assign N15296 = N14849 & N1415;
  assign N15297 = N14849 & idx_w_i[8];
  assign N15298 = N14851 & N1415;
  assign N15299 = N14851 & idx_w_i[8];
  assign N15300 = N14853 & N1415;
  assign N15301 = N14853 & idx_w_i[8];
  assign N15302 = N14855 & N1415;
  assign N15303 = N14855 & idx_w_i[8];
  assign N15304 = N14857 & N1415;
  assign N15305 = N14857 & idx_w_i[8];
  assign N15306 = N14859 & N1415;
  assign N15307 = N14859 & idx_w_i[8];
  assign N15308 = N14861 & N1415;
  assign N15309 = N14861 & idx_w_i[8];
  assign N15310 = N14863 & N1415;
  assign N15311 = N14863 & idx_w_i[8];
  assign N15312 = N14865 & N1415;
  assign N15313 = N14865 & idx_w_i[8];
  assign N15314 = N14867 & N1415;
  assign N15315 = N14867 & idx_w_i[8];
  assign N15316 = N14869 & N1415;
  assign N15317 = N14869 & idx_w_i[8];
  assign N15318 = N14871 & N1415;
  assign N15319 = N14871 & idx_w_i[8];
  assign N15320 = N14873 & N1415;
  assign N15321 = N14873 & idx_w_i[8];
  assign N15322 = N14875 & N1415;
  assign N15323 = N14875 & idx_w_i[8];
  assign N15324 = N14877 & N1415;
  assign N15325 = N14877 & idx_w_i[8];
  assign N15326 = N14879 & N1415;
  assign N15327 = N14879 & idx_w_i[8];
  assign N15328 = N14881 & N1415;
  assign N15329 = N14881 & idx_w_i[8];
  assign N15330 = N14883 & N1415;
  assign N15331 = N14883 & idx_w_i[8];
  assign N15332 = N14885 & N1415;
  assign N15333 = N14885 & idx_w_i[8];
  assign N15334 = N14887 & N1415;
  assign N15335 = N14887 & idx_w_i[8];
  assign N15336 = N14889 & N1415;
  assign N15337 = N14889 & idx_w_i[8];
  assign N15338 = N14891 & N1415;
  assign N15339 = N14891 & idx_w_i[8];
  assign N15340 = N14893 & N1415;
  assign N15341 = N14893 & idx_w_i[8];
  assign N15342 = N14895 & N1415;
  assign N15343 = N14895 & idx_w_i[8];
  assign N15344 = N14897 & N1415;
  assign N15345 = N14897 & idx_w_i[8];
  assign N15346 = N14899 & N1415;
  assign N15347 = N14899 & idx_w_i[8];
  assign N15348 = N14901 & N1415;
  assign N15349 = N14901 & idx_w_i[8];
  assign N15350 = N14903 & N1415;
  assign N15351 = N14903 & idx_w_i[8];
  assign N15352 = N14905 & N1415;
  assign N15353 = N14905 & idx_w_i[8];
  assign N15354 = N14907 & N1415;
  assign N15355 = N14907 & idx_w_i[8];
  assign N15356 = N14909 & N1415;
  assign N15357 = N14909 & idx_w_i[8];
  assign N15358 = N14911 & N1415;
  assign N15359 = N14911 & idx_w_i[8];
  assign N15360 = N14913 & N1415;
  assign N15361 = N14913 & idx_w_i[8];
  assign N15362 = N14915 & N1415;
  assign N15363 = N14915 & idx_w_i[8];
  assign N15364 = N14917 & N1415;
  assign N15365 = N14917 & idx_w_i[8];
  assign N15366 = N14919 & N1415;
  assign N15367 = N14919 & idx_w_i[8];
  assign N15368 = N14921 & N1415;
  assign N15369 = N14921 & idx_w_i[8];
  assign N15370 = N14923 & N1415;
  assign N15371 = N14923 & idx_w_i[8];
  assign N15372 = N14925 & N1415;
  assign N15373 = N14925 & idx_w_i[8];
  assign N15374 = N14927 & N1415;
  assign N15375 = N14927 & idx_w_i[8];
  assign N15376 = N14929 & N1415;
  assign N15377 = N14929 & idx_w_i[8];
  assign N15378 = N14931 & N1415;
  assign N15379 = N14931 & idx_w_i[8];
  assign N15380 = N14933 & N1415;
  assign N15381 = N14933 & idx_w_i[8];
  assign N15382 = N11473 & N1415;
  assign N15383 = N11475 & N1415;
  assign N15384 = N11477 & N1415;
  assign N15385 = N11479 & N1415;
  assign N15386 = N11481 & N1415;
  assign N15387 = N11483 & N1415;
  assign N15388 = N11485 & N1415;
  assign N15389 = N11487 & N1415;
  assign N15390 = N11489 & N1415;
  assign N15391 = N11491 & N1415;
  assign N15392 = N11493 & N1415;
  assign N15393 = N11495 & N1415;
  assign N15394 = N11497 & N1415;
  assign N15395 = N11499 & N1415;
  assign N15396 = N11501 & N1415;
  assign N15397 = N11503 & N1415;
  assign N15398 = N11505 & N1415;
  assign N15399 = N11507 & N1415;
  assign N15400 = N11509 & N1415;
  assign N15401 = N11511 & N1415;
  assign N15402 = N11513 & N1415;
  assign N15403 = N11515 & N1415;
  assign N15404 = N11517 & N1415;
  assign N15405 = N11519 & N1415;
  assign N15406 = N11521 & N1415;
  assign N15407 = N11523 & N1415;
  assign N15408 = N11525 & N1415;
  assign N15409 = N11527 & N1415;
  assign N15410 = N11529 & N1415;
  assign N15411 = N11531 & N1415;
  assign N15412 = N11533 & N1415;
  assign N15413 = N11535 & N1415;
  assign N15414 = N11537 & N1415;
  assign N15415 = N11539 & N1415;
  assign N15416 = N11541 & N1415;
  assign N15417 = N11543 & N1415;
  assign N15418 = N11545 & N1415;
  assign N15419 = N11547 & N1415;
  assign N15420 = N11549 & N1415;
  assign N15421 = N11551 & N1415;
  assign N15422 = N11553 & N1415;
  assign N15423 = N11555 & N1415;
  assign N15424 = N11557 & N1415;
  assign N15425 = N11559 & N1415;
  assign N15426 = N11561 & N1415;
  assign N15427 = N11563 & N1415;
  assign N15428 = N11565 & N1415;
  assign N15429 = N11567 & N1415;
  assign N15430 = N11569 & N1415;
  assign N15431 = N11571 & N1415;
  assign N15432 = N11573 & N1415;
  assign N15433 = N11575 & N1415;
  assign N15434 = N11577 & N1415;
  assign N15435 = N11579 & N1415;
  assign N15436 = N11581 & N1415;
  assign N15437 = N11583 & N1415;
  assign N15438 = N11585 & N1415;
  assign N15439 = N11587 & N1415;
  assign N15440 = N11589 & N1415;
  assign N15441 = N11591 & N1415;
  assign N15442 = N11593 & N1415;
  assign N15443 = N11595 & N1415;
  assign N15444 = N11597 & N1415;
  assign N15445 = N11599 & N1415;
  assign N15447 = ~N15446;
  assign N16496 = ~reset_i;
  assign N16497 = w_v_i & N16496;

endmodule