module bsg_mux_one_hot_width_p542_els_p2
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [1083:0] data_i;
  input [1:0] sel_one_hot_i;
  output [541:0] data_o;
  wire [541:0] data_o;
  wire [1083:0] data_masked;
  assign data_masked[541] = data_i[541] & sel_one_hot_i[0];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[0];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[0];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[0];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[0];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[0];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[0];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[0];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[0];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[0];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[0];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[0];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[0];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[0];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[0];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[0];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[0];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[0];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[0];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[0];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[0];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[0];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[0];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[0];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[0];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[0];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[0];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[0];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[0];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[0];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[0];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[0];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[0];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[0];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[0];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[0];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[0];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[0];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[0];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[0];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[0];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[0];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[0];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[0];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[0];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[0];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[0];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[0];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[0];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[0];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[0];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[0];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[0];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[0];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[0];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[0];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[0];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[0];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[0];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[0];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[0];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[0];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[0];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[0];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[0];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[0];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[0];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[0];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[0];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[0];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[0];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[0];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[0];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[0];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[0];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[0];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[0];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[0];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[0];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[0];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[0];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[0];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[0];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[0];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[0];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[0];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[0];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[0];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[0];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[0];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[0];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[0];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[0];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[0];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[0];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[0];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[0];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[0];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[0];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[0];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[0];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[0];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[0];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[0];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[0];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[0];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[0];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[0];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[0];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[0];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[0];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[0];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[0];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[0];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[0];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[0];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[0];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[0];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[0];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[0];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[0];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[0];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[0];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[0];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[0];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[0];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[0];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[0];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[0];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[0];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[0];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[0];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[0];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[0];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[0];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[0];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[0];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[0];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[0];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[0];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[0];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[0];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[0];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[0];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[0];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[0];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[0];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[0];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[0];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[0];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[0];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[0];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[0];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[0];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[0];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[0];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[0];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[0];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[0];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[0];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[0];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[0];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[0];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[0];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[0];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[0];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[0];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[0];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[0];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[0];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[0];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[0];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[0];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[0];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[0];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[0];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[0];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[0];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[0];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[0];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[0];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[0];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[0];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[0];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[0];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[0];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[0];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[0];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[0];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[0];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[0];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[0];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[0];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[0];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[0];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[0];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[0];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[0];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[0];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[0];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[0];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[0];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[0];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[0];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[0];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[0];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[0];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[0];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[0];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[0];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[0];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[0];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[0];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[0];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[0];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[0];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[0];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[0];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[0];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[0];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[0];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[0];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[0];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[0];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[0];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[0];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[0];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[0];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[0];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[0];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[0];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[0];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[0];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[0];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[0];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[0];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[0];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[0];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[0];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[0];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[0];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[0];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[0];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[0];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[0];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[0];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[0];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[0];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[0];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[0];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[0];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[0];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[0];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[0];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[0];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[0];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[0];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[0];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[0];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[0];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[0];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[0];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[0];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[0];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[0];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[0];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[0];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[0];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[0];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[0];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[0];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[0];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[0];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[0];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[0];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[0];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[0];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[0];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[0];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[0];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[0];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[0];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[0];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[0];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[0];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[0];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[0];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[0];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[0];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[0];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[0];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[0];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[0];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[0];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[0];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[0];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[0];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[0];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[0];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[0];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[0];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[0];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[0];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[0];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[0];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[0];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[0];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[0];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[0];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[0];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[0];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[0];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[0];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[0];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[0];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[0];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[0];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[0];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[0];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[0];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[0];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[0];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[0];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[0];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[0];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[0];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[0];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[0];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[0];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[0];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[0];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[0];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[0];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[0];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[0];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[0];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[0];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[0];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[0];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[0];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[0];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[0];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[0];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[0];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[0];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[0];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[0];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[0];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[0];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[0];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[0];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[0];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[0];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[0];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[0];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[0];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[0];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[0];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[0];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[0];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[0];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[0];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[0];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[0];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[0];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[0];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[0];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[0];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[0];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[0];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[0];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[0];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[0];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[0];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[0];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[0];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[0];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[0];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[0];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[0];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[0];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[0];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[0];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[0];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[0];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[0];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[0];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[0];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[0];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[0];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[0];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[0];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[0];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[0];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[0];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[0];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[0];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[0];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[0];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[0];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[0];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[0];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[0];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[0];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[0];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[0];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[0];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[0];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[0];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[0];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[0];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[0];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[0];
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[1083] = data_i[1083] & sel_one_hot_i[1];
  assign data_masked[1082] = data_i[1082] & sel_one_hot_i[1];
  assign data_masked[1081] = data_i[1081] & sel_one_hot_i[1];
  assign data_masked[1080] = data_i[1080] & sel_one_hot_i[1];
  assign data_masked[1079] = data_i[1079] & sel_one_hot_i[1];
  assign data_masked[1078] = data_i[1078] & sel_one_hot_i[1];
  assign data_masked[1077] = data_i[1077] & sel_one_hot_i[1];
  assign data_masked[1076] = data_i[1076] & sel_one_hot_i[1];
  assign data_masked[1075] = data_i[1075] & sel_one_hot_i[1];
  assign data_masked[1074] = data_i[1074] & sel_one_hot_i[1];
  assign data_masked[1073] = data_i[1073] & sel_one_hot_i[1];
  assign data_masked[1072] = data_i[1072] & sel_one_hot_i[1];
  assign data_masked[1071] = data_i[1071] & sel_one_hot_i[1];
  assign data_masked[1070] = data_i[1070] & sel_one_hot_i[1];
  assign data_masked[1069] = data_i[1069] & sel_one_hot_i[1];
  assign data_masked[1068] = data_i[1068] & sel_one_hot_i[1];
  assign data_masked[1067] = data_i[1067] & sel_one_hot_i[1];
  assign data_masked[1066] = data_i[1066] & sel_one_hot_i[1];
  assign data_masked[1065] = data_i[1065] & sel_one_hot_i[1];
  assign data_masked[1064] = data_i[1064] & sel_one_hot_i[1];
  assign data_masked[1063] = data_i[1063] & sel_one_hot_i[1];
  assign data_masked[1062] = data_i[1062] & sel_one_hot_i[1];
  assign data_masked[1061] = data_i[1061] & sel_one_hot_i[1];
  assign data_masked[1060] = data_i[1060] & sel_one_hot_i[1];
  assign data_masked[1059] = data_i[1059] & sel_one_hot_i[1];
  assign data_masked[1058] = data_i[1058] & sel_one_hot_i[1];
  assign data_masked[1057] = data_i[1057] & sel_one_hot_i[1];
  assign data_masked[1056] = data_i[1056] & sel_one_hot_i[1];
  assign data_masked[1055] = data_i[1055] & sel_one_hot_i[1];
  assign data_masked[1054] = data_i[1054] & sel_one_hot_i[1];
  assign data_masked[1053] = data_i[1053] & sel_one_hot_i[1];
  assign data_masked[1052] = data_i[1052] & sel_one_hot_i[1];
  assign data_masked[1051] = data_i[1051] & sel_one_hot_i[1];
  assign data_masked[1050] = data_i[1050] & sel_one_hot_i[1];
  assign data_masked[1049] = data_i[1049] & sel_one_hot_i[1];
  assign data_masked[1048] = data_i[1048] & sel_one_hot_i[1];
  assign data_masked[1047] = data_i[1047] & sel_one_hot_i[1];
  assign data_masked[1046] = data_i[1046] & sel_one_hot_i[1];
  assign data_masked[1045] = data_i[1045] & sel_one_hot_i[1];
  assign data_masked[1044] = data_i[1044] & sel_one_hot_i[1];
  assign data_masked[1043] = data_i[1043] & sel_one_hot_i[1];
  assign data_masked[1042] = data_i[1042] & sel_one_hot_i[1];
  assign data_masked[1041] = data_i[1041] & sel_one_hot_i[1];
  assign data_masked[1040] = data_i[1040] & sel_one_hot_i[1];
  assign data_masked[1039] = data_i[1039] & sel_one_hot_i[1];
  assign data_masked[1038] = data_i[1038] & sel_one_hot_i[1];
  assign data_masked[1037] = data_i[1037] & sel_one_hot_i[1];
  assign data_masked[1036] = data_i[1036] & sel_one_hot_i[1];
  assign data_masked[1035] = data_i[1035] & sel_one_hot_i[1];
  assign data_masked[1034] = data_i[1034] & sel_one_hot_i[1];
  assign data_masked[1033] = data_i[1033] & sel_one_hot_i[1];
  assign data_masked[1032] = data_i[1032] & sel_one_hot_i[1];
  assign data_masked[1031] = data_i[1031] & sel_one_hot_i[1];
  assign data_masked[1030] = data_i[1030] & sel_one_hot_i[1];
  assign data_masked[1029] = data_i[1029] & sel_one_hot_i[1];
  assign data_masked[1028] = data_i[1028] & sel_one_hot_i[1];
  assign data_masked[1027] = data_i[1027] & sel_one_hot_i[1];
  assign data_masked[1026] = data_i[1026] & sel_one_hot_i[1];
  assign data_masked[1025] = data_i[1025] & sel_one_hot_i[1];
  assign data_masked[1024] = data_i[1024] & sel_one_hot_i[1];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[1];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[1];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[1];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[1];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[1];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[1];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[1];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[1];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[1];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[1];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[1];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[1];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[1];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[1];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[1];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[1];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[1];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[1];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[1];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[1];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[1];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[1];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[1];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[1];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[1];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[1];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[1];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[1];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[1];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[1];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[1];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[1];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[1];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[1];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[1];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[1];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[1];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[1];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[1];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[1];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[1];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[1];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[1];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[1];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[1];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[1];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[1];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[1];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[1];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[1];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[1];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[1];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[1];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[1];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[1];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[1];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[1];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[1];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[1];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[1];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[1];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[1];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[1];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[1];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[1];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[1];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[1];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[1];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[1];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[1];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[1];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[1];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[1];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[1];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[1];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[1];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[1];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[1];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[1];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[1];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[1];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[1];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[1];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[1];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[1];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[1];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[1];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[1];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[1];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[1];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[1];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[1];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[1];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[1];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[1];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[1];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[1];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[1];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[1];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[1];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[1];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[1];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[1];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[1];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[1];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[1];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[1];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[1];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[1];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[1];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[1];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[1];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[1];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[1];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[1];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[1];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[1];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[1];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[1];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[1];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[1];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[1];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[1];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[1];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[1];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[1];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[1];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[1];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[1];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[1];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[1];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[1];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[1];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[1];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[1];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[1];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[1];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[1];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[1];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[1];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[1];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[1];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[1];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[1];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[1];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[1];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[1];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[1];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[1];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[1];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[1];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[1];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[1];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[1];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[1];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[1];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[1];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[1];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[1];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[1];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[1];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[1];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[1];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[1];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[1];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[1];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[1];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[1];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[1];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[1];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[1];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[1];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[1];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[1];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[1];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[1];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[1];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[1];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[1];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[1];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[1];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[1];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[1];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[1];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[1];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[1];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[1];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[1];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[1];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[1];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[1];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[1];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[1];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[1];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[1];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[1];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[1];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[1];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[1];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[1];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[1];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[1];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[1];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[1];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[1];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[1];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[1];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[1];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[1];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[1];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[1];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[1];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[1];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[1];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[1];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[1];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[1];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[1];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[1];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[1];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[1];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[1];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[1];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[1];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[1];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[1];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[1];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[1];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[1];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[1];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[1];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[1];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[1];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[1];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[1];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[1];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[1];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[1];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[1];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[1];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[1];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[1];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[1];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[1];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[1];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[1];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[1];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[1];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[1];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[1];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[1];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[1];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[1];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[1];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[1];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[1];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[1];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[1];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[1];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[1];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[1];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[1];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[1];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[1];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[1];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[1];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[1];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[1];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[1];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[1];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[1];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[1];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[1];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[1];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[1];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[1];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[1];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[1];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[1];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[1];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[1];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[1];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[1];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[1];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[1];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[1];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[1];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[1];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[1];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[1];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[1];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[1];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[1];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[1];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[1];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[1];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[1];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[1];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[1];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[1];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[1];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[1];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[1];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[1];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[1];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[1];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[1];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[1];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[1];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[1];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[1];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[1];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[1];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[1];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[1];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[1];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[1];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[1];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[1];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[1];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[1];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[1];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[1];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[1];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[1];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[1];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[1];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[1];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[1];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[1];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[1];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[1];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[1];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[1];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[1];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[1];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[1];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[1];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[1];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[1];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[1];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[1];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[1];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[1];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[1];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[1];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[1];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[1];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[1];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[1];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[1];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[1];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[1];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[1];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[1];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[1];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[1];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[1];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[1];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[1];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[1];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[1];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[1];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[1];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[1];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[1];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[1];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[1];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[1];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[1];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[1];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[1];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[1];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[1];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[1];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[1];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[1];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[1];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[1];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[1];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[1];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[1];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[1];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[1];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[1];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[1];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[1];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[1];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[1];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[1];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[1];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[1];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[1];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[1];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[1];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[1];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[1];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[1];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[1];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[1];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[1];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[1];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[1];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[1];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[1];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[1];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[1];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[1];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[1];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[1];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[1];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[1];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[1];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[1];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[1];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[1];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[1];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[1];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[1];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[1];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[1];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[1];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[1];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[1];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[1];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[1];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[1];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[1];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[1];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[1];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[1];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[1];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[1];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[1];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[1];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[1];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[1];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[1];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[1];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[1];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[1];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[1];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[1];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[1];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[1];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[1];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[1];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[1];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[1];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[1];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[1];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[1];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[1];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[1];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[1];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[1];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[1];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[1];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[1];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[1];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[1];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[1];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[1];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[1];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[1];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[1];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[1];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[1];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[1];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[1];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[1];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[1];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[1];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[1];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[1];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[1];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[1];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[1];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[1];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[1];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[1];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[1];
  assign data_o[0] = data_masked[542] | data_masked[0];
  assign data_o[1] = data_masked[543] | data_masked[1];
  assign data_o[2] = data_masked[544] | data_masked[2];
  assign data_o[3] = data_masked[545] | data_masked[3];
  assign data_o[4] = data_masked[546] | data_masked[4];
  assign data_o[5] = data_masked[547] | data_masked[5];
  assign data_o[6] = data_masked[548] | data_masked[6];
  assign data_o[7] = data_masked[549] | data_masked[7];
  assign data_o[8] = data_masked[550] | data_masked[8];
  assign data_o[9] = data_masked[551] | data_masked[9];
  assign data_o[10] = data_masked[552] | data_masked[10];
  assign data_o[11] = data_masked[553] | data_masked[11];
  assign data_o[12] = data_masked[554] | data_masked[12];
  assign data_o[13] = data_masked[555] | data_masked[13];
  assign data_o[14] = data_masked[556] | data_masked[14];
  assign data_o[15] = data_masked[557] | data_masked[15];
  assign data_o[16] = data_masked[558] | data_masked[16];
  assign data_o[17] = data_masked[559] | data_masked[17];
  assign data_o[18] = data_masked[560] | data_masked[18];
  assign data_o[19] = data_masked[561] | data_masked[19];
  assign data_o[20] = data_masked[562] | data_masked[20];
  assign data_o[21] = data_masked[563] | data_masked[21];
  assign data_o[22] = data_masked[564] | data_masked[22];
  assign data_o[23] = data_masked[565] | data_masked[23];
  assign data_o[24] = data_masked[566] | data_masked[24];
  assign data_o[25] = data_masked[567] | data_masked[25];
  assign data_o[26] = data_masked[568] | data_masked[26];
  assign data_o[27] = data_masked[569] | data_masked[27];
  assign data_o[28] = data_masked[570] | data_masked[28];
  assign data_o[29] = data_masked[571] | data_masked[29];
  assign data_o[30] = data_masked[572] | data_masked[30];
  assign data_o[31] = data_masked[573] | data_masked[31];
  assign data_o[32] = data_masked[574] | data_masked[32];
  assign data_o[33] = data_masked[575] | data_masked[33];
  assign data_o[34] = data_masked[576] | data_masked[34];
  assign data_o[35] = data_masked[577] | data_masked[35];
  assign data_o[36] = data_masked[578] | data_masked[36];
  assign data_o[37] = data_masked[579] | data_masked[37];
  assign data_o[38] = data_masked[580] | data_masked[38];
  assign data_o[39] = data_masked[581] | data_masked[39];
  assign data_o[40] = data_masked[582] | data_masked[40];
  assign data_o[41] = data_masked[583] | data_masked[41];
  assign data_o[42] = data_masked[584] | data_masked[42];
  assign data_o[43] = data_masked[585] | data_masked[43];
  assign data_o[44] = data_masked[586] | data_masked[44];
  assign data_o[45] = data_masked[587] | data_masked[45];
  assign data_o[46] = data_masked[588] | data_masked[46];
  assign data_o[47] = data_masked[589] | data_masked[47];
  assign data_o[48] = data_masked[590] | data_masked[48];
  assign data_o[49] = data_masked[591] | data_masked[49];
  assign data_o[50] = data_masked[592] | data_masked[50];
  assign data_o[51] = data_masked[593] | data_masked[51];
  assign data_o[52] = data_masked[594] | data_masked[52];
  assign data_o[53] = data_masked[595] | data_masked[53];
  assign data_o[54] = data_masked[596] | data_masked[54];
  assign data_o[55] = data_masked[597] | data_masked[55];
  assign data_o[56] = data_masked[598] | data_masked[56];
  assign data_o[57] = data_masked[599] | data_masked[57];
  assign data_o[58] = data_masked[600] | data_masked[58];
  assign data_o[59] = data_masked[601] | data_masked[59];
  assign data_o[60] = data_masked[602] | data_masked[60];
  assign data_o[61] = data_masked[603] | data_masked[61];
  assign data_o[62] = data_masked[604] | data_masked[62];
  assign data_o[63] = data_masked[605] | data_masked[63];
  assign data_o[64] = data_masked[606] | data_masked[64];
  assign data_o[65] = data_masked[607] | data_masked[65];
  assign data_o[66] = data_masked[608] | data_masked[66];
  assign data_o[67] = data_masked[609] | data_masked[67];
  assign data_o[68] = data_masked[610] | data_masked[68];
  assign data_o[69] = data_masked[611] | data_masked[69];
  assign data_o[70] = data_masked[612] | data_masked[70];
  assign data_o[71] = data_masked[613] | data_masked[71];
  assign data_o[72] = data_masked[614] | data_masked[72];
  assign data_o[73] = data_masked[615] | data_masked[73];
  assign data_o[74] = data_masked[616] | data_masked[74];
  assign data_o[75] = data_masked[617] | data_masked[75];
  assign data_o[76] = data_masked[618] | data_masked[76];
  assign data_o[77] = data_masked[619] | data_masked[77];
  assign data_o[78] = data_masked[620] | data_masked[78];
  assign data_o[79] = data_masked[621] | data_masked[79];
  assign data_o[80] = data_masked[622] | data_masked[80];
  assign data_o[81] = data_masked[623] | data_masked[81];
  assign data_o[82] = data_masked[624] | data_masked[82];
  assign data_o[83] = data_masked[625] | data_masked[83];
  assign data_o[84] = data_masked[626] | data_masked[84];
  assign data_o[85] = data_masked[627] | data_masked[85];
  assign data_o[86] = data_masked[628] | data_masked[86];
  assign data_o[87] = data_masked[629] | data_masked[87];
  assign data_o[88] = data_masked[630] | data_masked[88];
  assign data_o[89] = data_masked[631] | data_masked[89];
  assign data_o[90] = data_masked[632] | data_masked[90];
  assign data_o[91] = data_masked[633] | data_masked[91];
  assign data_o[92] = data_masked[634] | data_masked[92];
  assign data_o[93] = data_masked[635] | data_masked[93];
  assign data_o[94] = data_masked[636] | data_masked[94];
  assign data_o[95] = data_masked[637] | data_masked[95];
  assign data_o[96] = data_masked[638] | data_masked[96];
  assign data_o[97] = data_masked[639] | data_masked[97];
  assign data_o[98] = data_masked[640] | data_masked[98];
  assign data_o[99] = data_masked[641] | data_masked[99];
  assign data_o[100] = data_masked[642] | data_masked[100];
  assign data_o[101] = data_masked[643] | data_masked[101];
  assign data_o[102] = data_masked[644] | data_masked[102];
  assign data_o[103] = data_masked[645] | data_masked[103];
  assign data_o[104] = data_masked[646] | data_masked[104];
  assign data_o[105] = data_masked[647] | data_masked[105];
  assign data_o[106] = data_masked[648] | data_masked[106];
  assign data_o[107] = data_masked[649] | data_masked[107];
  assign data_o[108] = data_masked[650] | data_masked[108];
  assign data_o[109] = data_masked[651] | data_masked[109];
  assign data_o[110] = data_masked[652] | data_masked[110];
  assign data_o[111] = data_masked[653] | data_masked[111];
  assign data_o[112] = data_masked[654] | data_masked[112];
  assign data_o[113] = data_masked[655] | data_masked[113];
  assign data_o[114] = data_masked[656] | data_masked[114];
  assign data_o[115] = data_masked[657] | data_masked[115];
  assign data_o[116] = data_masked[658] | data_masked[116];
  assign data_o[117] = data_masked[659] | data_masked[117];
  assign data_o[118] = data_masked[660] | data_masked[118];
  assign data_o[119] = data_masked[661] | data_masked[119];
  assign data_o[120] = data_masked[662] | data_masked[120];
  assign data_o[121] = data_masked[663] | data_masked[121];
  assign data_o[122] = data_masked[664] | data_masked[122];
  assign data_o[123] = data_masked[665] | data_masked[123];
  assign data_o[124] = data_masked[666] | data_masked[124];
  assign data_o[125] = data_masked[667] | data_masked[125];
  assign data_o[126] = data_masked[668] | data_masked[126];
  assign data_o[127] = data_masked[669] | data_masked[127];
  assign data_o[128] = data_masked[670] | data_masked[128];
  assign data_o[129] = data_masked[671] | data_masked[129];
  assign data_o[130] = data_masked[672] | data_masked[130];
  assign data_o[131] = data_masked[673] | data_masked[131];
  assign data_o[132] = data_masked[674] | data_masked[132];
  assign data_o[133] = data_masked[675] | data_masked[133];
  assign data_o[134] = data_masked[676] | data_masked[134];
  assign data_o[135] = data_masked[677] | data_masked[135];
  assign data_o[136] = data_masked[678] | data_masked[136];
  assign data_o[137] = data_masked[679] | data_masked[137];
  assign data_o[138] = data_masked[680] | data_masked[138];
  assign data_o[139] = data_masked[681] | data_masked[139];
  assign data_o[140] = data_masked[682] | data_masked[140];
  assign data_o[141] = data_masked[683] | data_masked[141];
  assign data_o[142] = data_masked[684] | data_masked[142];
  assign data_o[143] = data_masked[685] | data_masked[143];
  assign data_o[144] = data_masked[686] | data_masked[144];
  assign data_o[145] = data_masked[687] | data_masked[145];
  assign data_o[146] = data_masked[688] | data_masked[146];
  assign data_o[147] = data_masked[689] | data_masked[147];
  assign data_o[148] = data_masked[690] | data_masked[148];
  assign data_o[149] = data_masked[691] | data_masked[149];
  assign data_o[150] = data_masked[692] | data_masked[150];
  assign data_o[151] = data_masked[693] | data_masked[151];
  assign data_o[152] = data_masked[694] | data_masked[152];
  assign data_o[153] = data_masked[695] | data_masked[153];
  assign data_o[154] = data_masked[696] | data_masked[154];
  assign data_o[155] = data_masked[697] | data_masked[155];
  assign data_o[156] = data_masked[698] | data_masked[156];
  assign data_o[157] = data_masked[699] | data_masked[157];
  assign data_o[158] = data_masked[700] | data_masked[158];
  assign data_o[159] = data_masked[701] | data_masked[159];
  assign data_o[160] = data_masked[702] | data_masked[160];
  assign data_o[161] = data_masked[703] | data_masked[161];
  assign data_o[162] = data_masked[704] | data_masked[162];
  assign data_o[163] = data_masked[705] | data_masked[163];
  assign data_o[164] = data_masked[706] | data_masked[164];
  assign data_o[165] = data_masked[707] | data_masked[165];
  assign data_o[166] = data_masked[708] | data_masked[166];
  assign data_o[167] = data_masked[709] | data_masked[167];
  assign data_o[168] = data_masked[710] | data_masked[168];
  assign data_o[169] = data_masked[711] | data_masked[169];
  assign data_o[170] = data_masked[712] | data_masked[170];
  assign data_o[171] = data_masked[713] | data_masked[171];
  assign data_o[172] = data_masked[714] | data_masked[172];
  assign data_o[173] = data_masked[715] | data_masked[173];
  assign data_o[174] = data_masked[716] | data_masked[174];
  assign data_o[175] = data_masked[717] | data_masked[175];
  assign data_o[176] = data_masked[718] | data_masked[176];
  assign data_o[177] = data_masked[719] | data_masked[177];
  assign data_o[178] = data_masked[720] | data_masked[178];
  assign data_o[179] = data_masked[721] | data_masked[179];
  assign data_o[180] = data_masked[722] | data_masked[180];
  assign data_o[181] = data_masked[723] | data_masked[181];
  assign data_o[182] = data_masked[724] | data_masked[182];
  assign data_o[183] = data_masked[725] | data_masked[183];
  assign data_o[184] = data_masked[726] | data_masked[184];
  assign data_o[185] = data_masked[727] | data_masked[185];
  assign data_o[186] = data_masked[728] | data_masked[186];
  assign data_o[187] = data_masked[729] | data_masked[187];
  assign data_o[188] = data_masked[730] | data_masked[188];
  assign data_o[189] = data_masked[731] | data_masked[189];
  assign data_o[190] = data_masked[732] | data_masked[190];
  assign data_o[191] = data_masked[733] | data_masked[191];
  assign data_o[192] = data_masked[734] | data_masked[192];
  assign data_o[193] = data_masked[735] | data_masked[193];
  assign data_o[194] = data_masked[736] | data_masked[194];
  assign data_o[195] = data_masked[737] | data_masked[195];
  assign data_o[196] = data_masked[738] | data_masked[196];
  assign data_o[197] = data_masked[739] | data_masked[197];
  assign data_o[198] = data_masked[740] | data_masked[198];
  assign data_o[199] = data_masked[741] | data_masked[199];
  assign data_o[200] = data_masked[742] | data_masked[200];
  assign data_o[201] = data_masked[743] | data_masked[201];
  assign data_o[202] = data_masked[744] | data_masked[202];
  assign data_o[203] = data_masked[745] | data_masked[203];
  assign data_o[204] = data_masked[746] | data_masked[204];
  assign data_o[205] = data_masked[747] | data_masked[205];
  assign data_o[206] = data_masked[748] | data_masked[206];
  assign data_o[207] = data_masked[749] | data_masked[207];
  assign data_o[208] = data_masked[750] | data_masked[208];
  assign data_o[209] = data_masked[751] | data_masked[209];
  assign data_o[210] = data_masked[752] | data_masked[210];
  assign data_o[211] = data_masked[753] | data_masked[211];
  assign data_o[212] = data_masked[754] | data_masked[212];
  assign data_o[213] = data_masked[755] | data_masked[213];
  assign data_o[214] = data_masked[756] | data_masked[214];
  assign data_o[215] = data_masked[757] | data_masked[215];
  assign data_o[216] = data_masked[758] | data_masked[216];
  assign data_o[217] = data_masked[759] | data_masked[217];
  assign data_o[218] = data_masked[760] | data_masked[218];
  assign data_o[219] = data_masked[761] | data_masked[219];
  assign data_o[220] = data_masked[762] | data_masked[220];
  assign data_o[221] = data_masked[763] | data_masked[221];
  assign data_o[222] = data_masked[764] | data_masked[222];
  assign data_o[223] = data_masked[765] | data_masked[223];
  assign data_o[224] = data_masked[766] | data_masked[224];
  assign data_o[225] = data_masked[767] | data_masked[225];
  assign data_o[226] = data_masked[768] | data_masked[226];
  assign data_o[227] = data_masked[769] | data_masked[227];
  assign data_o[228] = data_masked[770] | data_masked[228];
  assign data_o[229] = data_masked[771] | data_masked[229];
  assign data_o[230] = data_masked[772] | data_masked[230];
  assign data_o[231] = data_masked[773] | data_masked[231];
  assign data_o[232] = data_masked[774] | data_masked[232];
  assign data_o[233] = data_masked[775] | data_masked[233];
  assign data_o[234] = data_masked[776] | data_masked[234];
  assign data_o[235] = data_masked[777] | data_masked[235];
  assign data_o[236] = data_masked[778] | data_masked[236];
  assign data_o[237] = data_masked[779] | data_masked[237];
  assign data_o[238] = data_masked[780] | data_masked[238];
  assign data_o[239] = data_masked[781] | data_masked[239];
  assign data_o[240] = data_masked[782] | data_masked[240];
  assign data_o[241] = data_masked[783] | data_masked[241];
  assign data_o[242] = data_masked[784] | data_masked[242];
  assign data_o[243] = data_masked[785] | data_masked[243];
  assign data_o[244] = data_masked[786] | data_masked[244];
  assign data_o[245] = data_masked[787] | data_masked[245];
  assign data_o[246] = data_masked[788] | data_masked[246];
  assign data_o[247] = data_masked[789] | data_masked[247];
  assign data_o[248] = data_masked[790] | data_masked[248];
  assign data_o[249] = data_masked[791] | data_masked[249];
  assign data_o[250] = data_masked[792] | data_masked[250];
  assign data_o[251] = data_masked[793] | data_masked[251];
  assign data_o[252] = data_masked[794] | data_masked[252];
  assign data_o[253] = data_masked[795] | data_masked[253];
  assign data_o[254] = data_masked[796] | data_masked[254];
  assign data_o[255] = data_masked[797] | data_masked[255];
  assign data_o[256] = data_masked[798] | data_masked[256];
  assign data_o[257] = data_masked[799] | data_masked[257];
  assign data_o[258] = data_masked[800] | data_masked[258];
  assign data_o[259] = data_masked[801] | data_masked[259];
  assign data_o[260] = data_masked[802] | data_masked[260];
  assign data_o[261] = data_masked[803] | data_masked[261];
  assign data_o[262] = data_masked[804] | data_masked[262];
  assign data_o[263] = data_masked[805] | data_masked[263];
  assign data_o[264] = data_masked[806] | data_masked[264];
  assign data_o[265] = data_masked[807] | data_masked[265];
  assign data_o[266] = data_masked[808] | data_masked[266];
  assign data_o[267] = data_masked[809] | data_masked[267];
  assign data_o[268] = data_masked[810] | data_masked[268];
  assign data_o[269] = data_masked[811] | data_masked[269];
  assign data_o[270] = data_masked[812] | data_masked[270];
  assign data_o[271] = data_masked[813] | data_masked[271];
  assign data_o[272] = data_masked[814] | data_masked[272];
  assign data_o[273] = data_masked[815] | data_masked[273];
  assign data_o[274] = data_masked[816] | data_masked[274];
  assign data_o[275] = data_masked[817] | data_masked[275];
  assign data_o[276] = data_masked[818] | data_masked[276];
  assign data_o[277] = data_masked[819] | data_masked[277];
  assign data_o[278] = data_masked[820] | data_masked[278];
  assign data_o[279] = data_masked[821] | data_masked[279];
  assign data_o[280] = data_masked[822] | data_masked[280];
  assign data_o[281] = data_masked[823] | data_masked[281];
  assign data_o[282] = data_masked[824] | data_masked[282];
  assign data_o[283] = data_masked[825] | data_masked[283];
  assign data_o[284] = data_masked[826] | data_masked[284];
  assign data_o[285] = data_masked[827] | data_masked[285];
  assign data_o[286] = data_masked[828] | data_masked[286];
  assign data_o[287] = data_masked[829] | data_masked[287];
  assign data_o[288] = data_masked[830] | data_masked[288];
  assign data_o[289] = data_masked[831] | data_masked[289];
  assign data_o[290] = data_masked[832] | data_masked[290];
  assign data_o[291] = data_masked[833] | data_masked[291];
  assign data_o[292] = data_masked[834] | data_masked[292];
  assign data_o[293] = data_masked[835] | data_masked[293];
  assign data_o[294] = data_masked[836] | data_masked[294];
  assign data_o[295] = data_masked[837] | data_masked[295];
  assign data_o[296] = data_masked[838] | data_masked[296];
  assign data_o[297] = data_masked[839] | data_masked[297];
  assign data_o[298] = data_masked[840] | data_masked[298];
  assign data_o[299] = data_masked[841] | data_masked[299];
  assign data_o[300] = data_masked[842] | data_masked[300];
  assign data_o[301] = data_masked[843] | data_masked[301];
  assign data_o[302] = data_masked[844] | data_masked[302];
  assign data_o[303] = data_masked[845] | data_masked[303];
  assign data_o[304] = data_masked[846] | data_masked[304];
  assign data_o[305] = data_masked[847] | data_masked[305];
  assign data_o[306] = data_masked[848] | data_masked[306];
  assign data_o[307] = data_masked[849] | data_masked[307];
  assign data_o[308] = data_masked[850] | data_masked[308];
  assign data_o[309] = data_masked[851] | data_masked[309];
  assign data_o[310] = data_masked[852] | data_masked[310];
  assign data_o[311] = data_masked[853] | data_masked[311];
  assign data_o[312] = data_masked[854] | data_masked[312];
  assign data_o[313] = data_masked[855] | data_masked[313];
  assign data_o[314] = data_masked[856] | data_masked[314];
  assign data_o[315] = data_masked[857] | data_masked[315];
  assign data_o[316] = data_masked[858] | data_masked[316];
  assign data_o[317] = data_masked[859] | data_masked[317];
  assign data_o[318] = data_masked[860] | data_masked[318];
  assign data_o[319] = data_masked[861] | data_masked[319];
  assign data_o[320] = data_masked[862] | data_masked[320];
  assign data_o[321] = data_masked[863] | data_masked[321];
  assign data_o[322] = data_masked[864] | data_masked[322];
  assign data_o[323] = data_masked[865] | data_masked[323];
  assign data_o[324] = data_masked[866] | data_masked[324];
  assign data_o[325] = data_masked[867] | data_masked[325];
  assign data_o[326] = data_masked[868] | data_masked[326];
  assign data_o[327] = data_masked[869] | data_masked[327];
  assign data_o[328] = data_masked[870] | data_masked[328];
  assign data_o[329] = data_masked[871] | data_masked[329];
  assign data_o[330] = data_masked[872] | data_masked[330];
  assign data_o[331] = data_masked[873] | data_masked[331];
  assign data_o[332] = data_masked[874] | data_masked[332];
  assign data_o[333] = data_masked[875] | data_masked[333];
  assign data_o[334] = data_masked[876] | data_masked[334];
  assign data_o[335] = data_masked[877] | data_masked[335];
  assign data_o[336] = data_masked[878] | data_masked[336];
  assign data_o[337] = data_masked[879] | data_masked[337];
  assign data_o[338] = data_masked[880] | data_masked[338];
  assign data_o[339] = data_masked[881] | data_masked[339];
  assign data_o[340] = data_masked[882] | data_masked[340];
  assign data_o[341] = data_masked[883] | data_masked[341];
  assign data_o[342] = data_masked[884] | data_masked[342];
  assign data_o[343] = data_masked[885] | data_masked[343];
  assign data_o[344] = data_masked[886] | data_masked[344];
  assign data_o[345] = data_masked[887] | data_masked[345];
  assign data_o[346] = data_masked[888] | data_masked[346];
  assign data_o[347] = data_masked[889] | data_masked[347];
  assign data_o[348] = data_masked[890] | data_masked[348];
  assign data_o[349] = data_masked[891] | data_masked[349];
  assign data_o[350] = data_masked[892] | data_masked[350];
  assign data_o[351] = data_masked[893] | data_masked[351];
  assign data_o[352] = data_masked[894] | data_masked[352];
  assign data_o[353] = data_masked[895] | data_masked[353];
  assign data_o[354] = data_masked[896] | data_masked[354];
  assign data_o[355] = data_masked[897] | data_masked[355];
  assign data_o[356] = data_masked[898] | data_masked[356];
  assign data_o[357] = data_masked[899] | data_masked[357];
  assign data_o[358] = data_masked[900] | data_masked[358];
  assign data_o[359] = data_masked[901] | data_masked[359];
  assign data_o[360] = data_masked[902] | data_masked[360];
  assign data_o[361] = data_masked[903] | data_masked[361];
  assign data_o[362] = data_masked[904] | data_masked[362];
  assign data_o[363] = data_masked[905] | data_masked[363];
  assign data_o[364] = data_masked[906] | data_masked[364];
  assign data_o[365] = data_masked[907] | data_masked[365];
  assign data_o[366] = data_masked[908] | data_masked[366];
  assign data_o[367] = data_masked[909] | data_masked[367];
  assign data_o[368] = data_masked[910] | data_masked[368];
  assign data_o[369] = data_masked[911] | data_masked[369];
  assign data_o[370] = data_masked[912] | data_masked[370];
  assign data_o[371] = data_masked[913] | data_masked[371];
  assign data_o[372] = data_masked[914] | data_masked[372];
  assign data_o[373] = data_masked[915] | data_masked[373];
  assign data_o[374] = data_masked[916] | data_masked[374];
  assign data_o[375] = data_masked[917] | data_masked[375];
  assign data_o[376] = data_masked[918] | data_masked[376];
  assign data_o[377] = data_masked[919] | data_masked[377];
  assign data_o[378] = data_masked[920] | data_masked[378];
  assign data_o[379] = data_masked[921] | data_masked[379];
  assign data_o[380] = data_masked[922] | data_masked[380];
  assign data_o[381] = data_masked[923] | data_masked[381];
  assign data_o[382] = data_masked[924] | data_masked[382];
  assign data_o[383] = data_masked[925] | data_masked[383];
  assign data_o[384] = data_masked[926] | data_masked[384];
  assign data_o[385] = data_masked[927] | data_masked[385];
  assign data_o[386] = data_masked[928] | data_masked[386];
  assign data_o[387] = data_masked[929] | data_masked[387];
  assign data_o[388] = data_masked[930] | data_masked[388];
  assign data_o[389] = data_masked[931] | data_masked[389];
  assign data_o[390] = data_masked[932] | data_masked[390];
  assign data_o[391] = data_masked[933] | data_masked[391];
  assign data_o[392] = data_masked[934] | data_masked[392];
  assign data_o[393] = data_masked[935] | data_masked[393];
  assign data_o[394] = data_masked[936] | data_masked[394];
  assign data_o[395] = data_masked[937] | data_masked[395];
  assign data_o[396] = data_masked[938] | data_masked[396];
  assign data_o[397] = data_masked[939] | data_masked[397];
  assign data_o[398] = data_masked[940] | data_masked[398];
  assign data_o[399] = data_masked[941] | data_masked[399];
  assign data_o[400] = data_masked[942] | data_masked[400];
  assign data_o[401] = data_masked[943] | data_masked[401];
  assign data_o[402] = data_masked[944] | data_masked[402];
  assign data_o[403] = data_masked[945] | data_masked[403];
  assign data_o[404] = data_masked[946] | data_masked[404];
  assign data_o[405] = data_masked[947] | data_masked[405];
  assign data_o[406] = data_masked[948] | data_masked[406];
  assign data_o[407] = data_masked[949] | data_masked[407];
  assign data_o[408] = data_masked[950] | data_masked[408];
  assign data_o[409] = data_masked[951] | data_masked[409];
  assign data_o[410] = data_masked[952] | data_masked[410];
  assign data_o[411] = data_masked[953] | data_masked[411];
  assign data_o[412] = data_masked[954] | data_masked[412];
  assign data_o[413] = data_masked[955] | data_masked[413];
  assign data_o[414] = data_masked[956] | data_masked[414];
  assign data_o[415] = data_masked[957] | data_masked[415];
  assign data_o[416] = data_masked[958] | data_masked[416];
  assign data_o[417] = data_masked[959] | data_masked[417];
  assign data_o[418] = data_masked[960] | data_masked[418];
  assign data_o[419] = data_masked[961] | data_masked[419];
  assign data_o[420] = data_masked[962] | data_masked[420];
  assign data_o[421] = data_masked[963] | data_masked[421];
  assign data_o[422] = data_masked[964] | data_masked[422];
  assign data_o[423] = data_masked[965] | data_masked[423];
  assign data_o[424] = data_masked[966] | data_masked[424];
  assign data_o[425] = data_masked[967] | data_masked[425];
  assign data_o[426] = data_masked[968] | data_masked[426];
  assign data_o[427] = data_masked[969] | data_masked[427];
  assign data_o[428] = data_masked[970] | data_masked[428];
  assign data_o[429] = data_masked[971] | data_masked[429];
  assign data_o[430] = data_masked[972] | data_masked[430];
  assign data_o[431] = data_masked[973] | data_masked[431];
  assign data_o[432] = data_masked[974] | data_masked[432];
  assign data_o[433] = data_masked[975] | data_masked[433];
  assign data_o[434] = data_masked[976] | data_masked[434];
  assign data_o[435] = data_masked[977] | data_masked[435];
  assign data_o[436] = data_masked[978] | data_masked[436];
  assign data_o[437] = data_masked[979] | data_masked[437];
  assign data_o[438] = data_masked[980] | data_masked[438];
  assign data_o[439] = data_masked[981] | data_masked[439];
  assign data_o[440] = data_masked[982] | data_masked[440];
  assign data_o[441] = data_masked[983] | data_masked[441];
  assign data_o[442] = data_masked[984] | data_masked[442];
  assign data_o[443] = data_masked[985] | data_masked[443];
  assign data_o[444] = data_masked[986] | data_masked[444];
  assign data_o[445] = data_masked[987] | data_masked[445];
  assign data_o[446] = data_masked[988] | data_masked[446];
  assign data_o[447] = data_masked[989] | data_masked[447];
  assign data_o[448] = data_masked[990] | data_masked[448];
  assign data_o[449] = data_masked[991] | data_masked[449];
  assign data_o[450] = data_masked[992] | data_masked[450];
  assign data_o[451] = data_masked[993] | data_masked[451];
  assign data_o[452] = data_masked[994] | data_masked[452];
  assign data_o[453] = data_masked[995] | data_masked[453];
  assign data_o[454] = data_masked[996] | data_masked[454];
  assign data_o[455] = data_masked[997] | data_masked[455];
  assign data_o[456] = data_masked[998] | data_masked[456];
  assign data_o[457] = data_masked[999] | data_masked[457];
  assign data_o[458] = data_masked[1000] | data_masked[458];
  assign data_o[459] = data_masked[1001] | data_masked[459];
  assign data_o[460] = data_masked[1002] | data_masked[460];
  assign data_o[461] = data_masked[1003] | data_masked[461];
  assign data_o[462] = data_masked[1004] | data_masked[462];
  assign data_o[463] = data_masked[1005] | data_masked[463];
  assign data_o[464] = data_masked[1006] | data_masked[464];
  assign data_o[465] = data_masked[1007] | data_masked[465];
  assign data_o[466] = data_masked[1008] | data_masked[466];
  assign data_o[467] = data_masked[1009] | data_masked[467];
  assign data_o[468] = data_masked[1010] | data_masked[468];
  assign data_o[469] = data_masked[1011] | data_masked[469];
  assign data_o[470] = data_masked[1012] | data_masked[470];
  assign data_o[471] = data_masked[1013] | data_masked[471];
  assign data_o[472] = data_masked[1014] | data_masked[472];
  assign data_o[473] = data_masked[1015] | data_masked[473];
  assign data_o[474] = data_masked[1016] | data_masked[474];
  assign data_o[475] = data_masked[1017] | data_masked[475];
  assign data_o[476] = data_masked[1018] | data_masked[476];
  assign data_o[477] = data_masked[1019] | data_masked[477];
  assign data_o[478] = data_masked[1020] | data_masked[478];
  assign data_o[479] = data_masked[1021] | data_masked[479];
  assign data_o[480] = data_masked[1022] | data_masked[480];
  assign data_o[481] = data_masked[1023] | data_masked[481];
  assign data_o[482] = data_masked[1024] | data_masked[482];
  assign data_o[483] = data_masked[1025] | data_masked[483];
  assign data_o[484] = data_masked[1026] | data_masked[484];
  assign data_o[485] = data_masked[1027] | data_masked[485];
  assign data_o[486] = data_masked[1028] | data_masked[486];
  assign data_o[487] = data_masked[1029] | data_masked[487];
  assign data_o[488] = data_masked[1030] | data_masked[488];
  assign data_o[489] = data_masked[1031] | data_masked[489];
  assign data_o[490] = data_masked[1032] | data_masked[490];
  assign data_o[491] = data_masked[1033] | data_masked[491];
  assign data_o[492] = data_masked[1034] | data_masked[492];
  assign data_o[493] = data_masked[1035] | data_masked[493];
  assign data_o[494] = data_masked[1036] | data_masked[494];
  assign data_o[495] = data_masked[1037] | data_masked[495];
  assign data_o[496] = data_masked[1038] | data_masked[496];
  assign data_o[497] = data_masked[1039] | data_masked[497];
  assign data_o[498] = data_masked[1040] | data_masked[498];
  assign data_o[499] = data_masked[1041] | data_masked[499];
  assign data_o[500] = data_masked[1042] | data_masked[500];
  assign data_o[501] = data_masked[1043] | data_masked[501];
  assign data_o[502] = data_masked[1044] | data_masked[502];
  assign data_o[503] = data_masked[1045] | data_masked[503];
  assign data_o[504] = data_masked[1046] | data_masked[504];
  assign data_o[505] = data_masked[1047] | data_masked[505];
  assign data_o[506] = data_masked[1048] | data_masked[506];
  assign data_o[507] = data_masked[1049] | data_masked[507];
  assign data_o[508] = data_masked[1050] | data_masked[508];
  assign data_o[509] = data_masked[1051] | data_masked[509];
  assign data_o[510] = data_masked[1052] | data_masked[510];
  assign data_o[511] = data_masked[1053] | data_masked[511];
  assign data_o[512] = data_masked[1054] | data_masked[512];
  assign data_o[513] = data_masked[1055] | data_masked[513];
  assign data_o[514] = data_masked[1056] | data_masked[514];
  assign data_o[515] = data_masked[1057] | data_masked[515];
  assign data_o[516] = data_masked[1058] | data_masked[516];
  assign data_o[517] = data_masked[1059] | data_masked[517];
  assign data_o[518] = data_masked[1060] | data_masked[518];
  assign data_o[519] = data_masked[1061] | data_masked[519];
  assign data_o[520] = data_masked[1062] | data_masked[520];
  assign data_o[521] = data_masked[1063] | data_masked[521];
  assign data_o[522] = data_masked[1064] | data_masked[522];
  assign data_o[523] = data_masked[1065] | data_masked[523];
  assign data_o[524] = data_masked[1066] | data_masked[524];
  assign data_o[525] = data_masked[1067] | data_masked[525];
  assign data_o[526] = data_masked[1068] | data_masked[526];
  assign data_o[527] = data_masked[1069] | data_masked[527];
  assign data_o[528] = data_masked[1070] | data_masked[528];
  assign data_o[529] = data_masked[1071] | data_masked[529];
  assign data_o[530] = data_masked[1072] | data_masked[530];
  assign data_o[531] = data_masked[1073] | data_masked[531];
  assign data_o[532] = data_masked[1074] | data_masked[532];
  assign data_o[533] = data_masked[1075] | data_masked[533];
  assign data_o[534] = data_masked[1076] | data_masked[534];
  assign data_o[535] = data_masked[1077] | data_masked[535];
  assign data_o[536] = data_masked[1078] | data_masked[536];
  assign data_o[537] = data_masked[1079] | data_masked[537];
  assign data_o[538] = data_masked[1080] | data_masked[538];
  assign data_o[539] = data_masked[1081] | data_masked[539];
  assign data_o[540] = data_masked[1082] | data_masked[540];
  assign data_o[541] = data_masked[1083] | data_masked[541];

endmodule