module DCacheModuleanon3( // @[:freechips.rocketchip.system.TinyConfig.fir@103149.2]
  input         io_in_0_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [7:0]  io_in_0_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input         io_in_0_bits_write, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [31:0] io_in_0_bits_wdata, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [3:0]  io_in_0_bits_eccMask, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output        io_in_1_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input         io_in_1_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [7:0]  io_in_1_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input         io_in_1_bits_write, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [31:0] io_in_1_bits_wdata, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [3:0]  io_in_1_bits_eccMask, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output        io_in_3_ready, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input         io_in_3_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [7:0]  io_in_3_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [31:0] io_in_3_bits_wdata, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  input  [3:0]  io_in_3_bits_eccMask, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output        io_out_valid, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output [7:0]  io_out_bits_addr, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output        io_out_bits_write, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output [31:0] io_out_bits_wdata, // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
  output [3:0]  io_out_bits_eccMask // @[:freechips.rocketchip.system.TinyConfig.fir@103152.4]
);
  wire [3:0] _GEN_9; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  wire [31:0] _GEN_11; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  wire  _GEN_12; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  wire [7:0] _GEN_13; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  wire  _T; // @[Arbiter.scala 31:68:freechips.rocketchip.system.TinyConfig.fir@103188.4]
  wire  _T_3; // @[Arbiter.scala 31:78:freechips.rocketchip.system.TinyConfig.fir@103191.4]
  wire  _T_9; // @[Arbiter.scala 135:19:freechips.rocketchip.system.TinyConfig.fir@103201.4]
  assign _GEN_9 = io_in_1_valid ? io_in_1_bits_eccMask : io_in_3_bits_eccMask; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  assign _GEN_11 = io_in_1_valid ? io_in_1_bits_wdata : io_in_3_bits_wdata; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  assign _GEN_12 = io_in_1_valid ? io_in_1_bits_write : 1'h0; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  assign _GEN_13 = io_in_1_valid ? io_in_1_bits_addr : io_in_3_bits_addr; // @[Arbiter.scala 126:27:freechips.rocketchip.system.TinyConfig.fir@103170.4]
  assign _T = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68:freechips.rocketchip.system.TinyConfig.fir@103188.4]
  assign _T_3 = _T == 1'h0; // @[Arbiter.scala 31:78:freechips.rocketchip.system.TinyConfig.fir@103191.4]
  assign _T_9 = _T_3 == 1'h0; // @[Arbiter.scala 135:19:freechips.rocketchip.system.TinyConfig.fir@103201.4]
  assign io_in_1_ready = io_in_0_valid == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.TinyConfig.fir@103196.4]
  assign io_in_3_ready = _T == 1'h0; // @[Arbiter.scala 134:14:freechips.rocketchip.system.TinyConfig.fir@103200.4]
  assign io_out_valid = _T_9 | io_in_3_valid; // @[Arbiter.scala 135:16:freechips.rocketchip.system.TinyConfig.fir@103203.4]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : _GEN_13; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@103160.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103168.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103177.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103186.6]
  assign io_out_bits_write = io_in_0_valid ? io_in_0_bits_write : _GEN_12; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@103159.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103167.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103176.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103185.6]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : _GEN_11; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@103158.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103166.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103175.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103184.6]
  assign io_out_bits_eccMask = io_in_0_valid ? io_in_0_bits_eccMask : _GEN_9; // @[Arbiter.scala 124:15:freechips.rocketchip.system.TinyConfig.fir@103156.4 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103164.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103173.6 Arbiter.scala 128:19:freechips.rocketchip.system.TinyConfig.fir@103182.6]
endmodule