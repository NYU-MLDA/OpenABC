module core_debug_0(clk, rst, dmi_addr, dmi_din, dmi_req, dmi_wr, terminate, core_stopped, nia, msr, dbg_gpr_ack, dbg_gpr_data, log_data, log_read_addr, dmi_dout, dmi_ack, core_stop, core_rst, icache_rst, dbg_gpr_req, dbg_gpr_addr, log_read_data, log_write_addr, terminated_out);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  wire _06_;
  wire _07_;
  wire _08_;
  wire _09_;
  wire _10_;
  wire [63:0] _11_;
  wire _12_;
  wire _13_;
  wire _14_;
  wire [31:0] _15_;
  wire _16_;
  wire [7:0] _17_;
  wire _18_;
  wire [7:0] _19_;
  wire _20_;
  wire _21_;
  wire _22_;
  wire _23_;
  wire _24_;
  wire _25_;
  wire _26_;
  wire _27_;
  wire _28_;
  wire _29_;
  wire _30_;
  wire _31_;
  wire _32_;
  wire _33_;
  wire [63:0] _34_;
  wire [31:0] _35_;
  wire [63:0] _36_;
  wire [6:0] _37_;
  wire [31:0] _38_;
  wire [63:0] _39_;
  wire _40_;
  wire _41_;
  wire _42_;
  wire _43_;
  wire _44_;
  wire [6:0] _45_;
  wire [31:0] _46_;
  wire [63:0] _47_;
  wire _48_;
  wire _49_;
  wire _50_;
  wire _51_;
  wire _52_;
  wire [6:0] _53_;
  wire [31:0] _54_;
  wire [63:0] _55_;
  wire _56_;
  wire _57_;
  wire [1:0] _58_;
  wire [1:0] _59_;
  wire _60_;
  wire _61_;
  wire _62_;
  wire _63_;
  wire _64_;
  wire _65_;
  wire [1:0] _66_;
  wire [29:0] _67_;
  wire [63:0] _68_;
  wire _69_;
  wire _70_;
  wire _71_;
  wire _72_;
  wire _73_;
  wire _74_;
  wire _75_;
  wire _76_;
  wire _77_;
  wire _78_;
  wire _79_;
  wire [6:0] _80_;
  wire [31:0] _81_;
  wire [63:0] _82_;
  wire _83_;
  wire _84_;
  wire [7:0] _85_;
  reg _86_;
  reg _87_;
  reg _88_;
  reg _89_;
  reg _90_;
  reg _91_;
  reg [6:0] _92_;
  reg [31:0] _93_ = 32'd0;
  reg [63:0] _94_ = 64'h0000000000000000;
  reg _95_;
  reg _96_;
  reg [7:0] _97_ = 8'h00;
  wire _98_;
  wire _99_;
  input clk;
  wire clk;
  output core_rst;
  wire core_rst;
  output core_stop;
  wire core_stop;
  input core_stopped;
  wire core_stopped;
  input dbg_gpr_ack;
  wire dbg_gpr_ack;
  output [6:0] dbg_gpr_addr;
  wire [6:0] dbg_gpr_addr;
  input [63:0] dbg_gpr_data;
  wire [63:0] dbg_gpr_data;
  output dbg_gpr_req;
  wire dbg_gpr_req;
  output dmi_ack;
  wire dmi_ack;
  input [3:0] dmi_addr;
  wire [3:0] dmi_addr;
  input [63:0] dmi_din;
  wire [63:0] dmi_din;
  output [63:0] dmi_dout;
  wire [63:0] dmi_dout;
  wire dmi_read_log_data;
  wire dmi_read_log_data_1;
  input dmi_req;
  wire dmi_req;
  wire dmi_req_1;
  input dmi_wr;
  wire dmi_wr;
  wire do_icreset;
  wire do_log_trigger;
  wire do_reset;
  wire do_step;
  wire [6:0] gspr_index;
  output icache_rst;
  wire icache_rst;
  input [255:0] log_data;
  wire [255:0] log_data;
  wire [31:0] log_dmi_addr;
  wire [63:0] log_dmi_data;
  wire [63:0] log_dmi_trigger;
  input [31:0] log_read_addr;
  wire [31:0] log_read_addr;
  output [63:0] log_read_data;
  wire [63:0] log_read_data;
  wire [7:0] log_trigger_delay;
  output [31:0] log_write_addr;
  wire [31:0] log_write_addr;
  input [63:0] msr;
  wire [63:0] msr;
  input [63:0] nia;
  wire [63:0] nia;
  input rst;
  wire rst;
  wire [63:0] stat_reg;
  wire stopping;
  input terminate;
  wire terminate;
  wire terminated;
  output terminated_out;
  wire terminated_out;
  assign _00_ = dmi_addr != 4'h5;
  assign _01_ = _00_ ? dmi_req : dbg_gpr_ack;
  assign _02_ = dmi_addr == 4'h5;
  assign _03_ = _02_ ? dmi_req : 1'h0;
  assign _04_ = dmi_addr == 4'h1;
  assign _05_ = dmi_addr == 4'h2;
  assign _06_ = dmi_addr == 4'h3;
  assign _07_ = dmi_addr == 4'h5;
  assign _08_ = dmi_addr == 4'h6;
  assign _09_ = dmi_addr == 4'h7;
  assign _10_ = dmi_addr == 4'h8;
  function [63:0] \26470 ;
    input [63:0] a;
    input [447:0] b;
    input [6:0] s;
    (* parallel_case *)
    casez (s)
      7'b??????1:
        \26470  = b[63:0];
      7'b?????1?:
        \26470  = b[127:64];
      7'b????1??:
        \26470  = b[191:128];
      7'b???1???:
        \26470  = b[255:192];
      7'b??1????:
        \26470  = b[319:256];
      7'b?1?????:
        \26470  = b[383:320];
      7'b1??????:
        \26470  = b[447:384];
      default:
        \26470  = a;
    endcase
  endfunction
  assign _11_ = \26470 (64'h0000000000000000, { log_dmi_trigger, log_dmi_data, 32'h00000001, log_dmi_addr, dbg_gpr_data, msr, nia, stat_reg }, { _10_, _09_, _08_, _07_, _06_, _05_, _04_ });
  assign _12_ = { 24'h000000, log_trigger_delay } != 32'd0;
  assign _13_ = do_log_trigger | _12_;
  assign _14_ = { 24'h000000, log_trigger_delay } == 32'd255;
  assign _15_ = { 24'h000000, log_trigger_delay } + 32'd1;
  assign _16_ = _18_ ? 1'h1 : log_dmi_trigger[1];
  assign _17_ = _14_ ? 8'h00 : _15_[7:0];
  assign _18_ = _13_ & _14_;
  assign _19_ = _13_ ? _17_ : log_trigger_delay;
  assign _20_ = ~ dmi_req_1;
  assign _21_ = dmi_req & _20_;
  assign _22_ = dmi_addr == 4'h0;
  assign _23_ = dmi_din[1] ? 1'h1 : 1'h0;
  assign _24_ = dmi_din[1] ? 1'h0 : terminated;
  assign _25_ = dmi_din[0] ? 1'h1 : stopping;
  assign _26_ = dmi_din[3] ? 1'h1 : 1'h0;
  assign _27_ = dmi_din[3] ? 1'h0 : _24_;
  assign _28_ = dmi_din[2] ? 1'h1 : 1'h0;
  assign _29_ = dmi_din[4] ? 1'h0 : _25_;
  assign _30_ = dmi_din[4] ? 1'h0 : _27_;
  assign _31_ = dmi_addr == 4'h4;
  assign _32_ = dmi_addr == 4'h6;
  assign _33_ = dmi_addr == 4'h8;
  assign _34_ = _33_ ? dmi_din : { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] };
  assign _35_ = _32_ ? dmi_din[31:0] : log_dmi_addr;
  assign _36_ = _32_ ? { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] } : _34_;
  assign _37_ = _31_ ? dmi_din[6:0] : gspr_index;
  assign _38_ = _31_ ? log_dmi_addr : _35_;
  assign _39_ = _31_ ? { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] } : _36_;
  assign _40_ = _60_ ? _29_ : stopping;
  assign _41_ = _22_ ? _26_ : 1'h0;
  assign _42_ = _22_ ? _23_ : 1'h0;
  assign _43_ = _22_ ? _28_ : 1'h0;
  assign _44_ = _64_ ? _30_ : terminated;
  assign _45_ = _22_ ? gspr_index : _37_;
  assign _46_ = _22_ ? log_dmi_addr : _38_;
  assign _47_ = _22_ ? { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] } : _39_;
  assign _48_ = dmi_wr & _22_;
  assign _49_ = dmi_wr ? _41_ : 1'h0;
  assign _50_ = dmi_wr ? _42_ : 1'h0;
  assign _51_ = dmi_wr ? _43_ : 1'h0;
  assign _52_ = dmi_wr & _22_;
  assign _53_ = _65_ ? _45_ : gspr_index;
  assign _54_ = dmi_wr ? _46_ : log_dmi_addr;
  assign _55_ = dmi_wr ? _47_ : { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] };
  assign _56_ = ~ dmi_read_log_data;
  assign _57_ = _56_ & dmi_read_log_data_1;
  assign _58_ = log_dmi_addr[1:0] + 2'h1;
  assign _59_ = _57_ ? _58_ : log_dmi_addr[1:0];
  assign _60_ = _21_ & _48_;
  assign _61_ = _21_ ? _49_ : 1'h0;
  assign _62_ = _21_ ? _50_ : 1'h0;
  assign _63_ = _21_ ? _51_ : 1'h0;
  assign _64_ = _21_ & _52_;
  assign _65_ = _21_ & dmi_wr;
  assign _66_ = _21_ ? _54_[1:0] : _59_;
  assign _67_ = _21_ ? _54_[31:2] : log_dmi_addr[31:2];
  assign _68_ = _21_ ? _55_ : { log_dmi_trigger[63:2], _16_, log_dmi_trigger[0] };
  assign _69_ = dmi_addr == 4'h7;
  assign _70_ = dmi_req & _69_;
  assign _71_ = _70_ ? 1'h1 : 1'h0;
  assign _72_ = terminate ? 1'h1 : _40_;
  assign _73_ = terminate ? 1'h1 : _44_;
  assign _74_ = rst ? dmi_req_1 : dmi_req;
  assign _75_ = rst ? 1'h0 : _72_;
  assign _76_ = rst ? 1'h0 : _61_;
  assign _77_ = rst ? 1'h0 : _62_;
  assign _78_ = rst ? 1'h0 : _63_;
  assign _79_ = rst ? 1'h0 : _73_;
  assign _80_ = rst ? gspr_index : _53_;
  assign _81_ = rst ? log_dmi_addr : { _67_, _66_ };
  assign _82_ = rst ? log_dmi_trigger : _68_;
  assign _83_ = rst ? dmi_read_log_data : _71_;
  assign _84_ = rst ? dmi_read_log_data_1 : dmi_read_log_data;
  assign _85_ = rst ? 8'h00 : _19_;
  always @(posedge clk)
    _86_ <= _74_;
  always @(posedge clk)
    _87_ <= _75_;
  always @(posedge clk)
    _88_ <= _76_;
  always @(posedge clk)
    _89_ <= _77_;
  always @(posedge clk)
    _90_ <= _78_;
  always @(posedge clk)
    _91_ <= _79_;
  always @(posedge clk)
    _92_ <= _80_;
  always @(posedge clk)
    _93_ <= _81_;
  always @(posedge clk)
    _94_ <= _82_;
  always @(posedge clk)
    _95_ <= _83_;
  always @(posedge clk)
    _96_ <= _84_;
  always @(posedge clk)
    _97_ <= _85_;
  assign _98_ = ~ do_step;
  assign _99_ = stopping & _98_;
  assign dmi_req_1 = _86_;
  assign stat_reg = { 61'h0000000000000000, terminated, core_stopped, stopping };
  assign stopping = _87_;
  assign do_step = _88_;
  assign do_reset = _89_;
  assign do_icreset = _90_;
  assign terminated = _91_;
  assign gspr_index = _92_;
  assign log_dmi_addr = _93_;
  assign log_dmi_data = 64'h0000000000000000;
  assign log_dmi_trigger = _94_;
  assign do_log_trigger = 1'h0;
  assign dmi_read_log_data = _95_;
  assign dmi_read_log_data_1 = _96_;
  assign log_trigger_delay = _97_;
  assign dmi_dout = _11_;
  assign dmi_ack = _01_;
  assign core_stop = _99_;
  assign core_rst = do_reset;
  assign icache_rst = do_icreset;
  assign dbg_gpr_req = _03_;
  assign dbg_gpr_addr = gspr_index;
  assign log_read_data = 64'h0000000000000000;
  assign log_write_addr = 32'd1;
  assign terminated_out = terminated;
endmodule