module bsg_mem_1r1w_synth_width_p64_els_p8_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [2:0] w_addr_i;
  input [63:0] w_data_i;
  input [2:0] r_addr_i;
  output [63:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [63:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45;
  wire [511:0] mem;
  reg mem_511_sv2v_reg,mem_510_sv2v_reg,mem_509_sv2v_reg,mem_508_sv2v_reg,
  mem_507_sv2v_reg,mem_506_sv2v_reg,mem_505_sv2v_reg,mem_504_sv2v_reg,mem_503_sv2v_reg,
  mem_502_sv2v_reg,mem_501_sv2v_reg,mem_500_sv2v_reg,mem_499_sv2v_reg,mem_498_sv2v_reg,
  mem_497_sv2v_reg,mem_496_sv2v_reg,mem_495_sv2v_reg,mem_494_sv2v_reg,
  mem_493_sv2v_reg,mem_492_sv2v_reg,mem_491_sv2v_reg,mem_490_sv2v_reg,mem_489_sv2v_reg,
  mem_488_sv2v_reg,mem_487_sv2v_reg,mem_486_sv2v_reg,mem_485_sv2v_reg,mem_484_sv2v_reg,
  mem_483_sv2v_reg,mem_482_sv2v_reg,mem_481_sv2v_reg,mem_480_sv2v_reg,
  mem_479_sv2v_reg,mem_478_sv2v_reg,mem_477_sv2v_reg,mem_476_sv2v_reg,mem_475_sv2v_reg,
  mem_474_sv2v_reg,mem_473_sv2v_reg,mem_472_sv2v_reg,mem_471_sv2v_reg,mem_470_sv2v_reg,
  mem_469_sv2v_reg,mem_468_sv2v_reg,mem_467_sv2v_reg,mem_466_sv2v_reg,mem_465_sv2v_reg,
  mem_464_sv2v_reg,mem_463_sv2v_reg,mem_462_sv2v_reg,mem_461_sv2v_reg,
  mem_460_sv2v_reg,mem_459_sv2v_reg,mem_458_sv2v_reg,mem_457_sv2v_reg,mem_456_sv2v_reg,
  mem_455_sv2v_reg,mem_454_sv2v_reg,mem_453_sv2v_reg,mem_452_sv2v_reg,mem_451_sv2v_reg,
  mem_450_sv2v_reg,mem_449_sv2v_reg,mem_448_sv2v_reg,mem_447_sv2v_reg,
  mem_446_sv2v_reg,mem_445_sv2v_reg,mem_444_sv2v_reg,mem_443_sv2v_reg,mem_442_sv2v_reg,
  mem_441_sv2v_reg,mem_440_sv2v_reg,mem_439_sv2v_reg,mem_438_sv2v_reg,mem_437_sv2v_reg,
  mem_436_sv2v_reg,mem_435_sv2v_reg,mem_434_sv2v_reg,mem_433_sv2v_reg,mem_432_sv2v_reg,
  mem_431_sv2v_reg,mem_430_sv2v_reg,mem_429_sv2v_reg,mem_428_sv2v_reg,
  mem_427_sv2v_reg,mem_426_sv2v_reg,mem_425_sv2v_reg,mem_424_sv2v_reg,mem_423_sv2v_reg,
  mem_422_sv2v_reg,mem_421_sv2v_reg,mem_420_sv2v_reg,mem_419_sv2v_reg,mem_418_sv2v_reg,
  mem_417_sv2v_reg,mem_416_sv2v_reg,mem_415_sv2v_reg,mem_414_sv2v_reg,
  mem_413_sv2v_reg,mem_412_sv2v_reg,mem_411_sv2v_reg,mem_410_sv2v_reg,mem_409_sv2v_reg,
  mem_408_sv2v_reg,mem_407_sv2v_reg,mem_406_sv2v_reg,mem_405_sv2v_reg,mem_404_sv2v_reg,
  mem_403_sv2v_reg,mem_402_sv2v_reg,mem_401_sv2v_reg,mem_400_sv2v_reg,
  mem_399_sv2v_reg,mem_398_sv2v_reg,mem_397_sv2v_reg,mem_396_sv2v_reg,mem_395_sv2v_reg,
  mem_394_sv2v_reg,mem_393_sv2v_reg,mem_392_sv2v_reg,mem_391_sv2v_reg,mem_390_sv2v_reg,
  mem_389_sv2v_reg,mem_388_sv2v_reg,mem_387_sv2v_reg,mem_386_sv2v_reg,mem_385_sv2v_reg,
  mem_384_sv2v_reg,mem_383_sv2v_reg,mem_382_sv2v_reg,mem_381_sv2v_reg,
  mem_380_sv2v_reg,mem_379_sv2v_reg,mem_378_sv2v_reg,mem_377_sv2v_reg,mem_376_sv2v_reg,
  mem_375_sv2v_reg,mem_374_sv2v_reg,mem_373_sv2v_reg,mem_372_sv2v_reg,mem_371_sv2v_reg,
  mem_370_sv2v_reg,mem_369_sv2v_reg,mem_368_sv2v_reg,mem_367_sv2v_reg,
  mem_366_sv2v_reg,mem_365_sv2v_reg,mem_364_sv2v_reg,mem_363_sv2v_reg,mem_362_sv2v_reg,
  mem_361_sv2v_reg,mem_360_sv2v_reg,mem_359_sv2v_reg,mem_358_sv2v_reg,mem_357_sv2v_reg,
  mem_356_sv2v_reg,mem_355_sv2v_reg,mem_354_sv2v_reg,mem_353_sv2v_reg,mem_352_sv2v_reg,
  mem_351_sv2v_reg,mem_350_sv2v_reg,mem_349_sv2v_reg,mem_348_sv2v_reg,
  mem_347_sv2v_reg,mem_346_sv2v_reg,mem_345_sv2v_reg,mem_344_sv2v_reg,mem_343_sv2v_reg,
  mem_342_sv2v_reg,mem_341_sv2v_reg,mem_340_sv2v_reg,mem_339_sv2v_reg,mem_338_sv2v_reg,
  mem_337_sv2v_reg,mem_336_sv2v_reg,mem_335_sv2v_reg,mem_334_sv2v_reg,
  mem_333_sv2v_reg,mem_332_sv2v_reg,mem_331_sv2v_reg,mem_330_sv2v_reg,mem_329_sv2v_reg,
  mem_328_sv2v_reg,mem_327_sv2v_reg,mem_326_sv2v_reg,mem_325_sv2v_reg,mem_324_sv2v_reg,
  mem_323_sv2v_reg,mem_322_sv2v_reg,mem_321_sv2v_reg,mem_320_sv2v_reg,
  mem_319_sv2v_reg,mem_318_sv2v_reg,mem_317_sv2v_reg,mem_316_sv2v_reg,mem_315_sv2v_reg,
  mem_314_sv2v_reg,mem_313_sv2v_reg,mem_312_sv2v_reg,mem_311_sv2v_reg,mem_310_sv2v_reg,
  mem_309_sv2v_reg,mem_308_sv2v_reg,mem_307_sv2v_reg,mem_306_sv2v_reg,mem_305_sv2v_reg,
  mem_304_sv2v_reg,mem_303_sv2v_reg,mem_302_sv2v_reg,mem_301_sv2v_reg,
  mem_300_sv2v_reg,mem_299_sv2v_reg,mem_298_sv2v_reg,mem_297_sv2v_reg,mem_296_sv2v_reg,
  mem_295_sv2v_reg,mem_294_sv2v_reg,mem_293_sv2v_reg,mem_292_sv2v_reg,mem_291_sv2v_reg,
  mem_290_sv2v_reg,mem_289_sv2v_reg,mem_288_sv2v_reg,mem_287_sv2v_reg,
  mem_286_sv2v_reg,mem_285_sv2v_reg,mem_284_sv2v_reg,mem_283_sv2v_reg,mem_282_sv2v_reg,
  mem_281_sv2v_reg,mem_280_sv2v_reg,mem_279_sv2v_reg,mem_278_sv2v_reg,mem_277_sv2v_reg,
  mem_276_sv2v_reg,mem_275_sv2v_reg,mem_274_sv2v_reg,mem_273_sv2v_reg,mem_272_sv2v_reg,
  mem_271_sv2v_reg,mem_270_sv2v_reg,mem_269_sv2v_reg,mem_268_sv2v_reg,
  mem_267_sv2v_reg,mem_266_sv2v_reg,mem_265_sv2v_reg,mem_264_sv2v_reg,mem_263_sv2v_reg,
  mem_262_sv2v_reg,mem_261_sv2v_reg,mem_260_sv2v_reg,mem_259_sv2v_reg,mem_258_sv2v_reg,
  mem_257_sv2v_reg,mem_256_sv2v_reg,mem_255_sv2v_reg,mem_254_sv2v_reg,
  mem_253_sv2v_reg,mem_252_sv2v_reg,mem_251_sv2v_reg,mem_250_sv2v_reg,mem_249_sv2v_reg,
  mem_248_sv2v_reg,mem_247_sv2v_reg,mem_246_sv2v_reg,mem_245_sv2v_reg,mem_244_sv2v_reg,
  mem_243_sv2v_reg,mem_242_sv2v_reg,mem_241_sv2v_reg,mem_240_sv2v_reg,
  mem_239_sv2v_reg,mem_238_sv2v_reg,mem_237_sv2v_reg,mem_236_sv2v_reg,mem_235_sv2v_reg,
  mem_234_sv2v_reg,mem_233_sv2v_reg,mem_232_sv2v_reg,mem_231_sv2v_reg,mem_230_sv2v_reg,
  mem_229_sv2v_reg,mem_228_sv2v_reg,mem_227_sv2v_reg,mem_226_sv2v_reg,mem_225_sv2v_reg,
  mem_224_sv2v_reg,mem_223_sv2v_reg,mem_222_sv2v_reg,mem_221_sv2v_reg,
  mem_220_sv2v_reg,mem_219_sv2v_reg,mem_218_sv2v_reg,mem_217_sv2v_reg,mem_216_sv2v_reg,
  mem_215_sv2v_reg,mem_214_sv2v_reg,mem_213_sv2v_reg,mem_212_sv2v_reg,mem_211_sv2v_reg,
  mem_210_sv2v_reg,mem_209_sv2v_reg,mem_208_sv2v_reg,mem_207_sv2v_reg,
  mem_206_sv2v_reg,mem_205_sv2v_reg,mem_204_sv2v_reg,mem_203_sv2v_reg,mem_202_sv2v_reg,
  mem_201_sv2v_reg,mem_200_sv2v_reg,mem_199_sv2v_reg,mem_198_sv2v_reg,mem_197_sv2v_reg,
  mem_196_sv2v_reg,mem_195_sv2v_reg,mem_194_sv2v_reg,mem_193_sv2v_reg,mem_192_sv2v_reg,
  mem_191_sv2v_reg,mem_190_sv2v_reg,mem_189_sv2v_reg,mem_188_sv2v_reg,
  mem_187_sv2v_reg,mem_186_sv2v_reg,mem_185_sv2v_reg,mem_184_sv2v_reg,mem_183_sv2v_reg,
  mem_182_sv2v_reg,mem_181_sv2v_reg,mem_180_sv2v_reg,mem_179_sv2v_reg,mem_178_sv2v_reg,
  mem_177_sv2v_reg,mem_176_sv2v_reg,mem_175_sv2v_reg,mem_174_sv2v_reg,
  mem_173_sv2v_reg,mem_172_sv2v_reg,mem_171_sv2v_reg,mem_170_sv2v_reg,mem_169_sv2v_reg,
  mem_168_sv2v_reg,mem_167_sv2v_reg,mem_166_sv2v_reg,mem_165_sv2v_reg,mem_164_sv2v_reg,
  mem_163_sv2v_reg,mem_162_sv2v_reg,mem_161_sv2v_reg,mem_160_sv2v_reg,
  mem_159_sv2v_reg,mem_158_sv2v_reg,mem_157_sv2v_reg,mem_156_sv2v_reg,mem_155_sv2v_reg,
  mem_154_sv2v_reg,mem_153_sv2v_reg,mem_152_sv2v_reg,mem_151_sv2v_reg,mem_150_sv2v_reg,
  mem_149_sv2v_reg,mem_148_sv2v_reg,mem_147_sv2v_reg,mem_146_sv2v_reg,mem_145_sv2v_reg,
  mem_144_sv2v_reg,mem_143_sv2v_reg,mem_142_sv2v_reg,mem_141_sv2v_reg,
  mem_140_sv2v_reg,mem_139_sv2v_reg,mem_138_sv2v_reg,mem_137_sv2v_reg,mem_136_sv2v_reg,
  mem_135_sv2v_reg,mem_134_sv2v_reg,mem_133_sv2v_reg,mem_132_sv2v_reg,mem_131_sv2v_reg,
  mem_130_sv2v_reg,mem_129_sv2v_reg,mem_128_sv2v_reg,mem_127_sv2v_reg,
  mem_126_sv2v_reg,mem_125_sv2v_reg,mem_124_sv2v_reg,mem_123_sv2v_reg,mem_122_sv2v_reg,
  mem_121_sv2v_reg,mem_120_sv2v_reg,mem_119_sv2v_reg,mem_118_sv2v_reg,mem_117_sv2v_reg,
  mem_116_sv2v_reg,mem_115_sv2v_reg,mem_114_sv2v_reg,mem_113_sv2v_reg,mem_112_sv2v_reg,
  mem_111_sv2v_reg,mem_110_sv2v_reg,mem_109_sv2v_reg,mem_108_sv2v_reg,
  mem_107_sv2v_reg,mem_106_sv2v_reg,mem_105_sv2v_reg,mem_104_sv2v_reg,mem_103_sv2v_reg,
  mem_102_sv2v_reg,mem_101_sv2v_reg,mem_100_sv2v_reg,mem_99_sv2v_reg,mem_98_sv2v_reg,
  mem_97_sv2v_reg,mem_96_sv2v_reg,mem_95_sv2v_reg,mem_94_sv2v_reg,mem_93_sv2v_reg,
  mem_92_sv2v_reg,mem_91_sv2v_reg,mem_90_sv2v_reg,mem_89_sv2v_reg,mem_88_sv2v_reg,
  mem_87_sv2v_reg,mem_86_sv2v_reg,mem_85_sv2v_reg,mem_84_sv2v_reg,mem_83_sv2v_reg,
  mem_82_sv2v_reg,mem_81_sv2v_reg,mem_80_sv2v_reg,mem_79_sv2v_reg,mem_78_sv2v_reg,
  mem_77_sv2v_reg,mem_76_sv2v_reg,mem_75_sv2v_reg,mem_74_sv2v_reg,mem_73_sv2v_reg,
  mem_72_sv2v_reg,mem_71_sv2v_reg,mem_70_sv2v_reg,mem_69_sv2v_reg,mem_68_sv2v_reg,
  mem_67_sv2v_reg,mem_66_sv2v_reg,mem_65_sv2v_reg,mem_64_sv2v_reg,mem_63_sv2v_reg,
  mem_62_sv2v_reg,mem_61_sv2v_reg,mem_60_sv2v_reg,mem_59_sv2v_reg,mem_58_sv2v_reg,
  mem_57_sv2v_reg,mem_56_sv2v_reg,mem_55_sv2v_reg,mem_54_sv2v_reg,mem_53_sv2v_reg,
  mem_52_sv2v_reg,mem_51_sv2v_reg,mem_50_sv2v_reg,mem_49_sv2v_reg,mem_48_sv2v_reg,
  mem_47_sv2v_reg,mem_46_sv2v_reg,mem_45_sv2v_reg,mem_44_sv2v_reg,mem_43_sv2v_reg,
  mem_42_sv2v_reg,mem_41_sv2v_reg,mem_40_sv2v_reg,mem_39_sv2v_reg,mem_38_sv2v_reg,
  mem_37_sv2v_reg,mem_36_sv2v_reg,mem_35_sv2v_reg,mem_34_sv2v_reg,mem_33_sv2v_reg,
  mem_32_sv2v_reg,mem_31_sv2v_reg,mem_30_sv2v_reg,mem_29_sv2v_reg,mem_28_sv2v_reg,
  mem_27_sv2v_reg,mem_26_sv2v_reg,mem_25_sv2v_reg,mem_24_sv2v_reg,mem_23_sv2v_reg,
  mem_22_sv2v_reg,mem_21_sv2v_reg,mem_20_sv2v_reg,mem_19_sv2v_reg,mem_18_sv2v_reg,
  mem_17_sv2v_reg,mem_16_sv2v_reg,mem_15_sv2v_reg,mem_14_sv2v_reg,mem_13_sv2v_reg,
  mem_12_sv2v_reg,mem_11_sv2v_reg,mem_10_sv2v_reg,mem_9_sv2v_reg,mem_8_sv2v_reg,
  mem_7_sv2v_reg,mem_6_sv2v_reg,mem_5_sv2v_reg,mem_4_sv2v_reg,mem_3_sv2v_reg,
  mem_2_sv2v_reg,mem_1_sv2v_reg,mem_0_sv2v_reg;
  assign mem[511] = mem_511_sv2v_reg;
  assign mem[510] = mem_510_sv2v_reg;
  assign mem[509] = mem_509_sv2v_reg;
  assign mem[508] = mem_508_sv2v_reg;
  assign mem[507] = mem_507_sv2v_reg;
  assign mem[506] = mem_506_sv2v_reg;
  assign mem[505] = mem_505_sv2v_reg;
  assign mem[504] = mem_504_sv2v_reg;
  assign mem[503] = mem_503_sv2v_reg;
  assign mem[502] = mem_502_sv2v_reg;
  assign mem[501] = mem_501_sv2v_reg;
  assign mem[500] = mem_500_sv2v_reg;
  assign mem[499] = mem_499_sv2v_reg;
  assign mem[498] = mem_498_sv2v_reg;
  assign mem[497] = mem_497_sv2v_reg;
  assign mem[496] = mem_496_sv2v_reg;
  assign mem[495] = mem_495_sv2v_reg;
  assign mem[494] = mem_494_sv2v_reg;
  assign mem[493] = mem_493_sv2v_reg;
  assign mem[492] = mem_492_sv2v_reg;
  assign mem[491] = mem_491_sv2v_reg;
  assign mem[490] = mem_490_sv2v_reg;
  assign mem[489] = mem_489_sv2v_reg;
  assign mem[488] = mem_488_sv2v_reg;
  assign mem[487] = mem_487_sv2v_reg;
  assign mem[486] = mem_486_sv2v_reg;
  assign mem[485] = mem_485_sv2v_reg;
  assign mem[484] = mem_484_sv2v_reg;
  assign mem[483] = mem_483_sv2v_reg;
  assign mem[482] = mem_482_sv2v_reg;
  assign mem[481] = mem_481_sv2v_reg;
  assign mem[480] = mem_480_sv2v_reg;
  assign mem[479] = mem_479_sv2v_reg;
  assign mem[478] = mem_478_sv2v_reg;
  assign mem[477] = mem_477_sv2v_reg;
  assign mem[476] = mem_476_sv2v_reg;
  assign mem[475] = mem_475_sv2v_reg;
  assign mem[474] = mem_474_sv2v_reg;
  assign mem[473] = mem_473_sv2v_reg;
  assign mem[472] = mem_472_sv2v_reg;
  assign mem[471] = mem_471_sv2v_reg;
  assign mem[470] = mem_470_sv2v_reg;
  assign mem[469] = mem_469_sv2v_reg;
  assign mem[468] = mem_468_sv2v_reg;
  assign mem[467] = mem_467_sv2v_reg;
  assign mem[466] = mem_466_sv2v_reg;
  assign mem[465] = mem_465_sv2v_reg;
  assign mem[464] = mem_464_sv2v_reg;
  assign mem[463] = mem_463_sv2v_reg;
  assign mem[462] = mem_462_sv2v_reg;
  assign mem[461] = mem_461_sv2v_reg;
  assign mem[460] = mem_460_sv2v_reg;
  assign mem[459] = mem_459_sv2v_reg;
  assign mem[458] = mem_458_sv2v_reg;
  assign mem[457] = mem_457_sv2v_reg;
  assign mem[456] = mem_456_sv2v_reg;
  assign mem[455] = mem_455_sv2v_reg;
  assign mem[454] = mem_454_sv2v_reg;
  assign mem[453] = mem_453_sv2v_reg;
  assign mem[452] = mem_452_sv2v_reg;
  assign mem[451] = mem_451_sv2v_reg;
  assign mem[450] = mem_450_sv2v_reg;
  assign mem[449] = mem_449_sv2v_reg;
  assign mem[448] = mem_448_sv2v_reg;
  assign mem[447] = mem_447_sv2v_reg;
  assign mem[446] = mem_446_sv2v_reg;
  assign mem[445] = mem_445_sv2v_reg;
  assign mem[444] = mem_444_sv2v_reg;
  assign mem[443] = mem_443_sv2v_reg;
  assign mem[442] = mem_442_sv2v_reg;
  assign mem[441] = mem_441_sv2v_reg;
  assign mem[440] = mem_440_sv2v_reg;
  assign mem[439] = mem_439_sv2v_reg;
  assign mem[438] = mem_438_sv2v_reg;
  assign mem[437] = mem_437_sv2v_reg;
  assign mem[436] = mem_436_sv2v_reg;
  assign mem[435] = mem_435_sv2v_reg;
  assign mem[434] = mem_434_sv2v_reg;
  assign mem[433] = mem_433_sv2v_reg;
  assign mem[432] = mem_432_sv2v_reg;
  assign mem[431] = mem_431_sv2v_reg;
  assign mem[430] = mem_430_sv2v_reg;
  assign mem[429] = mem_429_sv2v_reg;
  assign mem[428] = mem_428_sv2v_reg;
  assign mem[427] = mem_427_sv2v_reg;
  assign mem[426] = mem_426_sv2v_reg;
  assign mem[425] = mem_425_sv2v_reg;
  assign mem[424] = mem_424_sv2v_reg;
  assign mem[423] = mem_423_sv2v_reg;
  assign mem[422] = mem_422_sv2v_reg;
  assign mem[421] = mem_421_sv2v_reg;
  assign mem[420] = mem_420_sv2v_reg;
  assign mem[419] = mem_419_sv2v_reg;
  assign mem[418] = mem_418_sv2v_reg;
  assign mem[417] = mem_417_sv2v_reg;
  assign mem[416] = mem_416_sv2v_reg;
  assign mem[415] = mem_415_sv2v_reg;
  assign mem[414] = mem_414_sv2v_reg;
  assign mem[413] = mem_413_sv2v_reg;
  assign mem[412] = mem_412_sv2v_reg;
  assign mem[411] = mem_411_sv2v_reg;
  assign mem[410] = mem_410_sv2v_reg;
  assign mem[409] = mem_409_sv2v_reg;
  assign mem[408] = mem_408_sv2v_reg;
  assign mem[407] = mem_407_sv2v_reg;
  assign mem[406] = mem_406_sv2v_reg;
  assign mem[405] = mem_405_sv2v_reg;
  assign mem[404] = mem_404_sv2v_reg;
  assign mem[403] = mem_403_sv2v_reg;
  assign mem[402] = mem_402_sv2v_reg;
  assign mem[401] = mem_401_sv2v_reg;
  assign mem[400] = mem_400_sv2v_reg;
  assign mem[399] = mem_399_sv2v_reg;
  assign mem[398] = mem_398_sv2v_reg;
  assign mem[397] = mem_397_sv2v_reg;
  assign mem[396] = mem_396_sv2v_reg;
  assign mem[395] = mem_395_sv2v_reg;
  assign mem[394] = mem_394_sv2v_reg;
  assign mem[393] = mem_393_sv2v_reg;
  assign mem[392] = mem_392_sv2v_reg;
  assign mem[391] = mem_391_sv2v_reg;
  assign mem[390] = mem_390_sv2v_reg;
  assign mem[389] = mem_389_sv2v_reg;
  assign mem[388] = mem_388_sv2v_reg;
  assign mem[387] = mem_387_sv2v_reg;
  assign mem[386] = mem_386_sv2v_reg;
  assign mem[385] = mem_385_sv2v_reg;
  assign mem[384] = mem_384_sv2v_reg;
  assign mem[383] = mem_383_sv2v_reg;
  assign mem[382] = mem_382_sv2v_reg;
  assign mem[381] = mem_381_sv2v_reg;
  assign mem[380] = mem_380_sv2v_reg;
  assign mem[379] = mem_379_sv2v_reg;
  assign mem[378] = mem_378_sv2v_reg;
  assign mem[377] = mem_377_sv2v_reg;
  assign mem[376] = mem_376_sv2v_reg;
  assign mem[375] = mem_375_sv2v_reg;
  assign mem[374] = mem_374_sv2v_reg;
  assign mem[373] = mem_373_sv2v_reg;
  assign mem[372] = mem_372_sv2v_reg;
  assign mem[371] = mem_371_sv2v_reg;
  assign mem[370] = mem_370_sv2v_reg;
  assign mem[369] = mem_369_sv2v_reg;
  assign mem[368] = mem_368_sv2v_reg;
  assign mem[367] = mem_367_sv2v_reg;
  assign mem[366] = mem_366_sv2v_reg;
  assign mem[365] = mem_365_sv2v_reg;
  assign mem[364] = mem_364_sv2v_reg;
  assign mem[363] = mem_363_sv2v_reg;
  assign mem[362] = mem_362_sv2v_reg;
  assign mem[361] = mem_361_sv2v_reg;
  assign mem[360] = mem_360_sv2v_reg;
  assign mem[359] = mem_359_sv2v_reg;
  assign mem[358] = mem_358_sv2v_reg;
  assign mem[357] = mem_357_sv2v_reg;
  assign mem[356] = mem_356_sv2v_reg;
  assign mem[355] = mem_355_sv2v_reg;
  assign mem[354] = mem_354_sv2v_reg;
  assign mem[353] = mem_353_sv2v_reg;
  assign mem[352] = mem_352_sv2v_reg;
  assign mem[351] = mem_351_sv2v_reg;
  assign mem[350] = mem_350_sv2v_reg;
  assign mem[349] = mem_349_sv2v_reg;
  assign mem[348] = mem_348_sv2v_reg;
  assign mem[347] = mem_347_sv2v_reg;
  assign mem[346] = mem_346_sv2v_reg;
  assign mem[345] = mem_345_sv2v_reg;
  assign mem[344] = mem_344_sv2v_reg;
  assign mem[343] = mem_343_sv2v_reg;
  assign mem[342] = mem_342_sv2v_reg;
  assign mem[341] = mem_341_sv2v_reg;
  assign mem[340] = mem_340_sv2v_reg;
  assign mem[339] = mem_339_sv2v_reg;
  assign mem[338] = mem_338_sv2v_reg;
  assign mem[337] = mem_337_sv2v_reg;
  assign mem[336] = mem_336_sv2v_reg;
  assign mem[335] = mem_335_sv2v_reg;
  assign mem[334] = mem_334_sv2v_reg;
  assign mem[333] = mem_333_sv2v_reg;
  assign mem[332] = mem_332_sv2v_reg;
  assign mem[331] = mem_331_sv2v_reg;
  assign mem[330] = mem_330_sv2v_reg;
  assign mem[329] = mem_329_sv2v_reg;
  assign mem[328] = mem_328_sv2v_reg;
  assign mem[327] = mem_327_sv2v_reg;
  assign mem[326] = mem_326_sv2v_reg;
  assign mem[325] = mem_325_sv2v_reg;
  assign mem[324] = mem_324_sv2v_reg;
  assign mem[323] = mem_323_sv2v_reg;
  assign mem[322] = mem_322_sv2v_reg;
  assign mem[321] = mem_321_sv2v_reg;
  assign mem[320] = mem_320_sv2v_reg;
  assign mem[319] = mem_319_sv2v_reg;
  assign mem[318] = mem_318_sv2v_reg;
  assign mem[317] = mem_317_sv2v_reg;
  assign mem[316] = mem_316_sv2v_reg;
  assign mem[315] = mem_315_sv2v_reg;
  assign mem[314] = mem_314_sv2v_reg;
  assign mem[313] = mem_313_sv2v_reg;
  assign mem[312] = mem_312_sv2v_reg;
  assign mem[311] = mem_311_sv2v_reg;
  assign mem[310] = mem_310_sv2v_reg;
  assign mem[309] = mem_309_sv2v_reg;
  assign mem[308] = mem_308_sv2v_reg;
  assign mem[307] = mem_307_sv2v_reg;
  assign mem[306] = mem_306_sv2v_reg;
  assign mem[305] = mem_305_sv2v_reg;
  assign mem[304] = mem_304_sv2v_reg;
  assign mem[303] = mem_303_sv2v_reg;
  assign mem[302] = mem_302_sv2v_reg;
  assign mem[301] = mem_301_sv2v_reg;
  assign mem[300] = mem_300_sv2v_reg;
  assign mem[299] = mem_299_sv2v_reg;
  assign mem[298] = mem_298_sv2v_reg;
  assign mem[297] = mem_297_sv2v_reg;
  assign mem[296] = mem_296_sv2v_reg;
  assign mem[295] = mem_295_sv2v_reg;
  assign mem[294] = mem_294_sv2v_reg;
  assign mem[293] = mem_293_sv2v_reg;
  assign mem[292] = mem_292_sv2v_reg;
  assign mem[291] = mem_291_sv2v_reg;
  assign mem[290] = mem_290_sv2v_reg;
  assign mem[289] = mem_289_sv2v_reg;
  assign mem[288] = mem_288_sv2v_reg;
  assign mem[287] = mem_287_sv2v_reg;
  assign mem[286] = mem_286_sv2v_reg;
  assign mem[285] = mem_285_sv2v_reg;
  assign mem[284] = mem_284_sv2v_reg;
  assign mem[283] = mem_283_sv2v_reg;
  assign mem[282] = mem_282_sv2v_reg;
  assign mem[281] = mem_281_sv2v_reg;
  assign mem[280] = mem_280_sv2v_reg;
  assign mem[279] = mem_279_sv2v_reg;
  assign mem[278] = mem_278_sv2v_reg;
  assign mem[277] = mem_277_sv2v_reg;
  assign mem[276] = mem_276_sv2v_reg;
  assign mem[275] = mem_275_sv2v_reg;
  assign mem[274] = mem_274_sv2v_reg;
  assign mem[273] = mem_273_sv2v_reg;
  assign mem[272] = mem_272_sv2v_reg;
  assign mem[271] = mem_271_sv2v_reg;
  assign mem[270] = mem_270_sv2v_reg;
  assign mem[269] = mem_269_sv2v_reg;
  assign mem[268] = mem_268_sv2v_reg;
  assign mem[267] = mem_267_sv2v_reg;
  assign mem[266] = mem_266_sv2v_reg;
  assign mem[265] = mem_265_sv2v_reg;
  assign mem[264] = mem_264_sv2v_reg;
  assign mem[263] = mem_263_sv2v_reg;
  assign mem[262] = mem_262_sv2v_reg;
  assign mem[261] = mem_261_sv2v_reg;
  assign mem[260] = mem_260_sv2v_reg;
  assign mem[259] = mem_259_sv2v_reg;
  assign mem[258] = mem_258_sv2v_reg;
  assign mem[257] = mem_257_sv2v_reg;
  assign mem[256] = mem_256_sv2v_reg;
  assign mem[255] = mem_255_sv2v_reg;
  assign mem[254] = mem_254_sv2v_reg;
  assign mem[253] = mem_253_sv2v_reg;
  assign mem[252] = mem_252_sv2v_reg;
  assign mem[251] = mem_251_sv2v_reg;
  assign mem[250] = mem_250_sv2v_reg;
  assign mem[249] = mem_249_sv2v_reg;
  assign mem[248] = mem_248_sv2v_reg;
  assign mem[247] = mem_247_sv2v_reg;
  assign mem[246] = mem_246_sv2v_reg;
  assign mem[245] = mem_245_sv2v_reg;
  assign mem[244] = mem_244_sv2v_reg;
  assign mem[243] = mem_243_sv2v_reg;
  assign mem[242] = mem_242_sv2v_reg;
  assign mem[241] = mem_241_sv2v_reg;
  assign mem[240] = mem_240_sv2v_reg;
  assign mem[239] = mem_239_sv2v_reg;
  assign mem[238] = mem_238_sv2v_reg;
  assign mem[237] = mem_237_sv2v_reg;
  assign mem[236] = mem_236_sv2v_reg;
  assign mem[235] = mem_235_sv2v_reg;
  assign mem[234] = mem_234_sv2v_reg;
  assign mem[233] = mem_233_sv2v_reg;
  assign mem[232] = mem_232_sv2v_reg;
  assign mem[231] = mem_231_sv2v_reg;
  assign mem[230] = mem_230_sv2v_reg;
  assign mem[229] = mem_229_sv2v_reg;
  assign mem[228] = mem_228_sv2v_reg;
  assign mem[227] = mem_227_sv2v_reg;
  assign mem[226] = mem_226_sv2v_reg;
  assign mem[225] = mem_225_sv2v_reg;
  assign mem[224] = mem_224_sv2v_reg;
  assign mem[223] = mem_223_sv2v_reg;
  assign mem[222] = mem_222_sv2v_reg;
  assign mem[221] = mem_221_sv2v_reg;
  assign mem[220] = mem_220_sv2v_reg;
  assign mem[219] = mem_219_sv2v_reg;
  assign mem[218] = mem_218_sv2v_reg;
  assign mem[217] = mem_217_sv2v_reg;
  assign mem[216] = mem_216_sv2v_reg;
  assign mem[215] = mem_215_sv2v_reg;
  assign mem[214] = mem_214_sv2v_reg;
  assign mem[213] = mem_213_sv2v_reg;
  assign mem[212] = mem_212_sv2v_reg;
  assign mem[211] = mem_211_sv2v_reg;
  assign mem[210] = mem_210_sv2v_reg;
  assign mem[209] = mem_209_sv2v_reg;
  assign mem[208] = mem_208_sv2v_reg;
  assign mem[207] = mem_207_sv2v_reg;
  assign mem[206] = mem_206_sv2v_reg;
  assign mem[205] = mem_205_sv2v_reg;
  assign mem[204] = mem_204_sv2v_reg;
  assign mem[203] = mem_203_sv2v_reg;
  assign mem[202] = mem_202_sv2v_reg;
  assign mem[201] = mem_201_sv2v_reg;
  assign mem[200] = mem_200_sv2v_reg;
  assign mem[199] = mem_199_sv2v_reg;
  assign mem[198] = mem_198_sv2v_reg;
  assign mem[197] = mem_197_sv2v_reg;
  assign mem[196] = mem_196_sv2v_reg;
  assign mem[195] = mem_195_sv2v_reg;
  assign mem[194] = mem_194_sv2v_reg;
  assign mem[193] = mem_193_sv2v_reg;
  assign mem[192] = mem_192_sv2v_reg;
  assign mem[191] = mem_191_sv2v_reg;
  assign mem[190] = mem_190_sv2v_reg;
  assign mem[189] = mem_189_sv2v_reg;
  assign mem[188] = mem_188_sv2v_reg;
  assign mem[187] = mem_187_sv2v_reg;
  assign mem[186] = mem_186_sv2v_reg;
  assign mem[185] = mem_185_sv2v_reg;
  assign mem[184] = mem_184_sv2v_reg;
  assign mem[183] = mem_183_sv2v_reg;
  assign mem[182] = mem_182_sv2v_reg;
  assign mem[181] = mem_181_sv2v_reg;
  assign mem[180] = mem_180_sv2v_reg;
  assign mem[179] = mem_179_sv2v_reg;
  assign mem[178] = mem_178_sv2v_reg;
  assign mem[177] = mem_177_sv2v_reg;
  assign mem[176] = mem_176_sv2v_reg;
  assign mem[175] = mem_175_sv2v_reg;
  assign mem[174] = mem_174_sv2v_reg;
  assign mem[173] = mem_173_sv2v_reg;
  assign mem[172] = mem_172_sv2v_reg;
  assign mem[171] = mem_171_sv2v_reg;
  assign mem[170] = mem_170_sv2v_reg;
  assign mem[169] = mem_169_sv2v_reg;
  assign mem[168] = mem_168_sv2v_reg;
  assign mem[167] = mem_167_sv2v_reg;
  assign mem[166] = mem_166_sv2v_reg;
  assign mem[165] = mem_165_sv2v_reg;
  assign mem[164] = mem_164_sv2v_reg;
  assign mem[163] = mem_163_sv2v_reg;
  assign mem[162] = mem_162_sv2v_reg;
  assign mem[161] = mem_161_sv2v_reg;
  assign mem[160] = mem_160_sv2v_reg;
  assign mem[159] = mem_159_sv2v_reg;
  assign mem[158] = mem_158_sv2v_reg;
  assign mem[157] = mem_157_sv2v_reg;
  assign mem[156] = mem_156_sv2v_reg;
  assign mem[155] = mem_155_sv2v_reg;
  assign mem[154] = mem_154_sv2v_reg;
  assign mem[153] = mem_153_sv2v_reg;
  assign mem[152] = mem_152_sv2v_reg;
  assign mem[151] = mem_151_sv2v_reg;
  assign mem[150] = mem_150_sv2v_reg;
  assign mem[149] = mem_149_sv2v_reg;
  assign mem[148] = mem_148_sv2v_reg;
  assign mem[147] = mem_147_sv2v_reg;
  assign mem[146] = mem_146_sv2v_reg;
  assign mem[145] = mem_145_sv2v_reg;
  assign mem[144] = mem_144_sv2v_reg;
  assign mem[143] = mem_143_sv2v_reg;
  assign mem[142] = mem_142_sv2v_reg;
  assign mem[141] = mem_141_sv2v_reg;
  assign mem[140] = mem_140_sv2v_reg;
  assign mem[139] = mem_139_sv2v_reg;
  assign mem[138] = mem_138_sv2v_reg;
  assign mem[137] = mem_137_sv2v_reg;
  assign mem[136] = mem_136_sv2v_reg;
  assign mem[135] = mem_135_sv2v_reg;
  assign mem[134] = mem_134_sv2v_reg;
  assign mem[133] = mem_133_sv2v_reg;
  assign mem[132] = mem_132_sv2v_reg;
  assign mem[131] = mem_131_sv2v_reg;
  assign mem[130] = mem_130_sv2v_reg;
  assign mem[129] = mem_129_sv2v_reg;
  assign mem[128] = mem_128_sv2v_reg;
  assign mem[127] = mem_127_sv2v_reg;
  assign mem[126] = mem_126_sv2v_reg;
  assign mem[125] = mem_125_sv2v_reg;
  assign mem[124] = mem_124_sv2v_reg;
  assign mem[123] = mem_123_sv2v_reg;
  assign mem[122] = mem_122_sv2v_reg;
  assign mem[121] = mem_121_sv2v_reg;
  assign mem[120] = mem_120_sv2v_reg;
  assign mem[119] = mem_119_sv2v_reg;
  assign mem[118] = mem_118_sv2v_reg;
  assign mem[117] = mem_117_sv2v_reg;
  assign mem[116] = mem_116_sv2v_reg;
  assign mem[115] = mem_115_sv2v_reg;
  assign mem[114] = mem_114_sv2v_reg;
  assign mem[113] = mem_113_sv2v_reg;
  assign mem[112] = mem_112_sv2v_reg;
  assign mem[111] = mem_111_sv2v_reg;
  assign mem[110] = mem_110_sv2v_reg;
  assign mem[109] = mem_109_sv2v_reg;
  assign mem[108] = mem_108_sv2v_reg;
  assign mem[107] = mem_107_sv2v_reg;
  assign mem[106] = mem_106_sv2v_reg;
  assign mem[105] = mem_105_sv2v_reg;
  assign mem[104] = mem_104_sv2v_reg;
  assign mem[103] = mem_103_sv2v_reg;
  assign mem[102] = mem_102_sv2v_reg;
  assign mem[101] = mem_101_sv2v_reg;
  assign mem[100] = mem_100_sv2v_reg;
  assign mem[99] = mem_99_sv2v_reg;
  assign mem[98] = mem_98_sv2v_reg;
  assign mem[97] = mem_97_sv2v_reg;
  assign mem[96] = mem_96_sv2v_reg;
  assign mem[95] = mem_95_sv2v_reg;
  assign mem[94] = mem_94_sv2v_reg;
  assign mem[93] = mem_93_sv2v_reg;
  assign mem[92] = mem_92_sv2v_reg;
  assign mem[91] = mem_91_sv2v_reg;
  assign mem[90] = mem_90_sv2v_reg;
  assign mem[89] = mem_89_sv2v_reg;
  assign mem[88] = mem_88_sv2v_reg;
  assign mem[87] = mem_87_sv2v_reg;
  assign mem[86] = mem_86_sv2v_reg;
  assign mem[85] = mem_85_sv2v_reg;
  assign mem[84] = mem_84_sv2v_reg;
  assign mem[83] = mem_83_sv2v_reg;
  assign mem[82] = mem_82_sv2v_reg;
  assign mem[81] = mem_81_sv2v_reg;
  assign mem[80] = mem_80_sv2v_reg;
  assign mem[79] = mem_79_sv2v_reg;
  assign mem[78] = mem_78_sv2v_reg;
  assign mem[77] = mem_77_sv2v_reg;
  assign mem[76] = mem_76_sv2v_reg;
  assign mem[75] = mem_75_sv2v_reg;
  assign mem[74] = mem_74_sv2v_reg;
  assign mem[73] = mem_73_sv2v_reg;
  assign mem[72] = mem_72_sv2v_reg;
  assign mem[71] = mem_71_sv2v_reg;
  assign mem[70] = mem_70_sv2v_reg;
  assign mem[69] = mem_69_sv2v_reg;
  assign mem[68] = mem_68_sv2v_reg;
  assign mem[67] = mem_67_sv2v_reg;
  assign mem[66] = mem_66_sv2v_reg;
  assign mem[65] = mem_65_sv2v_reg;
  assign mem[64] = mem_64_sv2v_reg;
  assign mem[63] = mem_63_sv2v_reg;
  assign mem[62] = mem_62_sv2v_reg;
  assign mem[61] = mem_61_sv2v_reg;
  assign mem[60] = mem_60_sv2v_reg;
  assign mem[59] = mem_59_sv2v_reg;
  assign mem[58] = mem_58_sv2v_reg;
  assign mem[57] = mem_57_sv2v_reg;
  assign mem[56] = mem_56_sv2v_reg;
  assign mem[55] = mem_55_sv2v_reg;
  assign mem[54] = mem_54_sv2v_reg;
  assign mem[53] = mem_53_sv2v_reg;
  assign mem[52] = mem_52_sv2v_reg;
  assign mem[51] = mem_51_sv2v_reg;
  assign mem[50] = mem_50_sv2v_reg;
  assign mem[49] = mem_49_sv2v_reg;
  assign mem[48] = mem_48_sv2v_reg;
  assign mem[47] = mem_47_sv2v_reg;
  assign mem[46] = mem_46_sv2v_reg;
  assign mem[45] = mem_45_sv2v_reg;
  assign mem[44] = mem_44_sv2v_reg;
  assign mem[43] = mem_43_sv2v_reg;
  assign mem[42] = mem_42_sv2v_reg;
  assign mem[41] = mem_41_sv2v_reg;
  assign mem[40] = mem_40_sv2v_reg;
  assign mem[39] = mem_39_sv2v_reg;
  assign mem[38] = mem_38_sv2v_reg;
  assign mem[37] = mem_37_sv2v_reg;
  assign mem[36] = mem_36_sv2v_reg;
  assign mem[35] = mem_35_sv2v_reg;
  assign mem[34] = mem_34_sv2v_reg;
  assign mem[33] = mem_33_sv2v_reg;
  assign mem[32] = mem_32_sv2v_reg;
  assign mem[31] = mem_31_sv2v_reg;
  assign mem[30] = mem_30_sv2v_reg;
  assign mem[29] = mem_29_sv2v_reg;
  assign mem[28] = mem_28_sv2v_reg;
  assign mem[27] = mem_27_sv2v_reg;
  assign mem[26] = mem_26_sv2v_reg;
  assign mem[25] = mem_25_sv2v_reg;
  assign mem[24] = mem_24_sv2v_reg;
  assign mem[23] = mem_23_sv2v_reg;
  assign mem[22] = mem_22_sv2v_reg;
  assign mem[21] = mem_21_sv2v_reg;
  assign mem[20] = mem_20_sv2v_reg;
  assign mem[19] = mem_19_sv2v_reg;
  assign mem[18] = mem_18_sv2v_reg;
  assign mem[17] = mem_17_sv2v_reg;
  assign mem[16] = mem_16_sv2v_reg;
  assign mem[15] = mem_15_sv2v_reg;
  assign mem[14] = mem_14_sv2v_reg;
  assign mem[13] = mem_13_sv2v_reg;
  assign mem[12] = mem_12_sv2v_reg;
  assign mem[11] = mem_11_sv2v_reg;
  assign mem[10] = mem_10_sv2v_reg;
  assign mem[9] = mem_9_sv2v_reg;
  assign mem[8] = mem_8_sv2v_reg;
  assign mem[7] = mem_7_sv2v_reg;
  assign mem[6] = mem_6_sv2v_reg;
  assign mem[5] = mem_5_sv2v_reg;
  assign mem[4] = mem_4_sv2v_reg;
  assign mem[3] = mem_3_sv2v_reg;
  assign mem[2] = mem_2_sv2v_reg;
  assign mem[1] = mem_1_sv2v_reg;
  assign mem[0] = mem_0_sv2v_reg;
  assign r_data_o[63] = (N17)? mem[63] : 
                        (N19)? mem[127] : 
                        (N21)? mem[191] : 
                        (N23)? mem[255] : 
                        (N18)? mem[319] : 
                        (N20)? mem[383] : 
                        (N22)? mem[447] : 
                        (N24)? mem[511] : 1'b0;
  assign r_data_o[62] = (N17)? mem[62] : 
                        (N19)? mem[126] : 
                        (N21)? mem[190] : 
                        (N23)? mem[254] : 
                        (N18)? mem[318] : 
                        (N20)? mem[382] : 
                        (N22)? mem[446] : 
                        (N24)? mem[510] : 1'b0;
  assign r_data_o[61] = (N17)? mem[61] : 
                        (N19)? mem[125] : 
                        (N21)? mem[189] : 
                        (N23)? mem[253] : 
                        (N18)? mem[317] : 
                        (N20)? mem[381] : 
                        (N22)? mem[445] : 
                        (N24)? mem[509] : 1'b0;
  assign r_data_o[60] = (N17)? mem[60] : 
                        (N19)? mem[124] : 
                        (N21)? mem[188] : 
                        (N23)? mem[252] : 
                        (N18)? mem[316] : 
                        (N20)? mem[380] : 
                        (N22)? mem[444] : 
                        (N24)? mem[508] : 1'b0;
  assign r_data_o[59] = (N17)? mem[59] : 
                        (N19)? mem[123] : 
                        (N21)? mem[187] : 
                        (N23)? mem[251] : 
                        (N18)? mem[315] : 
                        (N20)? mem[379] : 
                        (N22)? mem[443] : 
                        (N24)? mem[507] : 1'b0;
  assign r_data_o[58] = (N17)? mem[58] : 
                        (N19)? mem[122] : 
                        (N21)? mem[186] : 
                        (N23)? mem[250] : 
                        (N18)? mem[314] : 
                        (N20)? mem[378] : 
                        (N22)? mem[442] : 
                        (N24)? mem[506] : 1'b0;
  assign r_data_o[57] = (N17)? mem[57] : 
                        (N19)? mem[121] : 
                        (N21)? mem[185] : 
                        (N23)? mem[249] : 
                        (N18)? mem[313] : 
                        (N20)? mem[377] : 
                        (N22)? mem[441] : 
                        (N24)? mem[505] : 1'b0;
  assign r_data_o[56] = (N17)? mem[56] : 
                        (N19)? mem[120] : 
                        (N21)? mem[184] : 
                        (N23)? mem[248] : 
                        (N18)? mem[312] : 
                        (N20)? mem[376] : 
                        (N22)? mem[440] : 
                        (N24)? mem[504] : 1'b0;
  assign r_data_o[55] = (N17)? mem[55] : 
                        (N19)? mem[119] : 
                        (N21)? mem[183] : 
                        (N23)? mem[247] : 
                        (N18)? mem[311] : 
                        (N20)? mem[375] : 
                        (N22)? mem[439] : 
                        (N24)? mem[503] : 1'b0;
  assign r_data_o[54] = (N17)? mem[54] : 
                        (N19)? mem[118] : 
                        (N21)? mem[182] : 
                        (N23)? mem[246] : 
                        (N18)? mem[310] : 
                        (N20)? mem[374] : 
                        (N22)? mem[438] : 
                        (N24)? mem[502] : 1'b0;
  assign r_data_o[53] = (N17)? mem[53] : 
                        (N19)? mem[117] : 
                        (N21)? mem[181] : 
                        (N23)? mem[245] : 
                        (N18)? mem[309] : 
                        (N20)? mem[373] : 
                        (N22)? mem[437] : 
                        (N24)? mem[501] : 1'b0;
  assign r_data_o[52] = (N17)? mem[52] : 
                        (N19)? mem[116] : 
                        (N21)? mem[180] : 
                        (N23)? mem[244] : 
                        (N18)? mem[308] : 
                        (N20)? mem[372] : 
                        (N22)? mem[436] : 
                        (N24)? mem[500] : 1'b0;
  assign r_data_o[51] = (N17)? mem[51] : 
                        (N19)? mem[115] : 
                        (N21)? mem[179] : 
                        (N23)? mem[243] : 
                        (N18)? mem[307] : 
                        (N20)? mem[371] : 
                        (N22)? mem[435] : 
                        (N24)? mem[499] : 1'b0;
  assign r_data_o[50] = (N17)? mem[50] : 
                        (N19)? mem[114] : 
                        (N21)? mem[178] : 
                        (N23)? mem[242] : 
                        (N18)? mem[306] : 
                        (N20)? mem[370] : 
                        (N22)? mem[434] : 
                        (N24)? mem[498] : 1'b0;
  assign r_data_o[49] = (N17)? mem[49] : 
                        (N19)? mem[113] : 
                        (N21)? mem[177] : 
                        (N23)? mem[241] : 
                        (N18)? mem[305] : 
                        (N20)? mem[369] : 
                        (N22)? mem[433] : 
                        (N24)? mem[497] : 1'b0;
  assign r_data_o[48] = (N17)? mem[48] : 
                        (N19)? mem[112] : 
                        (N21)? mem[176] : 
                        (N23)? mem[240] : 
                        (N18)? mem[304] : 
                        (N20)? mem[368] : 
                        (N22)? mem[432] : 
                        (N24)? mem[496] : 1'b0;
  assign r_data_o[47] = (N17)? mem[47] : 
                        (N19)? mem[111] : 
                        (N21)? mem[175] : 
                        (N23)? mem[239] : 
                        (N18)? mem[303] : 
                        (N20)? mem[367] : 
                        (N22)? mem[431] : 
                        (N24)? mem[495] : 1'b0;
  assign r_data_o[46] = (N17)? mem[46] : 
                        (N19)? mem[110] : 
                        (N21)? mem[174] : 
                        (N23)? mem[238] : 
                        (N18)? mem[302] : 
                        (N20)? mem[366] : 
                        (N22)? mem[430] : 
                        (N24)? mem[494] : 1'b0;
  assign r_data_o[45] = (N17)? mem[45] : 
                        (N19)? mem[109] : 
                        (N21)? mem[173] : 
                        (N23)? mem[237] : 
                        (N18)? mem[301] : 
                        (N20)? mem[365] : 
                        (N22)? mem[429] : 
                        (N24)? mem[493] : 1'b0;
  assign r_data_o[44] = (N17)? mem[44] : 
                        (N19)? mem[108] : 
                        (N21)? mem[172] : 
                        (N23)? mem[236] : 
                        (N18)? mem[300] : 
                        (N20)? mem[364] : 
                        (N22)? mem[428] : 
                        (N24)? mem[492] : 1'b0;
  assign r_data_o[43] = (N17)? mem[43] : 
                        (N19)? mem[107] : 
                        (N21)? mem[171] : 
                        (N23)? mem[235] : 
                        (N18)? mem[299] : 
                        (N20)? mem[363] : 
                        (N22)? mem[427] : 
                        (N24)? mem[491] : 1'b0;
  assign r_data_o[42] = (N17)? mem[42] : 
                        (N19)? mem[106] : 
                        (N21)? mem[170] : 
                        (N23)? mem[234] : 
                        (N18)? mem[298] : 
                        (N20)? mem[362] : 
                        (N22)? mem[426] : 
                        (N24)? mem[490] : 1'b0;
  assign r_data_o[41] = (N17)? mem[41] : 
                        (N19)? mem[105] : 
                        (N21)? mem[169] : 
                        (N23)? mem[233] : 
                        (N18)? mem[297] : 
                        (N20)? mem[361] : 
                        (N22)? mem[425] : 
                        (N24)? mem[489] : 1'b0;
  assign r_data_o[40] = (N17)? mem[40] : 
                        (N19)? mem[104] : 
                        (N21)? mem[168] : 
                        (N23)? mem[232] : 
                        (N18)? mem[296] : 
                        (N20)? mem[360] : 
                        (N22)? mem[424] : 
                        (N24)? mem[488] : 1'b0;
  assign r_data_o[39] = (N17)? mem[39] : 
                        (N19)? mem[103] : 
                        (N21)? mem[167] : 
                        (N23)? mem[231] : 
                        (N18)? mem[295] : 
                        (N20)? mem[359] : 
                        (N22)? mem[423] : 
                        (N24)? mem[487] : 1'b0;
  assign r_data_o[38] = (N17)? mem[38] : 
                        (N19)? mem[102] : 
                        (N21)? mem[166] : 
                        (N23)? mem[230] : 
                        (N18)? mem[294] : 
                        (N20)? mem[358] : 
                        (N22)? mem[422] : 
                        (N24)? mem[486] : 1'b0;
  assign r_data_o[37] = (N17)? mem[37] : 
                        (N19)? mem[101] : 
                        (N21)? mem[165] : 
                        (N23)? mem[229] : 
                        (N18)? mem[293] : 
                        (N20)? mem[357] : 
                        (N22)? mem[421] : 
                        (N24)? mem[485] : 1'b0;
  assign r_data_o[36] = (N17)? mem[36] : 
                        (N19)? mem[100] : 
                        (N21)? mem[164] : 
                        (N23)? mem[228] : 
                        (N18)? mem[292] : 
                        (N20)? mem[356] : 
                        (N22)? mem[420] : 
                        (N24)? mem[484] : 1'b0;
  assign r_data_o[35] = (N17)? mem[35] : 
                        (N19)? mem[99] : 
                        (N21)? mem[163] : 
                        (N23)? mem[227] : 
                        (N18)? mem[291] : 
                        (N20)? mem[355] : 
                        (N22)? mem[419] : 
                        (N24)? mem[483] : 1'b0;
  assign r_data_o[34] = (N17)? mem[34] : 
                        (N19)? mem[98] : 
                        (N21)? mem[162] : 
                        (N23)? mem[226] : 
                        (N18)? mem[290] : 
                        (N20)? mem[354] : 
                        (N22)? mem[418] : 
                        (N24)? mem[482] : 1'b0;
  assign r_data_o[33] = (N17)? mem[33] : 
                        (N19)? mem[97] : 
                        (N21)? mem[161] : 
                        (N23)? mem[225] : 
                        (N18)? mem[289] : 
                        (N20)? mem[353] : 
                        (N22)? mem[417] : 
                        (N24)? mem[481] : 1'b0;
  assign r_data_o[32] = (N17)? mem[32] : 
                        (N19)? mem[96] : 
                        (N21)? mem[160] : 
                        (N23)? mem[224] : 
                        (N18)? mem[288] : 
                        (N20)? mem[352] : 
                        (N22)? mem[416] : 
                        (N24)? mem[480] : 1'b0;
  assign r_data_o[31] = (N17)? mem[31] : 
                        (N19)? mem[95] : 
                        (N21)? mem[159] : 
                        (N23)? mem[223] : 
                        (N18)? mem[287] : 
                        (N20)? mem[351] : 
                        (N22)? mem[415] : 
                        (N24)? mem[479] : 1'b0;
  assign r_data_o[30] = (N17)? mem[30] : 
                        (N19)? mem[94] : 
                        (N21)? mem[158] : 
                        (N23)? mem[222] : 
                        (N18)? mem[286] : 
                        (N20)? mem[350] : 
                        (N22)? mem[414] : 
                        (N24)? mem[478] : 1'b0;
  assign r_data_o[29] = (N17)? mem[29] : 
                        (N19)? mem[93] : 
                        (N21)? mem[157] : 
                        (N23)? mem[221] : 
                        (N18)? mem[285] : 
                        (N20)? mem[349] : 
                        (N22)? mem[413] : 
                        (N24)? mem[477] : 1'b0;
  assign r_data_o[28] = (N17)? mem[28] : 
                        (N19)? mem[92] : 
                        (N21)? mem[156] : 
                        (N23)? mem[220] : 
                        (N18)? mem[284] : 
                        (N20)? mem[348] : 
                        (N22)? mem[412] : 
                        (N24)? mem[476] : 1'b0;
  assign r_data_o[27] = (N17)? mem[27] : 
                        (N19)? mem[91] : 
                        (N21)? mem[155] : 
                        (N23)? mem[219] : 
                        (N18)? mem[283] : 
                        (N20)? mem[347] : 
                        (N22)? mem[411] : 
                        (N24)? mem[475] : 1'b0;
  assign r_data_o[26] = (N17)? mem[26] : 
                        (N19)? mem[90] : 
                        (N21)? mem[154] : 
                        (N23)? mem[218] : 
                        (N18)? mem[282] : 
                        (N20)? mem[346] : 
                        (N22)? mem[410] : 
                        (N24)? mem[474] : 1'b0;
  assign r_data_o[25] = (N17)? mem[25] : 
                        (N19)? mem[89] : 
                        (N21)? mem[153] : 
                        (N23)? mem[217] : 
                        (N18)? mem[281] : 
                        (N20)? mem[345] : 
                        (N22)? mem[409] : 
                        (N24)? mem[473] : 1'b0;
  assign r_data_o[24] = (N17)? mem[24] : 
                        (N19)? mem[88] : 
                        (N21)? mem[152] : 
                        (N23)? mem[216] : 
                        (N18)? mem[280] : 
                        (N20)? mem[344] : 
                        (N22)? mem[408] : 
                        (N24)? mem[472] : 1'b0;
  assign r_data_o[23] = (N17)? mem[23] : 
                        (N19)? mem[87] : 
                        (N21)? mem[151] : 
                        (N23)? mem[215] : 
                        (N18)? mem[279] : 
                        (N20)? mem[343] : 
                        (N22)? mem[407] : 
                        (N24)? mem[471] : 1'b0;
  assign r_data_o[22] = (N17)? mem[22] : 
                        (N19)? mem[86] : 
                        (N21)? mem[150] : 
                        (N23)? mem[214] : 
                        (N18)? mem[278] : 
                        (N20)? mem[342] : 
                        (N22)? mem[406] : 
                        (N24)? mem[470] : 1'b0;
  assign r_data_o[21] = (N17)? mem[21] : 
                        (N19)? mem[85] : 
                        (N21)? mem[149] : 
                        (N23)? mem[213] : 
                        (N18)? mem[277] : 
                        (N20)? mem[341] : 
                        (N22)? mem[405] : 
                        (N24)? mem[469] : 1'b0;
  assign r_data_o[20] = (N17)? mem[20] : 
                        (N19)? mem[84] : 
                        (N21)? mem[148] : 
                        (N23)? mem[212] : 
                        (N18)? mem[276] : 
                        (N20)? mem[340] : 
                        (N22)? mem[404] : 
                        (N24)? mem[468] : 1'b0;
  assign r_data_o[19] = (N17)? mem[19] : 
                        (N19)? mem[83] : 
                        (N21)? mem[147] : 
                        (N23)? mem[211] : 
                        (N18)? mem[275] : 
                        (N20)? mem[339] : 
                        (N22)? mem[403] : 
                        (N24)? mem[467] : 1'b0;
  assign r_data_o[18] = (N17)? mem[18] : 
                        (N19)? mem[82] : 
                        (N21)? mem[146] : 
                        (N23)? mem[210] : 
                        (N18)? mem[274] : 
                        (N20)? mem[338] : 
                        (N22)? mem[402] : 
                        (N24)? mem[466] : 1'b0;
  assign r_data_o[17] = (N17)? mem[17] : 
                        (N19)? mem[81] : 
                        (N21)? mem[145] : 
                        (N23)? mem[209] : 
                        (N18)? mem[273] : 
                        (N20)? mem[337] : 
                        (N22)? mem[401] : 
                        (N24)? mem[465] : 1'b0;
  assign r_data_o[16] = (N17)? mem[16] : 
                        (N19)? mem[80] : 
                        (N21)? mem[144] : 
                        (N23)? mem[208] : 
                        (N18)? mem[272] : 
                        (N20)? mem[336] : 
                        (N22)? mem[400] : 
                        (N24)? mem[464] : 1'b0;
  assign r_data_o[15] = (N17)? mem[15] : 
                        (N19)? mem[79] : 
                        (N21)? mem[143] : 
                        (N23)? mem[207] : 
                        (N18)? mem[271] : 
                        (N20)? mem[335] : 
                        (N22)? mem[399] : 
                        (N24)? mem[463] : 1'b0;
  assign r_data_o[14] = (N17)? mem[14] : 
                        (N19)? mem[78] : 
                        (N21)? mem[142] : 
                        (N23)? mem[206] : 
                        (N18)? mem[270] : 
                        (N20)? mem[334] : 
                        (N22)? mem[398] : 
                        (N24)? mem[462] : 1'b0;
  assign r_data_o[13] = (N17)? mem[13] : 
                        (N19)? mem[77] : 
                        (N21)? mem[141] : 
                        (N23)? mem[205] : 
                        (N18)? mem[269] : 
                        (N20)? mem[333] : 
                        (N22)? mem[397] : 
                        (N24)? mem[461] : 1'b0;
  assign r_data_o[12] = (N17)? mem[12] : 
                        (N19)? mem[76] : 
                        (N21)? mem[140] : 
                        (N23)? mem[204] : 
                        (N18)? mem[268] : 
                        (N20)? mem[332] : 
                        (N22)? mem[396] : 
                        (N24)? mem[460] : 1'b0;
  assign r_data_o[11] = (N17)? mem[11] : 
                        (N19)? mem[75] : 
                        (N21)? mem[139] : 
                        (N23)? mem[203] : 
                        (N18)? mem[267] : 
                        (N20)? mem[331] : 
                        (N22)? mem[395] : 
                        (N24)? mem[459] : 1'b0;
  assign r_data_o[10] = (N17)? mem[10] : 
                        (N19)? mem[74] : 
                        (N21)? mem[138] : 
                        (N23)? mem[202] : 
                        (N18)? mem[266] : 
                        (N20)? mem[330] : 
                        (N22)? mem[394] : 
                        (N24)? mem[458] : 1'b0;
  assign r_data_o[9] = (N17)? mem[9] : 
                       (N19)? mem[73] : 
                       (N21)? mem[137] : 
                       (N23)? mem[201] : 
                       (N18)? mem[265] : 
                       (N20)? mem[329] : 
                       (N22)? mem[393] : 
                       (N24)? mem[457] : 1'b0;
  assign r_data_o[8] = (N17)? mem[8] : 
                       (N19)? mem[72] : 
                       (N21)? mem[136] : 
                       (N23)? mem[200] : 
                       (N18)? mem[264] : 
                       (N20)? mem[328] : 
                       (N22)? mem[392] : 
                       (N24)? mem[456] : 1'b0;
  assign r_data_o[7] = (N17)? mem[7] : 
                       (N19)? mem[71] : 
                       (N21)? mem[135] : 
                       (N23)? mem[199] : 
                       (N18)? mem[263] : 
                       (N20)? mem[327] : 
                       (N22)? mem[391] : 
                       (N24)? mem[455] : 1'b0;
  assign r_data_o[6] = (N17)? mem[6] : 
                       (N19)? mem[70] : 
                       (N21)? mem[134] : 
                       (N23)? mem[198] : 
                       (N18)? mem[262] : 
                       (N20)? mem[326] : 
                       (N22)? mem[390] : 
                       (N24)? mem[454] : 1'b0;
  assign r_data_o[5] = (N17)? mem[5] : 
                       (N19)? mem[69] : 
                       (N21)? mem[133] : 
                       (N23)? mem[197] : 
                       (N18)? mem[261] : 
                       (N20)? mem[325] : 
                       (N22)? mem[389] : 
                       (N24)? mem[453] : 1'b0;
  assign r_data_o[4] = (N17)? mem[4] : 
                       (N19)? mem[68] : 
                       (N21)? mem[132] : 
                       (N23)? mem[196] : 
                       (N18)? mem[260] : 
                       (N20)? mem[324] : 
                       (N22)? mem[388] : 
                       (N24)? mem[452] : 1'b0;
  assign r_data_o[3] = (N17)? mem[3] : 
                       (N19)? mem[67] : 
                       (N21)? mem[131] : 
                       (N23)? mem[195] : 
                       (N18)? mem[259] : 
                       (N20)? mem[323] : 
                       (N22)? mem[387] : 
                       (N24)? mem[451] : 1'b0;
  assign r_data_o[2] = (N17)? mem[2] : 
                       (N19)? mem[66] : 
                       (N21)? mem[130] : 
                       (N23)? mem[194] : 
                       (N18)? mem[258] : 
                       (N20)? mem[322] : 
                       (N22)? mem[386] : 
                       (N24)? mem[450] : 1'b0;
  assign r_data_o[1] = (N17)? mem[1] : 
                       (N19)? mem[65] : 
                       (N21)? mem[129] : 
                       (N23)? mem[193] : 
                       (N18)? mem[257] : 
                       (N20)? mem[321] : 
                       (N22)? mem[385] : 
                       (N24)? mem[449] : 1'b0;
  assign r_data_o[0] = (N17)? mem[0] : 
                       (N19)? mem[64] : 
                       (N21)? mem[128] : 
                       (N23)? mem[192] : 
                       (N18)? mem[256] : 
                       (N20)? mem[320] : 
                       (N22)? mem[384] : 
                       (N24)? mem[448] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_511_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_510_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_509_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_508_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_507_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_506_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_505_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_504_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_503_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_502_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_501_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_500_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_499_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_498_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_497_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_496_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_495_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_494_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_493_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_492_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_491_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_490_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_489_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_488_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_487_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_486_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_485_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_484_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_483_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_482_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_481_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_480_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_479_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_478_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_477_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_476_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_475_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_474_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_473_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_472_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_471_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_470_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_469_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_468_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_467_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_466_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_465_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_464_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_463_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_462_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_461_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_460_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_459_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_458_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_457_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_456_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_455_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_454_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_453_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_452_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_451_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_450_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_449_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N41) begin
      mem_448_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_447_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_446_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_445_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_444_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_443_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_442_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_441_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_440_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_439_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_438_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_437_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_436_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_435_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_434_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_433_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_432_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_431_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_430_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_429_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_428_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_427_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_426_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_425_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_424_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_423_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_422_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_421_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_420_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_419_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_418_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_417_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_416_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_415_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_414_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_413_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_412_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_411_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_410_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_409_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_408_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_407_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_406_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_405_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_404_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_403_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_402_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_401_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_400_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_399_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_398_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_397_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_396_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_395_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_394_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_393_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_392_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_391_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_390_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_389_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_388_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_387_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_386_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_385_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N40) begin
      mem_384_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_383_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_382_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_381_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_380_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_379_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_378_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_377_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_376_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_375_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_374_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_373_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_372_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_371_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_370_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_369_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_368_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_367_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_366_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_365_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_364_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_363_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_362_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_361_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_360_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_359_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_358_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_357_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_356_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_355_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_354_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_353_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_352_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_351_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_350_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_349_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_348_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_347_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_346_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_345_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_344_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_343_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_342_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_341_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_340_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_339_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_338_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_337_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_336_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_335_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_334_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_333_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_332_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_331_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_330_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_329_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_328_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_327_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_326_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_325_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_324_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_323_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_322_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_321_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N39) begin
      mem_320_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_319_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_318_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_317_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_316_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_315_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_314_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_313_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_312_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_311_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_310_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_309_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_308_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_307_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_306_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_305_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_304_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_303_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_302_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_301_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_300_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_299_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_298_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_297_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_296_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_295_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_294_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_293_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_292_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_291_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_290_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_289_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_288_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_287_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_286_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_285_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_284_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_283_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_282_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_281_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_280_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_279_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_278_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_277_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_276_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_275_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_274_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_273_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_272_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_271_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_270_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_269_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_268_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_267_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_266_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_265_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_264_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_263_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_262_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_261_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_260_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_259_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_258_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_257_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N38) begin
      mem_256_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_255_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_254_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_253_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_252_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_251_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_250_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_249_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_248_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_247_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_246_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_245_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_244_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_243_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_242_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_241_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_240_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_239_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_238_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_237_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_236_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_235_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_234_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_233_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_232_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_231_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_230_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_229_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_228_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_227_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_226_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_225_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_224_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_223_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_222_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_221_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_220_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_219_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_218_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_217_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_216_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_215_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_214_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_213_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_212_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_211_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_210_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_209_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_208_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_207_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_206_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_205_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_204_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_203_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_202_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_201_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_200_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_199_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_198_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_197_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_196_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_195_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_194_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_193_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N37) begin
      mem_192_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_191_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_190_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_189_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_188_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_187_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_186_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_185_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_184_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_183_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_182_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_181_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_180_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_179_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_178_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_177_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_176_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_175_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_174_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_173_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_172_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_171_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_170_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_169_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_168_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_167_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_166_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_165_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_164_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_163_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_162_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_161_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_160_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_159_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_158_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_157_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_156_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_155_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_154_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_153_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_152_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_151_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_150_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_149_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_148_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_147_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_146_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_145_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_144_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_143_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_142_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_141_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_140_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_139_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_138_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_137_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_136_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_135_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_134_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_133_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_132_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_131_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_130_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_129_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N36) begin
      mem_128_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_127_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_126_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_125_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_124_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_123_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_122_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_121_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_120_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_119_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_118_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_117_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_116_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_115_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_114_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_113_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_112_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_111_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_110_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_109_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_108_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_107_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_106_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_105_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_104_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_103_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_102_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_101_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_100_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_99_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_98_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_97_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_96_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_95_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_94_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_93_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_92_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_91_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_90_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_89_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_88_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_87_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_86_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_85_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_84_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_83_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_82_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_81_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_80_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_79_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_78_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_77_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_76_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_75_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_74_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_73_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_72_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_71_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_70_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_69_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_68_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_67_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_66_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_65_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N35) begin
      mem_64_sv2v_reg <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_63_sv2v_reg <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_62_sv2v_reg <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_61_sv2v_reg <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_60_sv2v_reg <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_59_sv2v_reg <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_58_sv2v_reg <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_57_sv2v_reg <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_56_sv2v_reg <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_55_sv2v_reg <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_54_sv2v_reg <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_53_sv2v_reg <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_52_sv2v_reg <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_51_sv2v_reg <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_50_sv2v_reg <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_49_sv2v_reg <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_48_sv2v_reg <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_47_sv2v_reg <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_46_sv2v_reg <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_45_sv2v_reg <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_44_sv2v_reg <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_43_sv2v_reg <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_42_sv2v_reg <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_41_sv2v_reg <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_40_sv2v_reg <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_39_sv2v_reg <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_38_sv2v_reg <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_37_sv2v_reg <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_36_sv2v_reg <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_35_sv2v_reg <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_34_sv2v_reg <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_33_sv2v_reg <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_32_sv2v_reg <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_31_sv2v_reg <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_30_sv2v_reg <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_29_sv2v_reg <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_28_sv2v_reg <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_27_sv2v_reg <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_26_sv2v_reg <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_25_sv2v_reg <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_24_sv2v_reg <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_23_sv2v_reg <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_22_sv2v_reg <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_21_sv2v_reg <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_20_sv2v_reg <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_19_sv2v_reg <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_18_sv2v_reg <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_17_sv2v_reg <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_16_sv2v_reg <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_15_sv2v_reg <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_14_sv2v_reg <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_13_sv2v_reg <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_12_sv2v_reg <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_11_sv2v_reg <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_10_sv2v_reg <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_9_sv2v_reg <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_8_sv2v_reg <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_7_sv2v_reg <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_6_sv2v_reg <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_5_sv2v_reg <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_4_sv2v_reg <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_3_sv2v_reg <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_2_sv2v_reg <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_1_sv2v_reg <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N34) begin
      mem_0_sv2v_reg <= w_data_i[0];
    end 
  end

  assign N42 = w_addr_i[0] & w_addr_i[1];
  assign N33 = N42 & w_addr_i[2];
  assign N43 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N32 = N43 & w_addr_i[2];
  assign N44 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N31 = N44 & w_addr_i[2];
  assign N45 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign N30 = N45 & w_addr_i[2];
  assign N29 = N42 & N4;
  assign N4 = ~w_addr_i[2];
  assign N28 = N43 & N5;
  assign N5 = ~w_addr_i[2];
  assign N27 = N44 & N6;
  assign N6 = ~w_addr_i[2];
  assign N26 = N45 & N7;
  assign N7 = ~w_addr_i[2];
  assign { N41, N40, N39, N38, N37, N36, N35, N34 } = (N8)? { N33, N32, N31, N30, N29, N28, N27, N26 } : 
                                                      (N9)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N8 = w_v_i;
  assign N9 = N25;
  assign N10 = ~r_addr_i[0];
  assign N11 = ~r_addr_i[1];
  assign N12 = N10 & N11;
  assign N13 = N10 & r_addr_i[1];
  assign N14 = r_addr_i[0] & N11;
  assign N15 = r_addr_i[0] & r_addr_i[1];
  assign N16 = ~r_addr_i[2];
  assign N17 = N12 & N16;
  assign N18 = N12 & r_addr_i[2];
  assign N19 = N14 & N16;
  assign N20 = N14 & r_addr_i[2];
  assign N21 = N13 & N16;
  assign N22 = N13 & r_addr_i[2];
  assign N23 = N15 & N16;
  assign N24 = N15 & r_addr_i[2];
  assign N25 = ~w_v_i;

endmodule