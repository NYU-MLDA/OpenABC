module MulDiv
(
  clk,
  reset,
  io_req_ready,
  io_req_valid,
  io_req_bits_fn,
  io_req_bits_dw,
  io_req_bits_in1,
  io_req_bits_in2,
  io_req_bits_tag,
  io_kill,
  io_resp_ready,
  io_resp_valid,
  io_resp_bits_data,
  io_resp_bits_tag
);

  input [3:0] io_req_bits_fn;
  input [63:0] io_req_bits_in1;
  input [63:0] io_req_bits_in2;
  input [4:0] io_req_bits_tag;
  output [63:0] io_resp_bits_data;
  output [4:0] io_resp_bits_tag;
  input clk;
  input reset;
  input io_req_valid;
  input io_req_bits_dw;
  input io_kill;
  input io_resp_ready;
  output io_req_ready;
  output io_resp_valid;
  wire io_req_ready,io_resp_valid,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,
  N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,
  N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,
  N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,
  N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,
  N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,
  N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,
  N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,
  N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,
  N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,
  N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,
  N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,
  N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,
  N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,
  N256,N257,N258,N259,N260,N261,N262,N263,T1,T179_32,T167,T162,T447_0,T153,T11,T12,
  cmdMul,T120,T118,T96,N264,T82,T31,T32,T41,T33,cmdHi,T36,T42,T45,T46,T51_0,
  rhsSigned,T55,T81,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,
  N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,
  N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,
  N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,
  N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,
  N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,
  N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,
  N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,T94,
  T83,N390,T84,lhsSigned,T85,T93,N391,T97,T99,T111,T113,T112,T121,T123,N392,T124,
  T125,N393,N394,T163,T168,T171,T169,T170,N395,T175_0,N396,N397,N398,N399,N400,N401,
  N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,
  N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,
  N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,
  N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,
  N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,
  N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,
  N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,
  N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
  N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
  N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,
  N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,
  N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,
  N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,
  N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,
  N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,
  N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,
  N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,
  N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
  N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,
  N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,
  N786,N787,N789,N790,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,SV2V_UNCONNECTED_1,
  SV2V_UNCONNECTED_2,SV2V_UNCONNECTED_3,SV2V_UNCONNECTED_4,SV2V_UNCONNECTED_5,
  SV2V_UNCONNECTED_6,SV2V_UNCONNECTED_7,SV2V_UNCONNECTED_8,
  SV2V_UNCONNECTED_9,SV2V_UNCONNECTED_10,SV2V_UNCONNECTED_11,SV2V_UNCONNECTED_12,
  SV2V_UNCONNECTED_13,SV2V_UNCONNECTED_14,SV2V_UNCONNECTED_15,
  SV2V_UNCONNECTED_16,SV2V_UNCONNECTED_17,SV2V_UNCONNECTED_18,
  SV2V_UNCONNECTED_19,SV2V_UNCONNECTED_20,SV2V_UNCONNECTED_21,SV2V_UNCONNECTED_22,
  SV2V_UNCONNECTED_23,SV2V_UNCONNECTED_24,SV2V_UNCONNECTED_25,
  SV2V_UNCONNECTED_26,SV2V_UNCONNECTED_27,SV2V_UNCONNECTED_28,
  SV2V_UNCONNECTED_29,SV2V_UNCONNECTED_30,SV2V_UNCONNECTED_31,SV2V_UNCONNECTED_32,
  SV2V_UNCONNECTED_33,SV2V_UNCONNECTED_34,SV2V_UNCONNECTED_35,
  SV2V_UNCONNECTED_36,SV2V_UNCONNECTED_37,SV2V_UNCONNECTED_38,
  SV2V_UNCONNECTED_39,SV2V_UNCONNECTED_40,SV2V_UNCONNECTED_41,SV2V_UNCONNECTED_42,
  SV2V_UNCONNECTED_43,SV2V_UNCONNECTED_44,SV2V_UNCONNECTED_45,
  SV2V_UNCONNECTED_46,SV2V_UNCONNECTED_47,SV2V_UNCONNECTED_48,
  SV2V_UNCONNECTED_49,SV2V_UNCONNECTED_50,SV2V_UNCONNECTED_51,SV2V_UNCONNECTED_52,
  SV2V_UNCONNECTED_53,SV2V_UNCONNECTED_54,SV2V_UNCONNECTED_55,
  SV2V_UNCONNECTED_56,SV2V_UNCONNECTED_57,SV2V_UNCONNECTED_58,
  SV2V_UNCONNECTED_59,SV2V_UNCONNECTED_60,SV2V_UNCONNECTED_61,SV2V_UNCONNECTED_62,
  SV2V_UNCONNECTED_63,SV2V_UNCONNECTED_64;
  wire [63:63] T179;
  wire [63:32] T449;
  wire [126:0] T448;
  wire [128:65] T447;
  wire [63:0] T130,T188,T101,T102,T103,T147;
  wire [1:0] T122,T252,T253,T377,T378;
  wire [2:0] T116,T248,T249,T250,T251,T373,T374,T375,T376;
  wire [2:1] T95;
  wire [0:0] T28,T117,T450;
  wire [64:0] subtractor;
  wire [64:32] T48;
  wire [31:31] T51,T175;
  wire [5:0] T191,T72,T77,T192,T193,T194,T195,T196,T197,T198,T199,T200,T201,T202,T203,T204,
  T205,T206,T207,T208,T209,T210,T211,T212,T213,T214,T215,T216,T217,T218,T219,T220,
  T221,T222,T223,T317,T318,T319,T320,T321,T322,T323,T324,T325,T326,T327,T328,T329,
  T330,T331,T332,T333,T334,T335,T336,T337,T338,T339,T340,T341,T342,T343,T344,T345,
  T346,T347,T348,T148;
  wire [6:0] T70,T69;
  wire [4:0] T224,T225,T226,T227,T228,T229,T230,T231,T232,T233,T234,T235,T236,T237,T238,T239,
  T349,T350,T351,T352,T353,T354,T355,T356,T357,T358,T359,T360,T361,T362,T363,T364;
  wire [3:0] T240,T241,T242,T243,T244,T245,T246,T247,T365,T366,T367,T368,T369,T370,T371,T372;
  wire [128:56] T136;
  wire [72:0] T142;
  wire [72:72] T444;
  reg [4:0] io_resp_bits_tag;
  reg [128:128] T108;
  reg [64:0] T63;
  reg T3_63_,T3_62_,T3_61_,T3_60_,T3_59_,T3_58_,T3_57_,T3_56_,T3_55_,T3_54_,T3_53_,
  T3_52_,T3_51_,T3_50_,T3_49_,T3_48_,T3_47_,T3_46_,T3_45_,T3_44_,T3_43_,T3_42_,
  T3_41_,T3_40_,T3_39_,T3_38_,T3_37_,T3_36_,T3_35_,T3_34_,T3_33_,T3_32_,isMul,neg_out,
  isHi,T184;
  reg [63:0] io_resp_bits_data,T79;
  reg [2:0] state;
  reg [64:64] T146;
  reg [9:6] T106;
  reg [5:3] T105;
  assign T81 = T192 < T317;
  assign T84 = T450[0] ^ T48[64];
  assign { SV2V_UNCONNECTED_1, T103 } = $signed({ 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 }) >>> { T105, 1'b0, 1'b0, 1'b0 };
  assign T448 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_, io_resp_bits_data[31:0] } << T191;
  assign T170 = 1'b0 < T72;

  always @(posedge clk) begin
    if(T1) begin
      io_resp_bits_tag[4] <= io_req_bits_tag[4];
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      io_resp_bits_tag[3] <= io_req_bits_tag[3];
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      io_resp_bits_tag[2] <= io_req_bits_tag[2];
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      io_resp_bits_tag[1] <= io_req_bits_tag[1];
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      io_resp_bits_tag[0] <= io_req_bits_tag[0];
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T108[128] <= N534;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[64] <= N533;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[63] <= N532;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[62] <= N531;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[61] <= N530;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[60] <= N529;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[59] <= N528;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[58] <= N527;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[57] <= N526;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[56] <= N525;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[55] <= N524;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[54] <= N523;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[53] <= N522;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[52] <= N521;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[51] <= N520;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[50] <= N519;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[49] <= N518;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[48] <= N517;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[47] <= N516;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[46] <= N515;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[45] <= N514;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[44] <= N513;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[43] <= N512;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[42] <= N511;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[41] <= N510;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[40] <= N509;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[39] <= N508;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[38] <= N507;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[37] <= N506;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[36] <= N505;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[35] <= N504;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[34] <= N503;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[33] <= N502;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[32] <= N501;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[31] <= N500;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[30] <= N499;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[29] <= N498;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[28] <= N497;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[27] <= N496;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[26] <= N495;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[25] <= N494;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[24] <= N493;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[23] <= N492;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[22] <= N491;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[21] <= N490;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[20] <= N489;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[19] <= N488;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[18] <= N487;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[17] <= N486;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[16] <= N485;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[15] <= N484;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[14] <= N483;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[13] <= N482;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[12] <= N481;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[11] <= N480;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[10] <= N479;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[9] <= N478;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[8] <= N477;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[7] <= N476;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[6] <= N475;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[5] <= N474;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[4] <= N473;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[3] <= N472;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[2] <= N471;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[1] <= N470;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T63[0] <= N469;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_63_ <= N468;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_62_ <= N467;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_61_ <= N466;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_60_ <= N465;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_59_ <= N464;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_58_ <= N463;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_57_ <= N462;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_56_ <= N461;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_55_ <= N460;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_54_ <= N459;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_53_ <= N458;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_52_ <= N457;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_51_ <= N456;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_50_ <= N455;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_49_ <= N454;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_48_ <= N453;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_47_ <= N452;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_46_ <= N451;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_45_ <= N450;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_44_ <= N449;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_43_ <= N448;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_42_ <= N447;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_41_ <= N446;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_40_ <= N445;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_39_ <= N444;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_38_ <= N443;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_37_ <= N442;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_36_ <= N441;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_35_ <= N440;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_34_ <= N439;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_33_ <= N438;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      T3_32_ <= N437;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      io_resp_bits_data[31] <= N436;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[30] <= N435;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[29] <= N434;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[28] <= N433;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[27] <= N432;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[26] <= N431;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[25] <= N430;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[24] <= N429;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[23] <= N428;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[22] <= N427;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[21] <= N426;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[20] <= N425;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[19] <= N424;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[18] <= N423;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[17] <= N422;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[16] <= N421;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[15] <= N420;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[14] <= N419;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[13] <= N418;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[12] <= N417;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[11] <= N416;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[10] <= N415;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[9] <= N414;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[8] <= N413;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[7] <= N412;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[6] <= N411;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[5] <= N410;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[4] <= N409;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[3] <= N408;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[2] <= N407;
    end 
  end


  always @(posedge clk) begin
    if(N405) begin
      io_resp_bits_data[1] <= N406;
    end 
  end


  always @(posedge clk) begin
    if(N403) begin
      io_resp_bits_data[0] <= N404;
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      isMul <= cmdMul;
    end 
  end


  always @(posedge clk) begin
    if(N543) begin
      state[2] <= N546;
    end 
  end


  always @(posedge clk) begin
    if(N543) begin
      state[1] <= N545;
    end 
  end


  always @(posedge clk) begin
    if(N543) begin
      state[0] <= N544;
    end 
  end


  always @(posedge clk) begin
    if(N549) begin
      neg_out <= N550;
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      isHi <= cmdHi;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T146[64] <= N618;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[63] <= N617;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[62] <= N616;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[61] <= N615;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[60] <= N614;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[59] <= N613;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[58] <= N612;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[57] <= N611;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[56] <= N610;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[55] <= N609;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[54] <= N608;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[53] <= N607;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[52] <= N606;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[51] <= N605;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[50] <= N604;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[49] <= N603;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[48] <= N602;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[47] <= N601;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[46] <= N600;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[45] <= N599;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[44] <= N598;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[43] <= N597;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[42] <= N596;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[41] <= N595;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[40] <= N594;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[39] <= N593;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[38] <= N592;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[37] <= N591;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[36] <= N590;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[35] <= N589;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[34] <= N588;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[33] <= N587;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[32] <= N586;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[31] <= N585;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[30] <= N584;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[29] <= N583;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[28] <= N582;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[27] <= N581;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[26] <= N580;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[25] <= N579;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[24] <= N578;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[23] <= N577;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[22] <= N576;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[21] <= N575;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[20] <= N574;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[19] <= N573;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[18] <= N572;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[17] <= N571;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[16] <= N570;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[15] <= N569;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[14] <= N568;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[13] <= N567;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[12] <= N566;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[11] <= N565;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[10] <= N564;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[9] <= N563;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[8] <= N562;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[7] <= N561;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[6] <= N560;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[5] <= N559;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[4] <= N558;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[3] <= N557;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[2] <= N556;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[1] <= N555;
    end 
  end


  always @(posedge clk) begin
    if(N553) begin
      T79[0] <= N554;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T106[9] <= N630;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T106[8] <= N629;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T106[7] <= N628;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T106[6] <= N627;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T105[5] <= N626;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T105[4] <= N625;
    end 
  end


  always @(posedge clk) begin
    if(N623) begin
      T105[3] <= N624;
    end 
  end


  always @(posedge clk) begin
    if(T1) begin
      T184 <= io_req_bits_dw;
    end 
  end

  assign N670 = ~T184;
  assign { SV2V_UNCONNECTED_2, SV2V_UNCONNECTED_3, SV2V_UNCONNECTED_4, SV2V_UNCONNECTED_5, SV2V_UNCONNECTED_6, SV2V_UNCONNECTED_7, SV2V_UNCONNECTED_8, SV2V_UNCONNECTED_9, SV2V_UNCONNECTED_10, SV2V_UNCONNECTED_11, SV2V_UNCONNECTED_12, SV2V_UNCONNECTED_13, SV2V_UNCONNECTED_14, SV2V_UNCONNECTED_15, SV2V_UNCONNECTED_16, SV2V_UNCONNECTED_17, SV2V_UNCONNECTED_18, SV2V_UNCONNECTED_19, SV2V_UNCONNECTED_20, SV2V_UNCONNECTED_21, SV2V_UNCONNECTED_22, SV2V_UNCONNECTED_23, SV2V_UNCONNECTED_24, SV2V_UNCONNECTED_25, SV2V_UNCONNECTED_26, SV2V_UNCONNECTED_27, SV2V_UNCONNECTED_28, SV2V_UNCONNECTED_29, SV2V_UNCONNECTED_30, SV2V_UNCONNECTED_31, SV2V_UNCONNECTED_32, SV2V_UNCONNECTED_33, SV2V_UNCONNECTED_34, SV2V_UNCONNECTED_35, SV2V_UNCONNECTED_36, SV2V_UNCONNECTED_37, SV2V_UNCONNECTED_38, SV2V_UNCONNECTED_39, SV2V_UNCONNECTED_40, SV2V_UNCONNECTED_41, SV2V_UNCONNECTED_42, SV2V_UNCONNECTED_43, SV2V_UNCONNECTED_44, SV2V_UNCONNECTED_45, SV2V_UNCONNECTED_46, SV2V_UNCONNECTED_47, SV2V_UNCONNECTED_48, SV2V_UNCONNECTED_49, SV2V_UNCONNECTED_50, SV2V_UNCONNECTED_51, SV2V_UNCONNECTED_52, SV2V_UNCONNECTED_53, SV2V_UNCONNECTED_54, SV2V_UNCONNECTED_55, SV2V_UNCONNECTED_56, SV2V_UNCONNECTED_57, SV2V_UNCONNECTED_58, SV2V_UNCONNECTED_59, SV2V_UNCONNECTED_60, SV2V_UNCONNECTED_61, SV2V_UNCONNECTED_62, SV2V_UNCONNECTED_63, SV2V_UNCONNECTED_64, T147 } = { T63[63:1], T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_, io_resp_bits_data[31:0] } >> T148;
  assign N671 = ~state[2];
  assign N672 = state[1] | N671;
  assign N673 = state[0] | N672;
  assign N674 = ~N673;
  assign N675 = ~state[0];
  assign N676 = state[1] | state[2];
  assign N677 = N675 | N676;
  assign N678 = ~N677;
  assign N679 = ~state[1];
  assign N680 = N679 | state[2];
  assign N681 = N675 | N680;
  assign N682 = ~N681;
  assign N683 = io_req_bits_fn[0] | io_req_bits_fn[1];
  assign N684 = ~N683;
  assign N685 = T106[8] | T106[9];
  assign N686 = T106[7] | N685;
  assign N687 = T106[6] | N686;
  assign N688 = T105[5] | N687;
  assign N689 = T105[4] | N688;
  assign N690 = T105[3] | N689;
  assign N691 = ~N690;
  assign N692 = ~io_req_bits_fn[0];
  assign N693 = N692 | io_req_bits_fn[2];
  assign N694 = ~N693;
  assign N695 = io_req_bits_fn[0] | io_req_bits_fn[3];
  assign N696 = ~N695;
  assign N697 = ~io_req_bits_fn[2];
  assign N698 = ~T106[9];
  assign N699 = T106[8] | N698;
  assign N700 = T106[7] | N699;
  assign N701 = T106[6] | N700;
  assign N702 = T105[5] | N701;
  assign N703 = T105[4] | N702;
  assign N704 = T105[3] | N703;
  assign N705 = ~N704;
  assign N706 = N679 | state[2];
  assign N707 = state[0] | N706;
  assign N708 = ~N707;
  assign N709 = ~T105[5];
  assign N710 = ~T105[4];
  assign N711 = ~T105[3];
  assign N712 = T106[8] | T106[9];
  assign N713 = T106[7] | N712;
  assign N714 = T106[6] | N713;
  assign N715 = N709 | N714;
  assign N716 = N710 | N715;
  assign N717 = N711 | N716;
  assign N718 = ~N717;
  assign N719 = T101[62] | T101[63];
  assign N720 = T101[61] | N719;
  assign N721 = T101[60] | N720;
  assign N722 = T101[59] | N721;
  assign N723 = T101[58] | N722;
  assign N724 = T101[57] | N723;
  assign N725 = T101[56] | N724;
  assign N726 = T101[55] | N725;
  assign N727 = T101[54] | N726;
  assign N728 = T101[53] | N727;
  assign N729 = T101[52] | N728;
  assign N730 = T101[51] | N729;
  assign N731 = T101[50] | N730;
  assign N732 = T101[49] | N731;
  assign N733 = T101[48] | N732;
  assign N734 = T101[47] | N733;
  assign N735 = T101[46] | N734;
  assign N736 = T101[45] | N735;
  assign N737 = T101[44] | N736;
  assign N738 = T101[43] | N737;
  assign N739 = T101[42] | N738;
  assign N740 = T101[41] | N739;
  assign N741 = T101[40] | N740;
  assign N742 = T101[39] | N741;
  assign N743 = T101[38] | N742;
  assign N744 = T101[37] | N743;
  assign N745 = T101[36] | N744;
  assign N746 = T101[35] | N745;
  assign N747 = T101[34] | N746;
  assign N748 = T101[33] | N747;
  assign N749 = T101[32] | N748;
  assign N750 = T101[31] | N749;
  assign N751 = T101[30] | N750;
  assign N752 = T101[29] | N751;
  assign N753 = T101[28] | N752;
  assign N754 = T101[27] | N753;
  assign N755 = T101[26] | N754;
  assign N756 = T101[25] | N755;
  assign N757 = T101[24] | N756;
  assign N758 = T101[23] | N757;
  assign N759 = T101[22] | N758;
  assign N760 = T101[21] | N759;
  assign N761 = T101[20] | N760;
  assign N762 = T101[19] | N761;
  assign N763 = T101[18] | N762;
  assign N764 = T101[17] | N763;
  assign N765 = T101[16] | N764;
  assign N766 = T101[15] | N765;
  assign N767 = T101[14] | N766;
  assign N768 = T101[13] | N767;
  assign N769 = T101[12] | N768;
  assign N770 = T101[11] | N769;
  assign N771 = T101[10] | N770;
  assign N772 = T101[9] | N771;
  assign N773 = T101[8] | N772;
  assign N774 = T101[7] | N773;
  assign N775 = T101[6] | N774;
  assign N776 = T101[5] | N775;
  assign N777 = T101[4] | N776;
  assign N778 = T101[3] | N777;
  assign N779 = T101[2] | N778;
  assign N780 = T101[1] | N779;
  assign N781 = T101[0] | N780;
  assign N782 = ~N781;
  assign N783 = N679 | state[2];
  assign N784 = state[0] | N783;
  assign N785 = ~N784;
  assign N786 = state[1] | state[2];
  assign N787 = state[0] | N786;
  assign io_req_ready = ~N787;
  assign N789 = state[1] | N671;
  assign N790 = N675 | N789;
  assign io_resp_valid = ~N790;
  assign N792 = T106[8] | T106[9];
  assign N793 = T106[7] | N792;
  assign N794 = T106[6] | N793;
  assign N795 = T105[5] | N794;
  assign N796 = T105[4] | N795;
  assign N797 = T105[3] | N796;
  assign N798 = ~N797;
  assign N799 = T106[8] | T106[9];
  assign N800 = T106[7] | N799;
  assign N801 = T106[6] | N800;
  assign N802 = N709 | N801;
  assign N803 = N710 | N802;
  assign N804 = N711 | N803;
  assign N805 = T106[8] | T106[9];
  assign N806 = T106[7] | N805;
  assign N807 = T106[6] | N806;
  assign N808 = T105[5] | N807;
  assign N809 = T105[4] | N808;
  assign N810 = T105[3] | N809;
  assign subtractor = T63 - { T146[64:64], T79 };
  assign { T179[63:63], T179_32 } = 1'b0 - io_resp_bits_data[31];
  assign T188 = 1'b0 - { T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_, io_resp_bits_data[31:0] };
  assign T142 = $signed({ T146[64:64], T79 }) * $signed({ 1'b0, io_resp_bits_data[7:0] });
  assign T69 = { T106, T105 } + 1'b1;
  assign T70 = { T106, T105 } + 1'b1;
  assign T148 = 1'b0 - { T105, 1'b0, 1'b0, 1'b0 };
  assign T136 = T142 + { T444[72:72], T444[72:72], T444[72:72], T444[72:72], T444[72:72], T444[72:72], T444[72:72], T444[72:72], T108[128:128], T63[64:1] };
  assign { T51[31:31], T51_0 } = 1'b0 - T48[64];
  assign { T175[31:31], T175_0 } = 1'b0 - T450[0];
  assign T77 = { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } + T317;
  assign T72 = T77 - T192;
  assign io_resp_bits_data[63:32] = (N0)? { T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179[63:63], T179_32 } : 
                                    (N1)? { T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_ } : 1'b0;
  assign N0 = N670;
  assign N1 = T184;
  assign T48[63:32] = (N2)? io_req_bits_in2[63:32] : 
                      (N3)? { T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51[31:31], T51_0 } : 1'b0;
  assign N2 = io_req_bits_dw;
  assign N3 = N395;
  assign T55 = (N2)? io_req_bits_in2[63] : 
               (N3)? io_req_bits_in2[31] : 1'b0;
  assign T191 = (N4)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N5)? T72 : 1'b0;
  assign N4 = T81;
  assign N5 = N265;
  assign T192 = (N6)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N7)? T193 : 1'b0;
  assign N6 = T3_63_;
  assign N7 = N266;
  assign T193 = (N8)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N9)? T194 : 1'b0;
  assign N8 = T3_62_;
  assign N9 = N267;
  assign T194 = (N10)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N11)? T195 : 1'b0;
  assign N10 = T3_61_;
  assign N11 = N268;
  assign T195 = (N12)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N13)? T196 : 1'b0;
  assign N12 = T3_60_;
  assign N13 = N269;
  assign T196 = (N14)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N15)? T197 : 1'b0;
  assign N14 = T3_59_;
  assign N15 = N270;
  assign T197 = (N16)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N17)? T198 : 1'b0;
  assign N16 = T3_58_;
  assign N17 = N271;
  assign T198 = (N18)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N19)? T199 : 1'b0;
  assign N18 = T3_57_;
  assign N19 = N272;
  assign T199 = (N20)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N21)? T200 : 1'b0;
  assign N20 = T3_56_;
  assign N21 = N273;
  assign T200 = (N22)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N23)? T201 : 1'b0;
  assign N22 = T3_55_;
  assign N23 = N274;
  assign T201 = (N24)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N25)? T202 : 1'b0;
  assign N24 = T3_54_;
  assign N25 = N275;
  assign T202 = (N26)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N27)? T203 : 1'b0;
  assign N26 = T3_53_;
  assign N27 = N276;
  assign T203 = (N28)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N29)? T204 : 1'b0;
  assign N28 = T3_52_;
  assign N29 = N277;
  assign T204 = (N30)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N31)? T205 : 1'b0;
  assign N30 = T3_51_;
  assign N31 = N278;
  assign T205 = (N32)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N33)? T206 : 1'b0;
  assign N32 = T3_50_;
  assign N33 = N279;
  assign T206 = (N34)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N35)? T207 : 1'b0;
  assign N34 = T3_49_;
  assign N35 = N280;
  assign T207 = (N36)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N37)? T208 : 1'b0;
  assign N36 = T3_48_;
  assign N37 = N281;
  assign T208 = (N38)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N39)? T209 : 1'b0;
  assign N38 = T3_47_;
  assign N39 = N282;
  assign T209 = (N40)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N41)? T210 : 1'b0;
  assign N40 = T3_46_;
  assign N41 = N283;
  assign T210 = (N42)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N43)? T211 : 1'b0;
  assign N42 = T3_45_;
  assign N43 = N284;
  assign T211 = (N44)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N45)? T212 : 1'b0;
  assign N44 = T3_44_;
  assign N45 = N285;
  assign T212 = (N46)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N47)? T213 : 1'b0;
  assign N46 = T3_43_;
  assign N47 = N286;
  assign T213 = (N48)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N49)? T214 : 1'b0;
  assign N48 = T3_42_;
  assign N49 = N287;
  assign T214 = (N50)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N51)? T215 : 1'b0;
  assign N50 = T3_41_;
  assign N51 = N288;
  assign T215 = (N52)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N53)? T216 : 1'b0;
  assign N52 = T3_40_;
  assign N53 = N289;
  assign T216 = (N54)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N55)? T217 : 1'b0;
  assign N54 = T3_39_;
  assign N55 = N290;
  assign T217 = (N56)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N57)? T218 : 1'b0;
  assign N56 = T3_38_;
  assign N57 = N291;
  assign T218 = (N58)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N59)? T219 : 1'b0;
  assign N58 = T3_37_;
  assign N59 = N292;
  assign T219 = (N60)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N61)? T220 : 1'b0;
  assign N60 = T3_36_;
  assign N61 = N293;
  assign T220 = (N62)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N63)? T221 : 1'b0;
  assign N62 = T3_35_;
  assign N63 = N294;
  assign T221 = (N64)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N65)? T222 : 1'b0;
  assign N64 = T3_34_;
  assign N65 = N295;
  assign T222 = (N66)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N67)? T223 : 1'b0;
  assign N66 = T3_33_;
  assign N67 = N296;
  assign T223[4:0] = (N68)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N69)? T224 : 1'b0;
  assign N68 = T223[5];
  assign N69 = N297;
  assign T224 = (N70)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N71)? T225 : 1'b0;
  assign N70 = io_resp_bits_data[31];
  assign N71 = N298;
  assign T225 = (N72)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N73)? T226 : 1'b0;
  assign N72 = io_resp_bits_data[30];
  assign N73 = N299;
  assign T226 = (N74)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N75)? T227 : 1'b0;
  assign N74 = io_resp_bits_data[29];
  assign N75 = N300;
  assign T227 = (N76)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N77)? T228 : 1'b0;
  assign N76 = io_resp_bits_data[28];
  assign N77 = N301;
  assign T228 = (N78)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N79)? T229 : 1'b0;
  assign N78 = io_resp_bits_data[27];
  assign N79 = N302;
  assign T229 = (N80)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N81)? T230 : 1'b0;
  assign N80 = io_resp_bits_data[26];
  assign N81 = N303;
  assign T230 = (N82)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N83)? T231 : 1'b0;
  assign N82 = io_resp_bits_data[25];
  assign N83 = N304;
  assign T231 = (N84)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N85)? T232 : 1'b0;
  assign N84 = io_resp_bits_data[24];
  assign N85 = N305;
  assign T232 = (N86)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N87)? T233 : 1'b0;
  assign N86 = io_resp_bits_data[23];
  assign N87 = N306;
  assign T233 = (N88)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N89)? T234 : 1'b0;
  assign N88 = io_resp_bits_data[22];
  assign N89 = N307;
  assign T234 = (N90)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N91)? T235 : 1'b0;
  assign N90 = io_resp_bits_data[21];
  assign N91 = N308;
  assign T235 = (N92)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N93)? T236 : 1'b0;
  assign N92 = io_resp_bits_data[20];
  assign N93 = N309;
  assign T236 = (N94)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N95)? T237 : 1'b0;
  assign N94 = io_resp_bits_data[19];
  assign N95 = N310;
  assign T237 = (N96)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N97)? T238 : 1'b0;
  assign N96 = io_resp_bits_data[18];
  assign N97 = N311;
  assign T238 = (N98)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N99)? T239 : 1'b0;
  assign N98 = io_resp_bits_data[17];
  assign N99 = N312;
  assign T239[3:0] = (N100)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N101)? T240 : 1'b0;
  assign N100 = T239[4];
  assign N101 = N313;
  assign T240 = (N102)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N103)? T241 : 1'b0;
  assign N102 = io_resp_bits_data[15];
  assign N103 = N314;
  assign T241 = (N104)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N105)? T242 : 1'b0;
  assign N104 = io_resp_bits_data[14];
  assign N105 = N315;
  assign T242 = (N106)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N107)? T243 : 1'b0;
  assign N106 = io_resp_bits_data[13];
  assign N107 = N316;
  assign T243 = (N108)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N109)? T244 : 1'b0;
  assign N108 = io_resp_bits_data[12];
  assign N109 = N317;
  assign T244 = (N110)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N111)? T245 : 1'b0;
  assign N110 = io_resp_bits_data[11];
  assign N111 = N318;
  assign T245 = (N112)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N113)? T246 : 1'b0;
  assign N112 = io_resp_bits_data[10];
  assign N113 = N319;
  assign T246 = (N114)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N115)? T247 : 1'b0;
  assign N114 = io_resp_bits_data[9];
  assign N115 = N320;
  assign T247[2:0] = (N116)? { 1'b0, 1'b0, 1'b0 } : 
                     (N117)? T248 : 1'b0;
  assign N116 = T247[3];
  assign N117 = N321;
  assign T248 = (N118)? { 1'b1, 1'b1, 1'b1 } : 
                (N119)? T249 : 1'b0;
  assign N118 = io_resp_bits_data[7];
  assign N119 = N322;
  assign T249 = (N120)? { 1'b1, 1'b1, 1'b0 } : 
                (N121)? T250 : 1'b0;
  assign N120 = io_resp_bits_data[6];
  assign N121 = N323;
  assign T250 = (N122)? { 1'b1, 1'b0, 1'b1 } : 
                (N123)? T251 : 1'b0;
  assign N122 = io_resp_bits_data[5];
  assign N123 = N324;
  assign T251[1:0] = (N124)? { 1'b0, 1'b0 } : 
                     (N125)? T252 : 1'b0;
  assign N124 = T251[2];
  assign N125 = N325;
  assign T252 = (N126)? { 1'b1, 1'b1 } : 
                (N127)? T253 : 1'b0;
  assign N126 = io_resp_bits_data[3];
  assign N127 = N326;
  assign T253[0] = (N128)? 1'b0 : 
                   (N129)? io_resp_bits_data[1] : 1'b0;
  assign N128 = T253[1];
  assign N129 = N327;
  assign T317 = (N130)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N131)? T318 : 1'b0;
  assign N130 = T79[63];
  assign N131 = N328;
  assign T318 = (N132)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N133)? T319 : 1'b0;
  assign N132 = T79[62];
  assign N133 = N329;
  assign T319 = (N134)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N135)? T320 : 1'b0;
  assign N134 = T79[61];
  assign N135 = N330;
  assign T320 = (N136)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N137)? T321 : 1'b0;
  assign N136 = T79[60];
  assign N137 = N331;
  assign T321 = (N138)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N139)? T322 : 1'b0;
  assign N138 = T79[59];
  assign N139 = N332;
  assign T322 = (N140)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N141)? T323 : 1'b0;
  assign N140 = T79[58];
  assign N141 = N333;
  assign T323 = (N142)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N143)? T324 : 1'b0;
  assign N142 = T79[57];
  assign N143 = N334;
  assign T324 = (N144)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N145)? T325 : 1'b0;
  assign N144 = T79[56];
  assign N145 = N335;
  assign T325 = (N146)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N147)? T326 : 1'b0;
  assign N146 = T79[55];
  assign N147 = N336;
  assign T326 = (N148)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N149)? T327 : 1'b0;
  assign N148 = T79[54];
  assign N149 = N337;
  assign T327 = (N150)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N151)? T328 : 1'b0;
  assign N150 = T79[53];
  assign N151 = N338;
  assign T328 = (N152)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N153)? T329 : 1'b0;
  assign N152 = T79[52];
  assign N153 = N339;
  assign T329 = (N154)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N155)? T330 : 1'b0;
  assign N154 = T79[51];
  assign N155 = N340;
  assign T330 = (N156)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N157)? T331 : 1'b0;
  assign N156 = T79[50];
  assign N157 = N341;
  assign T331 = (N158)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N159)? T332 : 1'b0;
  assign N158 = T79[49];
  assign N159 = N342;
  assign T332 = (N160)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N161)? T333 : 1'b0;
  assign N160 = T79[48];
  assign N161 = N343;
  assign T333 = (N162)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N163)? T334 : 1'b0;
  assign N162 = T79[47];
  assign N163 = N344;
  assign T334 = (N164)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N165)? T335 : 1'b0;
  assign N164 = T79[46];
  assign N165 = N345;
  assign T335 = (N166)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N167)? T336 : 1'b0;
  assign N166 = T79[45];
  assign N167 = N346;
  assign T336 = (N168)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N169)? T337 : 1'b0;
  assign N168 = T79[44];
  assign N169 = N347;
  assign T337 = (N170)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N171)? T338 : 1'b0;
  assign N170 = T79[43];
  assign N171 = N348;
  assign T338 = (N172)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N173)? T339 : 1'b0;
  assign N172 = T79[42];
  assign N173 = N349;
  assign T339 = (N174)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N175)? T340 : 1'b0;
  assign N174 = T79[41];
  assign N175 = N350;
  assign T340 = (N176)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N177)? T341 : 1'b0;
  assign N176 = T79[40];
  assign N177 = N351;
  assign T341 = (N178)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N179)? T342 : 1'b0;
  assign N178 = T79[39];
  assign N179 = N352;
  assign T342 = (N180)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N181)? T343 : 1'b0;
  assign N180 = T79[38];
  assign N181 = N353;
  assign T343 = (N182)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N183)? T344 : 1'b0;
  assign N182 = T79[37];
  assign N183 = N354;
  assign T344 = (N184)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N185)? T345 : 1'b0;
  assign N184 = T79[36];
  assign N185 = N355;
  assign T345 = (N186)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N187)? T346 : 1'b0;
  assign N186 = T79[35];
  assign N187 = N356;
  assign T346 = (N188)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N189)? T347 : 1'b0;
  assign N188 = T79[34];
  assign N189 = N357;
  assign T347 = (N190)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N191)? T348 : 1'b0;
  assign N190 = T79[33];
  assign N191 = N358;
  assign T348[4:0] = (N192)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N193)? T349 : 1'b0;
  assign N192 = T348[5];
  assign N193 = N359;
  assign T349 = (N194)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N195)? T350 : 1'b0;
  assign N194 = T79[31];
  assign N195 = N360;
  assign T350 = (N196)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N197)? T351 : 1'b0;
  assign N196 = T79[30];
  assign N197 = N361;
  assign T351 = (N198)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N199)? T352 : 1'b0;
  assign N198 = T79[29];
  assign N199 = N362;
  assign T352 = (N200)? { 1'b1, 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N201)? T353 : 1'b0;
  assign N200 = T79[28];
  assign N201 = N363;
  assign T353 = (N202)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N203)? T354 : 1'b0;
  assign N202 = T79[27];
  assign N203 = N364;
  assign T354 = (N204)? { 1'b1, 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N205)? T355 : 1'b0;
  assign N204 = T79[26];
  assign N205 = N365;
  assign T355 = (N206)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N207)? T356 : 1'b0;
  assign N206 = T79[25];
  assign N207 = N366;
  assign T356 = (N208)? { 1'b1, 1'b1, 1'b0, 1'b0, 1'b0 } : 
                (N209)? T357 : 1'b0;
  assign N208 = T79[24];
  assign N209 = N367;
  assign T357 = (N210)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b1 } : 
                (N211)? T358 : 1'b0;
  assign N210 = T79[23];
  assign N211 = N368;
  assign T358 = (N212)? { 1'b1, 1'b0, 1'b1, 1'b1, 1'b0 } : 
                (N213)? T359 : 1'b0;
  assign N212 = T79[22];
  assign N213 = N369;
  assign T359 = (N214)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b1 } : 
                (N215)? T360 : 1'b0;
  assign N214 = T79[21];
  assign N215 = N370;
  assign T360 = (N216)? { 1'b1, 1'b0, 1'b1, 1'b0, 1'b0 } : 
                (N217)? T361 : 1'b0;
  assign N216 = T79[20];
  assign N217 = N371;
  assign T361 = (N218)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b1 } : 
                (N219)? T362 : 1'b0;
  assign N218 = T79[19];
  assign N219 = N372;
  assign T362 = (N220)? { 1'b1, 1'b0, 1'b0, 1'b1, 1'b0 } : 
                (N221)? T363 : 1'b0;
  assign N220 = T79[18];
  assign N221 = N373;
  assign T363 = (N222)? { 1'b1, 1'b0, 1'b0, 1'b0, 1'b1 } : 
                (N223)? T364 : 1'b0;
  assign N222 = T79[17];
  assign N223 = N374;
  assign T364[3:0] = (N224)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 
                     (N225)? T365 : 1'b0;
  assign N224 = T364[4];
  assign N225 = N375;
  assign T365 = (N226)? { 1'b1, 1'b1, 1'b1, 1'b1 } : 
                (N227)? T366 : 1'b0;
  assign N226 = T79[15];
  assign N227 = N376;
  assign T366 = (N228)? { 1'b1, 1'b1, 1'b1, 1'b0 } : 
                (N229)? T367 : 1'b0;
  assign N228 = T79[14];
  assign N229 = N377;
  assign T367 = (N230)? { 1'b1, 1'b1, 1'b0, 1'b1 } : 
                (N231)? T368 : 1'b0;
  assign N230 = T79[13];
  assign N231 = N378;
  assign T368 = (N232)? { 1'b1, 1'b1, 1'b0, 1'b0 } : 
                (N233)? T369 : 1'b0;
  assign N232 = T79[12];
  assign N233 = N379;
  assign T369 = (N234)? { 1'b1, 1'b0, 1'b1, 1'b1 } : 
                (N235)? T370 : 1'b0;
  assign N234 = T79[11];
  assign N235 = N380;
  assign T370 = (N236)? { 1'b1, 1'b0, 1'b1, 1'b0 } : 
                (N237)? T371 : 1'b0;
  assign N236 = T79[10];
  assign N237 = N381;
  assign T371 = (N238)? { 1'b1, 1'b0, 1'b0, 1'b1 } : 
                (N239)? T372 : 1'b0;
  assign N238 = T79[9];
  assign N239 = N382;
  assign T372[2:0] = (N240)? { 1'b0, 1'b0, 1'b0 } : 
                     (N241)? T373 : 1'b0;
  assign N240 = T372[3];
  assign N241 = N383;
  assign T373 = (N242)? { 1'b1, 1'b1, 1'b1 } : 
                (N243)? T374 : 1'b0;
  assign N242 = T79[7];
  assign N243 = N384;
  assign T374 = (N244)? { 1'b1, 1'b1, 1'b0 } : 
                (N245)? T375 : 1'b0;
  assign N244 = T79[6];
  assign N245 = N385;
  assign T375 = (N246)? { 1'b1, 1'b0, 1'b1 } : 
                (N247)? T376 : 1'b0;
  assign N246 = T79[5];
  assign N247 = N386;
  assign T376[1:0] = (N248)? { 1'b0, 1'b0 } : 
                     (N249)? T377 : 1'b0;
  assign N248 = T376[2];
  assign N249 = N387;
  assign T377 = (N250)? { 1'b1, 1'b1 } : 
                (N251)? T378 : 1'b0;
  assign N250 = T79[3];
  assign N251 = N388;
  assign T378[0] = (N252)? 1'b0 : 
                   (N253)? T79[1] : 1'b0;
  assign N252 = T378[1];
  assign N253 = N389;
  assign T83 = (N254)? T450[0] : 
               (N255)? T84 : 1'b0;
  assign N254 = cmdHi;
  assign N255 = N390;
  assign T85 = (N2)? io_req_bits_in1[63] : 
               (N3)? io_req_bits_in1[31] : 1'b0;
  assign T116[0] = (N256)? 1'b1 : 
                   (N257)? T117[0] : 1'b0;
  assign N256 = T116[1];
  assign N257 = T116[2];
  assign T130 = (N258)? T147 : 
                (N259)? { T136[63:56], T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_, io_resp_bits_data[31:8] } : 1'b0;
  assign N258 = T99;
  assign N259 = N393;
  assign T447 = (N260)? T63[63:0] : 
                (N261)? subtractor[63:0] : 1'b0;
  assign N260 = subtractor[64];
  assign N261 = N394;
  assign T449 = (N2)? io_req_bits_in1[63:32] : 
                (N3)? { T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175[31:31], T175_0 } : 1'b0;
  assign { N405, N403 } = (N262)? { 1'b1, 1'b1 } : 
                          (N632)? { 1'b1, 1'b1 } : 
                          (N635)? { 1'b1, 1'b1 } : 
                          (N638)? { 1'b1, 1'b1 } : 
                          (N641)? { 1'b1, 1'b1 } : 
                          (N643)? { 1'b1, 1'b1 } : 
                          (N645)? { 1'b1, 1'b1 } : 
                          (N402)? { 1'b0, 1'b0 } : 1'b0;
  assign N262 = T1;
  assign { N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N404 } = (N262)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T449, io_req_bits_in1[31:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N632)? { 1'b0, 1'b0, 1'b0, T448 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N635)? { 1'b0, T447, T3_63_, T3_62_, T3_61_, T3_60_, T3_59_, T3_58_, T3_57_, T3_56_, T3_55_, T3_54_, T3_53_, T3_52_, T3_51_, T3_50_, T3_49_, T3_48_, T3_47_, T3_46_, T3_45_, T3_44_, T3_43_, T3_42_, T3_41_, T3_40_, T3_39_, T3_38_, T3_37_, T3_36_, T3_35_, T3_34_, T3_33_, T3_32_, io_resp_bits_data[31:0], T447_0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N638)? { T136[128:64], 1'b0, T130 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N641)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T63[64:1] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N643)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T188 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          (N645)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, T188 } : 1'b0;
  assign N543 = (N263)? 1'b1 : 
                (N647)? 1'b1 : 
                (N649)? 1'b1 : 
                (N652)? 1'b1 : 
                (N655)? 1'b1 : 
                (N658)? 1'b1 : 
                (N660)? 1'b1 : 
                (N662)? 1'b1 : 
                (N542)? 1'b0 : 1'b0;
  assign N263 = reset;
  assign { N546, N545, N544 } = (N263)? { 1'b0, 1'b0, 1'b0 } : 
                                (N647)? { 1'b0, T122 } : 
                                (N649)? { 1'b0, 1'b0, 1'b0 } : 
                                (N652)? T116 : 
                                (N655)? { T95, 1'b1 } : 
                                (N658)? { 1'b1, 1'b0, T28[0:0] } : 
                                (N660)? { 1'b1, 1'b0, 1'b1 } : 
                                (N662)? { 1'b0, 1'b1, 1'b0 } : 1'b0;
  assign N549 = (N262)? 1'b1 : 
                (N663)? 1'b1 : 
                (N548)? 1'b0 : 1'b0;
  assign N550 = (N262)? T82 : 
                (N663)? 1'b0 : 1'b0;
  assign N553 = (N262)? 1'b1 : 
                (N664)? 1'b1 : 
                (N552)? 1'b0 : 1'b0;
  assign { N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554 } = (N262)? { T48, io_req_bits_in2[31:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                    (N664)? subtractor : 1'b0;
  assign N623 = (N262)? 1'b1 : 
                (N665)? 1'b1 : 
                (N667)? 1'b1 : 
                (N669)? 1'b1 : 
                (N622)? 1'b0 : 1'b0;
  assign { N630, N629, N628, N627, N626, N625, N624 } = (N262)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N665)? { 1'b0, T191 } : 
                                                        (N667)? T70 : 
                                                        (N669)? T69 : 1'b0;
  assign T1 = io_req_ready & io_req_valid;
  assign T11 = N678 & T12;
  assign T12 = T3_63_ | isMul;
  assign cmdMul = N697 | io_req_bits_fn[3];
  assign N264 = ~neg_out;
  assign T28[0] = N264;
  assign T31 = T162 & T32;
  assign T32 = T41 & T33;
  assign T33 = ~isHi;
  assign cmdHi = T36 | io_req_bits_fn[3];
  assign T36 = N694 | io_req_bits_fn[1];
  assign T41 = N691 & T42;
  assign T42 = ~subtractor[64];
  assign T45 = N678 & T46;
  assign T46 = T79[63] | isMul;
  assign T48[64] = rhsSigned & T55;
  assign rhsSigned = N696 | N697;
  assign N265 = ~T81;
  assign N266 = ~T3_63_;
  assign N267 = ~T3_62_;
  assign N268 = ~T3_61_;
  assign N269 = ~T3_60_;
  assign N270 = ~T3_59_;
  assign N271 = ~T3_58_;
  assign N272 = ~T3_57_;
  assign N273 = ~T3_56_;
  assign N274 = ~T3_55_;
  assign N275 = ~T3_54_;
  assign N276 = ~T3_53_;
  assign N277 = ~T3_52_;
  assign N278 = ~T3_51_;
  assign N279 = ~T3_50_;
  assign N280 = ~T3_49_;
  assign N281 = ~T3_48_;
  assign N282 = ~T3_47_;
  assign N283 = ~T3_46_;
  assign N284 = ~T3_45_;
  assign N285 = ~T3_44_;
  assign N286 = ~T3_43_;
  assign N287 = ~T3_42_;
  assign N288 = ~T3_41_;
  assign N289 = ~T3_40_;
  assign N290 = ~T3_39_;
  assign N291 = ~T3_38_;
  assign N292 = ~T3_37_;
  assign N293 = ~T3_36_;
  assign N294 = ~T3_35_;
  assign N295 = ~T3_34_;
  assign N296 = ~T3_33_;
  assign N297 = ~T3_32_;
  assign T223[5] = T3_32_;
  assign N298 = ~io_resp_bits_data[31];
  assign N299 = ~io_resp_bits_data[30];
  assign N300 = ~io_resp_bits_data[29];
  assign N301 = ~io_resp_bits_data[28];
  assign N302 = ~io_resp_bits_data[27];
  assign N303 = ~io_resp_bits_data[26];
  assign N304 = ~io_resp_bits_data[25];
  assign N305 = ~io_resp_bits_data[24];
  assign N306 = ~io_resp_bits_data[23];
  assign N307 = ~io_resp_bits_data[22];
  assign N308 = ~io_resp_bits_data[21];
  assign N309 = ~io_resp_bits_data[20];
  assign N310 = ~io_resp_bits_data[19];
  assign N311 = ~io_resp_bits_data[18];
  assign N312 = ~io_resp_bits_data[17];
  assign N313 = ~io_resp_bits_data[16];
  assign T239[4] = io_resp_bits_data[16];
  assign N314 = ~io_resp_bits_data[15];
  assign N315 = ~io_resp_bits_data[14];
  assign N316 = ~io_resp_bits_data[13];
  assign N317 = ~io_resp_bits_data[12];
  assign N318 = ~io_resp_bits_data[11];
  assign N319 = ~io_resp_bits_data[10];
  assign N320 = ~io_resp_bits_data[9];
  assign N321 = ~io_resp_bits_data[8];
  assign T247[3] = io_resp_bits_data[8];
  assign N322 = ~io_resp_bits_data[7];
  assign N323 = ~io_resp_bits_data[6];
  assign N324 = ~io_resp_bits_data[5];
  assign N325 = ~io_resp_bits_data[4];
  assign T251[2] = io_resp_bits_data[4];
  assign N326 = ~io_resp_bits_data[3];
  assign N327 = ~io_resp_bits_data[2];
  assign T253[1] = io_resp_bits_data[2];
  assign N328 = ~T79[63];
  assign N329 = ~T79[62];
  assign N330 = ~T79[61];
  assign N331 = ~T79[60];
  assign N332 = ~T79[59];
  assign N333 = ~T79[58];
  assign N334 = ~T79[57];
  assign N335 = ~T79[56];
  assign N336 = ~T79[55];
  assign N337 = ~T79[54];
  assign N338 = ~T79[53];
  assign N339 = ~T79[52];
  assign N340 = ~T79[51];
  assign N341 = ~T79[50];
  assign N342 = ~T79[49];
  assign N343 = ~T79[48];
  assign N344 = ~T79[47];
  assign N345 = ~T79[46];
  assign N346 = ~T79[45];
  assign N347 = ~T79[44];
  assign N348 = ~T79[43];
  assign N349 = ~T79[42];
  assign N350 = ~T79[41];
  assign N351 = ~T79[40];
  assign N352 = ~T79[39];
  assign N353 = ~T79[38];
  assign N354 = ~T79[37];
  assign N355 = ~T79[36];
  assign N356 = ~T79[35];
  assign N357 = ~T79[34];
  assign N358 = ~T79[33];
  assign N359 = ~T79[32];
  assign T348[5] = T79[32];
  assign N360 = ~T79[31];
  assign N361 = ~T79[30];
  assign N362 = ~T79[29];
  assign N363 = ~T79[28];
  assign N364 = ~T79[27];
  assign N365 = ~T79[26];
  assign N366 = ~T79[25];
  assign N367 = ~T79[24];
  assign N368 = ~T79[23];
  assign N369 = ~T79[22];
  assign N370 = ~T79[21];
  assign N371 = ~T79[20];
  assign N372 = ~T79[19];
  assign N373 = ~T79[18];
  assign N374 = ~T79[17];
  assign N375 = ~T79[16];
  assign T364[4] = T79[16];
  assign N376 = ~T79[15];
  assign N377 = ~T79[14];
  assign N378 = ~T79[13];
  assign N379 = ~T79[12];
  assign N380 = ~T79[11];
  assign N381 = ~T79[10];
  assign N382 = ~T79[9];
  assign N383 = ~T79[8];
  assign T372[3] = T79[8];
  assign N384 = ~T79[7];
  assign N385 = ~T79[6];
  assign N386 = ~T79[5];
  assign N387 = ~T79[4];
  assign T376[2] = T79[4];
  assign N388 = ~T79[3];
  assign N389 = ~T79[2];
  assign T378[1] = T79[2];
  assign T82 = T94 & T83;
  assign N390 = ~cmdHi;
  assign T450[0] = lhsSigned & T85;
  assign lhsSigned = T93 | N684;
  assign T93 = N696 | N697;
  assign T94 = ~cmdMul;
  assign N391 = ~isHi;
  assign T95[1] = isHi;
  assign T95[2] = N391;
  assign T96 = T153 & T97;
  assign T97 = T99 | N718;
  assign T99 = T111 & N782;
  assign T101[63] = T3_63_ & T102[63];
  assign T101[62] = T3_62_ & T102[62];
  assign T101[61] = T3_61_ & T102[61];
  assign T101[60] = T3_60_ & T102[60];
  assign T101[59] = T3_59_ & T102[59];
  assign T101[58] = T3_58_ & T102[58];
  assign T101[57] = T3_57_ & T102[57];
  assign T101[56] = T3_56_ & T102[56];
  assign T101[55] = T3_55_ & T102[55];
  assign T101[54] = T3_54_ & T102[54];
  assign T101[53] = T3_53_ & T102[53];
  assign T101[52] = T3_52_ & T102[52];
  assign T101[51] = T3_51_ & T102[51];
  assign T101[50] = T3_50_ & T102[50];
  assign T101[49] = T3_49_ & T102[49];
  assign T101[48] = T3_48_ & T102[48];
  assign T101[47] = T3_47_ & T102[47];
  assign T101[46] = T3_46_ & T102[46];
  assign T101[45] = T3_45_ & T102[45];
  assign T101[44] = T3_44_ & T102[44];
  assign T101[43] = T3_43_ & T102[43];
  assign T101[42] = T3_42_ & T102[42];
  assign T101[41] = T3_41_ & T102[41];
  assign T101[40] = T3_40_ & T102[40];
  assign T101[39] = T3_39_ & T102[39];
  assign T101[38] = T3_38_ & T102[38];
  assign T101[37] = T3_37_ & T102[37];
  assign T101[36] = T3_36_ & T102[36];
  assign T101[35] = T3_35_ & T102[35];
  assign T101[34] = T3_34_ & T102[34];
  assign T101[33] = T3_33_ & T102[33];
  assign T101[32] = T3_32_ & T102[32];
  assign T101[31] = io_resp_bits_data[31] & T102[31];
  assign T101[30] = io_resp_bits_data[30] & T102[30];
  assign T101[29] = io_resp_bits_data[29] & T102[29];
  assign T101[28] = io_resp_bits_data[28] & T102[28];
  assign T101[27] = io_resp_bits_data[27] & T102[27];
  assign T101[26] = io_resp_bits_data[26] & T102[26];
  assign T101[25] = io_resp_bits_data[25] & T102[25];
  assign T101[24] = io_resp_bits_data[24] & T102[24];
  assign T101[23] = io_resp_bits_data[23] & T102[23];
  assign T101[22] = io_resp_bits_data[22] & T102[22];
  assign T101[21] = io_resp_bits_data[21] & T102[21];
  assign T101[20] = io_resp_bits_data[20] & T102[20];
  assign T101[19] = io_resp_bits_data[19] & T102[19];
  assign T101[18] = io_resp_bits_data[18] & T102[18];
  assign T101[17] = io_resp_bits_data[17] & T102[17];
  assign T101[16] = io_resp_bits_data[16] & T102[16];
  assign T101[15] = io_resp_bits_data[15] & T102[15];
  assign T101[14] = io_resp_bits_data[14] & T102[14];
  assign T101[13] = io_resp_bits_data[13] & T102[13];
  assign T101[12] = io_resp_bits_data[12] & T102[12];
  assign T101[11] = io_resp_bits_data[11] & T102[11];
  assign T101[10] = io_resp_bits_data[10] & T102[10];
  assign T101[9] = io_resp_bits_data[9] & T102[9];
  assign T101[8] = io_resp_bits_data[8] & T102[8];
  assign T101[7] = io_resp_bits_data[7] & T102[7];
  assign T101[6] = io_resp_bits_data[6] & T102[6];
  assign T101[5] = io_resp_bits_data[5] & T102[5];
  assign T101[4] = io_resp_bits_data[4] & T102[4];
  assign T101[3] = io_resp_bits_data[3] & T102[3];
  assign T101[2] = io_resp_bits_data[2] & T102[2];
  assign T101[1] = io_resp_bits_data[1] & T102[1];
  assign T101[0] = io_resp_bits_data[0] & T102[0];
  assign T102[63] = ~T103[63];
  assign T102[62] = ~T103[62];
  assign T102[61] = ~T103[61];
  assign T102[60] = ~T103[60];
  assign T102[59] = ~T103[59];
  assign T102[58] = ~T103[58];
  assign T102[57] = ~T103[57];
  assign T102[56] = ~T103[56];
  assign T102[55] = ~T103[55];
  assign T102[54] = ~T103[54];
  assign T102[53] = ~T103[53];
  assign T102[52] = ~T103[52];
  assign T102[51] = ~T103[51];
  assign T102[50] = ~T103[50];
  assign T102[49] = ~T103[49];
  assign T102[48] = ~T103[48];
  assign T102[47] = ~T103[47];
  assign T102[46] = ~T103[46];
  assign T102[45] = ~T103[45];
  assign T102[44] = ~T103[44];
  assign T102[43] = ~T103[43];
  assign T102[42] = ~T103[42];
  assign T102[41] = ~T103[41];
  assign T102[40] = ~T103[40];
  assign T102[39] = ~T103[39];
  assign T102[38] = ~T103[38];
  assign T102[37] = ~T103[37];
  assign T102[36] = ~T103[36];
  assign T102[35] = ~T103[35];
  assign T102[34] = ~T103[34];
  assign T102[33] = ~T103[33];
  assign T102[32] = ~T103[32];
  assign T102[31] = ~T103[31];
  assign T102[30] = ~T103[30];
  assign T102[29] = ~T103[29];
  assign T102[28] = ~T103[28];
  assign T102[27] = ~T103[27];
  assign T102[26] = ~T103[26];
  assign T102[25] = ~T103[25];
  assign T102[24] = ~T103[24];
  assign T102[23] = ~T103[23];
  assign T102[22] = ~T103[22];
  assign T102[21] = ~T103[21];
  assign T102[20] = ~T103[20];
  assign T102[19] = ~T103[19];
  assign T102[18] = ~T103[18];
  assign T102[17] = ~T103[17];
  assign T102[16] = ~T103[16];
  assign T102[15] = ~T103[15];
  assign T102[14] = ~T103[14];
  assign T102[13] = ~T103[13];
  assign T102[12] = ~T103[12];
  assign T102[11] = ~T103[11];
  assign T102[10] = ~T103[10];
  assign T102[9] = ~T103[9];
  assign T102[8] = ~T103[8];
  assign T102[7] = ~T103[7];
  assign T102[6] = ~T103[6];
  assign T102[5] = ~T103[5];
  assign T102[4] = ~T103[4];
  assign T102[3] = ~T103[3];
  assign T102[2] = ~T103[2];
  assign T102[1] = ~T103[1];
  assign T102[0] = ~T103[0];
  assign T111 = T113 & T112;
  assign T112 = ~isHi;
  assign T113 = N804 & N810;
  assign T116[1] = isHi;
  assign T116[2] = N391;
  assign T117[0] = N264;
  assign T118 = T162 & N705;
  assign T120 = T121 | io_kill;
  assign T121 = io_resp_ready & io_resp_valid;
  assign N392 = ~T123;
  assign T122[0] = T123;
  assign T122[1] = N392;
  assign T123 = T450[0] | T124;
  assign T124 = T48[64] & T125;
  assign T125 = ~cmdMul;
  assign N393 = ~T99;
  assign T444[72] = T108[128];
  assign T153 = N708 & isMul;
  assign T447_0 = ~subtractor[64];
  assign N394 = ~subtractor[64];
  assign T162 = N785 & T163;
  assign T163 = ~isMul;
  assign T167 = T162 & T168;
  assign T168 = T171 & T169;
  assign T169 = T170 | T81;
  assign T171 = N798 & subtractor[64];
  assign N395 = ~io_req_bits_dw;
  assign N396 = T167 | T1;
  assign N397 = T162 | N396;
  assign N398 = T153 | N397;
  assign N399 = N682 | N398;
  assign N400 = N674 | N399;
  assign N401 = T11 | N400;
  assign N402 = ~N401;
  assign N535 = T1 | reset;
  assign N536 = T120 | N535;
  assign N537 = T118 | N536;
  assign N538 = T96 | N537;
  assign N539 = N682 | N538;
  assign N540 = N674 | N539;
  assign N541 = N678 | N540;
  assign N542 = ~N541;
  assign N547 = T31 | T1;
  assign N548 = ~N547;
  assign N551 = T45 | T1;
  assign N552 = ~N551;
  assign N619 = T167 | T1;
  assign N620 = T162 | N619;
  assign N621 = T153 | N620;
  assign N622 = ~N621;
  assign N631 = ~T1;
  assign N632 = T167 & N631;
  assign N633 = ~T167;
  assign N634 = N631 & N633;
  assign N635 = T162 & N634;
  assign N636 = ~T162;
  assign N637 = N634 & N636;
  assign N638 = T153 & N637;
  assign N639 = ~T153;
  assign N640 = N637 & N639;
  assign N641 = N682 & N640;
  assign N642 = N640 & N681;
  assign N643 = N674 & N642;
  assign N644 = N642 & N673;
  assign N645 = T11 & N644;
  assign N646 = ~reset;
  assign N647 = T1 & N646;
  assign N648 = N646 & N631;
  assign N649 = T120 & N648;
  assign N650 = ~T120;
  assign N651 = N648 & N650;
  assign N652 = T118 & N651;
  assign N653 = ~T118;
  assign N654 = N651 & N653;
  assign N655 = T96 & N654;
  assign N656 = ~T96;
  assign N657 = N654 & N656;
  assign N658 = N682 & N657;
  assign N659 = N657 & N681;
  assign N660 = N674 & N659;
  assign N661 = N659 & N673;
  assign N662 = N678 & N661;
  assign N663 = T31 & N631;
  assign N664 = T45 & N631;
  assign N665 = T167 & N631;
  assign N666 = N631 & N633;
  assign N667 = T162 & N666;
  assign N668 = N666 & N636;
  assign N669 = T153 & N668;

endmodule