module bp_cce_reg_05
(
  clk_i,
  reset_i,
  decoded_inst_i,
  lce_req_i,
  null_wb_flag_i,
  lce_resp_type_i,
  mem_resp_type_i,
  alu_res_i,
  mov_src_i,
  pending_o_i,
  pending_v_o_i,
  dir_lru_v_i,
  dir_lru_cached_excl_i,
  dir_lru_tag_i,
  dir_tag_i,
  gad_req_addr_way_i,
  gad_transfer_lce_i,
  gad_transfer_lce_way_i,
  gad_transfer_flag_i,
  gad_replacement_flag_i,
  gad_upgrade_flag_i,
  gad_invalidate_flag_i,
  gad_cached_flag_i,
  gad_cached_exclusive_flag_i,
  gad_cached_owned_flag_i,
  gad_cached_dirty_flag_i,
  mshr_o,
  gpr_o,
  coh_state_o,
  nc_data_o
);

  input [211:0] decoded_inst_i;
  input [118:0] lce_req_i;
  input [2:0] lce_resp_type_i;
  input [3:0] mem_resp_type_i;
  input [47:0] alu_res_i;
  input [47:0] mov_src_i;
  input [27:0] dir_lru_tag_i;
  input [27:0] dir_tag_i;
  input [2:0] gad_req_addr_way_i;
  input [2:0] gad_transfer_lce_i;
  input [2:0] gad_transfer_lce_way_i;
  output [121:0] mshr_o;
  output [383:0] gpr_o;
  output [2:0] coh_state_o;
  output [63:0] nc_data_o;
  input clk_i;
  input reset_i;
  input null_wb_flag_i;
  input pending_o_i;
  input pending_v_o_i;
  input dir_lru_v_i;
  input dir_lru_cached_excl_i;
  input gad_transfer_flag_i;
  input gad_replacement_flag_i;
  input gad_upgrade_flag_i;
  input gad_invalidate_flag_i;
  input gad_cached_flag_i;
  input gad_cached_exclusive_flag_i;
  input gad_cached_owned_flag_i;
  input gad_cached_dirty_flag_i;
  wire [121:0] mshr_o;
  wire [383:0] gpr_o,gpr_n;
  wire [2:0] coh_state_o;
  wire [63:0] nc_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,
  uc_req,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,
  N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,
  N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
  N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,
  N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,
  N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,
  N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,
  N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,
  N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,
  N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,
  N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,
  N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,
  N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,
  N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,
  N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,
  N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,
  N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,
  N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,
  N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,
  N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,
  N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,
  N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,
  N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,
  N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,
  N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,
  N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,
  N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,
  N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,
  N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,
  N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,
  N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,
  N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,
  N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,
  N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,
  N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,
  N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,
  N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,
  N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,
  N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,
  N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,
  N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,
  N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,
  N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,
  N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,
  N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,
  N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,
  N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,
  N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,
  N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,
  N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,
  N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,
  N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,
  N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,
  N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,
  N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,
  N1330,N1331,N1332,mshr_n_lce_id__5_,mshr_n_lce_id__4_,mshr_n_lce_id__3_,
  mshr_n_lce_id__2_,mshr_n_lce_id__1_,mshr_n_lce_id__0_,mshr_n_paddr__39_,mshr_n_paddr__38_,
  mshr_n_paddr__37_,mshr_n_paddr__36_,mshr_n_paddr__35_,mshr_n_paddr__34_,
  mshr_n_paddr__33_,mshr_n_paddr__32_,mshr_n_paddr__31_,mshr_n_paddr__30_,
  mshr_n_paddr__29_,mshr_n_paddr__28_,mshr_n_paddr__27_,mshr_n_paddr__26_,mshr_n_paddr__25_,
  mshr_n_paddr__24_,mshr_n_paddr__23_,mshr_n_paddr__22_,mshr_n_paddr__21_,
  mshr_n_paddr__20_,mshr_n_paddr__19_,mshr_n_paddr__18_,mshr_n_paddr__17_,mshr_n_paddr__16_,
  mshr_n_paddr__15_,mshr_n_paddr__14_,mshr_n_paddr__13_,mshr_n_paddr__12_,
  mshr_n_paddr__11_,mshr_n_paddr__10_,mshr_n_paddr__9_,mshr_n_paddr__8_,mshr_n_paddr__7_,
  mshr_n_paddr__6_,mshr_n_paddr__5_,mshr_n_paddr__4_,mshr_n_paddr__3_,mshr_n_paddr__2_,
  mshr_n_paddr__1_,mshr_n_paddr__0_,mshr_n_way_id__2_,mshr_n_way_id__1_,
  mshr_n_way_id__0_,mshr_n_lru_paddr__39_,mshr_n_lru_paddr__38_,mshr_n_lru_paddr__37_,
  mshr_n_lru_paddr__36_,mshr_n_lru_paddr__35_,mshr_n_lru_paddr__34_,
  mshr_n_lru_paddr__33_,mshr_n_lru_paddr__32_,mshr_n_lru_paddr__31_,mshr_n_lru_paddr__30_,
  mshr_n_lru_paddr__29_,mshr_n_lru_paddr__28_,mshr_n_lru_paddr__27_,mshr_n_lru_paddr__26_,
  mshr_n_lru_paddr__25_,mshr_n_lru_paddr__24_,mshr_n_lru_paddr__23_,
  mshr_n_lru_paddr__22_,mshr_n_lru_paddr__21_,mshr_n_lru_paddr__20_,mshr_n_lru_paddr__19_,
  mshr_n_lru_paddr__18_,mshr_n_lru_paddr__17_,mshr_n_lru_paddr__16_,mshr_n_lru_paddr__15_,
  mshr_n_lru_paddr__14_,mshr_n_lru_paddr__13_,mshr_n_lru_paddr__12_,
  mshr_n_lru_paddr__11_,mshr_n_lru_paddr__10_,mshr_n_lru_paddr__9_,mshr_n_lru_paddr__8_,
  mshr_n_lru_paddr__7_,mshr_n_lru_paddr__6_,mshr_n_lru_way_id__2_,mshr_n_lru_way_id__1_,
  mshr_n_lru_way_id__0_,mshr_n_tr_lce_id__2_,mshr_n_tr_lce_id__1_,mshr_n_tr_lce_id__0_,
  mshr_n_tr_way_id__2_,mshr_n_tr_way_id__1_,mshr_n_tr_way_id__0_,
  mshr_n_next_coh_state__2_,mshr_n_next_coh_state__1_,mshr_n_next_coh_state__0_,mshr_n_flags__15_,
  mshr_n_flags__14_,mshr_n_flags__13_,mshr_n_flags__12_,mshr_n_flags__11_,
  mshr_n_flags__10_,mshr_n_flags__9_,mshr_n_flags__8_,mshr_n_flags__7_,mshr_n_flags__6_,
  mshr_n_flags__5_,mshr_n_flags__4_,mshr_n_flags__3_,mshr_n_flags__2_,
  mshr_n_flags__1_,mshr_n_flags__0_,mshr_n_uc_req_size__1_,mshr_n_uc_req_size__0_,N1333,N1334,
  N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,
  N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,
  N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,
  N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,
  N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,
  N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,
  N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,
  N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,
  N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,
  N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,
  N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,
  N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,
  N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,
  N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,
  N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,
  N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,
  N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,
  N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,
  N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,
  N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,
  N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,
  N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,
  N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,
  N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,
  N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,
  N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,
  N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,
  N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,
  N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,
  N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,
  N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,
  N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,
  N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,
  N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,
  N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,
  N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,
  N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,
  N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,
  N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,
  N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,
  N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,
  N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,
  N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,
  N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,
  N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,
  N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,
  N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,
  N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,
  N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,
  N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,
  N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,
  N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,
  N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,
  N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,
  N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,
  N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,
  N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,
  N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,
  N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,
  N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,
  N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,
  N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156;
  reg coh_state_o_2_sv2v_reg,coh_state_o_1_sv2v_reg,coh_state_o_0_sv2v_reg,
  mshr_o_121_sv2v_reg,mshr_o_120_sv2v_reg,mshr_o_119_sv2v_reg,mshr_o_118_sv2v_reg,
  mshr_o_117_sv2v_reg,mshr_o_116_sv2v_reg,mshr_o_115_sv2v_reg,mshr_o_114_sv2v_reg,
  mshr_o_113_sv2v_reg,mshr_o_112_sv2v_reg,mshr_o_111_sv2v_reg,mshr_o_110_sv2v_reg,
  mshr_o_109_sv2v_reg,mshr_o_108_sv2v_reg,mshr_o_107_sv2v_reg,mshr_o_106_sv2v_reg,
  mshr_o_105_sv2v_reg,mshr_o_104_sv2v_reg,mshr_o_103_sv2v_reg,mshr_o_102_sv2v_reg,
  mshr_o_101_sv2v_reg,mshr_o_100_sv2v_reg,mshr_o_99_sv2v_reg,mshr_o_98_sv2v_reg,
  mshr_o_97_sv2v_reg,mshr_o_96_sv2v_reg,mshr_o_95_sv2v_reg,mshr_o_94_sv2v_reg,
  mshr_o_93_sv2v_reg,mshr_o_92_sv2v_reg,mshr_o_91_sv2v_reg,mshr_o_90_sv2v_reg,mshr_o_89_sv2v_reg,
  mshr_o_88_sv2v_reg,mshr_o_87_sv2v_reg,mshr_o_86_sv2v_reg,mshr_o_85_sv2v_reg,
  mshr_o_84_sv2v_reg,mshr_o_83_sv2v_reg,mshr_o_82_sv2v_reg,mshr_o_81_sv2v_reg,
  mshr_o_80_sv2v_reg,mshr_o_79_sv2v_reg,mshr_o_78_sv2v_reg,mshr_o_77_sv2v_reg,
  mshr_o_76_sv2v_reg,mshr_o_75_sv2v_reg,mshr_o_74_sv2v_reg,mshr_o_73_sv2v_reg,
  mshr_o_72_sv2v_reg,mshr_o_71_sv2v_reg,mshr_o_70_sv2v_reg,mshr_o_69_sv2v_reg,mshr_o_68_sv2v_reg,
  mshr_o_67_sv2v_reg,mshr_o_66_sv2v_reg,mshr_o_65_sv2v_reg,mshr_o_64_sv2v_reg,
  mshr_o_63_sv2v_reg,mshr_o_62_sv2v_reg,mshr_o_61_sv2v_reg,mshr_o_60_sv2v_reg,
  mshr_o_59_sv2v_reg,mshr_o_58_sv2v_reg,mshr_o_57_sv2v_reg,mshr_o_56_sv2v_reg,
  mshr_o_55_sv2v_reg,mshr_o_54_sv2v_reg,mshr_o_53_sv2v_reg,mshr_o_52_sv2v_reg,mshr_o_51_sv2v_reg,
  mshr_o_50_sv2v_reg,mshr_o_49_sv2v_reg,mshr_o_48_sv2v_reg,mshr_o_47_sv2v_reg,
  mshr_o_46_sv2v_reg,mshr_o_45_sv2v_reg,mshr_o_44_sv2v_reg,mshr_o_43_sv2v_reg,
  mshr_o_42_sv2v_reg,mshr_o_41_sv2v_reg,mshr_o_40_sv2v_reg,mshr_o_39_sv2v_reg,
  mshr_o_38_sv2v_reg,mshr_o_37_sv2v_reg,mshr_o_36_sv2v_reg,mshr_o_35_sv2v_reg,
  mshr_o_34_sv2v_reg,mshr_o_33_sv2v_reg,mshr_o_32_sv2v_reg,mshr_o_31_sv2v_reg,mshr_o_30_sv2v_reg,
  mshr_o_29_sv2v_reg,mshr_o_28_sv2v_reg,mshr_o_27_sv2v_reg,mshr_o_26_sv2v_reg,
  mshr_o_25_sv2v_reg,mshr_o_24_sv2v_reg,mshr_o_23_sv2v_reg,mshr_o_22_sv2v_reg,
  mshr_o_21_sv2v_reg,mshr_o_20_sv2v_reg,mshr_o_19_sv2v_reg,mshr_o_18_sv2v_reg,
  mshr_o_17_sv2v_reg,mshr_o_16_sv2v_reg,mshr_o_15_sv2v_reg,mshr_o_14_sv2v_reg,
  mshr_o_13_sv2v_reg,mshr_o_12_sv2v_reg,mshr_o_11_sv2v_reg,mshr_o_10_sv2v_reg,mshr_o_9_sv2v_reg,
  mshr_o_8_sv2v_reg,mshr_o_7_sv2v_reg,mshr_o_6_sv2v_reg,mshr_o_5_sv2v_reg,
  mshr_o_4_sv2v_reg,mshr_o_3_sv2v_reg,mshr_o_2_sv2v_reg,mshr_o_1_sv2v_reg,mshr_o_0_sv2v_reg,
  gpr_o_383_sv2v_reg,gpr_o_382_sv2v_reg,gpr_o_381_sv2v_reg,gpr_o_380_sv2v_reg,
  gpr_o_379_sv2v_reg,gpr_o_378_sv2v_reg,gpr_o_377_sv2v_reg,gpr_o_376_sv2v_reg,
  gpr_o_375_sv2v_reg,gpr_o_374_sv2v_reg,gpr_o_373_sv2v_reg,gpr_o_372_sv2v_reg,
  gpr_o_371_sv2v_reg,gpr_o_370_sv2v_reg,gpr_o_369_sv2v_reg,gpr_o_368_sv2v_reg,
  gpr_o_367_sv2v_reg,gpr_o_366_sv2v_reg,gpr_o_365_sv2v_reg,gpr_o_364_sv2v_reg,gpr_o_363_sv2v_reg,
  gpr_o_362_sv2v_reg,gpr_o_361_sv2v_reg,gpr_o_360_sv2v_reg,gpr_o_359_sv2v_reg,
  gpr_o_358_sv2v_reg,gpr_o_357_sv2v_reg,gpr_o_356_sv2v_reg,gpr_o_355_sv2v_reg,
  gpr_o_354_sv2v_reg,gpr_o_353_sv2v_reg,gpr_o_352_sv2v_reg,gpr_o_351_sv2v_reg,
  gpr_o_350_sv2v_reg,gpr_o_349_sv2v_reg,gpr_o_348_sv2v_reg,gpr_o_347_sv2v_reg,
  gpr_o_346_sv2v_reg,gpr_o_345_sv2v_reg,gpr_o_344_sv2v_reg,gpr_o_343_sv2v_reg,gpr_o_342_sv2v_reg,
  gpr_o_341_sv2v_reg,gpr_o_340_sv2v_reg,gpr_o_339_sv2v_reg,gpr_o_338_sv2v_reg,
  gpr_o_337_sv2v_reg,gpr_o_336_sv2v_reg,gpr_o_335_sv2v_reg,gpr_o_334_sv2v_reg,
  gpr_o_333_sv2v_reg,gpr_o_332_sv2v_reg,gpr_o_331_sv2v_reg,gpr_o_330_sv2v_reg,
  gpr_o_329_sv2v_reg,gpr_o_328_sv2v_reg,gpr_o_327_sv2v_reg,gpr_o_326_sv2v_reg,gpr_o_325_sv2v_reg,
  gpr_o_324_sv2v_reg,gpr_o_323_sv2v_reg,gpr_o_322_sv2v_reg,gpr_o_321_sv2v_reg,
  gpr_o_320_sv2v_reg,gpr_o_319_sv2v_reg,gpr_o_318_sv2v_reg,gpr_o_317_sv2v_reg,
  gpr_o_316_sv2v_reg,gpr_o_315_sv2v_reg,gpr_o_314_sv2v_reg,gpr_o_313_sv2v_reg,
  gpr_o_312_sv2v_reg,gpr_o_311_sv2v_reg,gpr_o_310_sv2v_reg,gpr_o_309_sv2v_reg,
  gpr_o_308_sv2v_reg,gpr_o_307_sv2v_reg,gpr_o_306_sv2v_reg,gpr_o_305_sv2v_reg,gpr_o_304_sv2v_reg,
  gpr_o_303_sv2v_reg,gpr_o_302_sv2v_reg,gpr_o_301_sv2v_reg,gpr_o_300_sv2v_reg,
  gpr_o_299_sv2v_reg,gpr_o_298_sv2v_reg,gpr_o_297_sv2v_reg,gpr_o_296_sv2v_reg,
  gpr_o_295_sv2v_reg,gpr_o_294_sv2v_reg,gpr_o_293_sv2v_reg,gpr_o_292_sv2v_reg,
  gpr_o_291_sv2v_reg,gpr_o_290_sv2v_reg,gpr_o_289_sv2v_reg,gpr_o_288_sv2v_reg,
  gpr_o_287_sv2v_reg,gpr_o_286_sv2v_reg,gpr_o_285_sv2v_reg,gpr_o_284_sv2v_reg,gpr_o_283_sv2v_reg,
  gpr_o_282_sv2v_reg,gpr_o_281_sv2v_reg,gpr_o_280_sv2v_reg,gpr_o_279_sv2v_reg,
  gpr_o_278_sv2v_reg,gpr_o_277_sv2v_reg,gpr_o_276_sv2v_reg,gpr_o_275_sv2v_reg,
  gpr_o_274_sv2v_reg,gpr_o_273_sv2v_reg,gpr_o_272_sv2v_reg,gpr_o_271_sv2v_reg,
  gpr_o_270_sv2v_reg,gpr_o_269_sv2v_reg,gpr_o_268_sv2v_reg,gpr_o_267_sv2v_reg,
  gpr_o_266_sv2v_reg,gpr_o_265_sv2v_reg,gpr_o_264_sv2v_reg,gpr_o_263_sv2v_reg,gpr_o_262_sv2v_reg,
  gpr_o_261_sv2v_reg,gpr_o_260_sv2v_reg,gpr_o_259_sv2v_reg,gpr_o_258_sv2v_reg,
  gpr_o_257_sv2v_reg,gpr_o_256_sv2v_reg,gpr_o_255_sv2v_reg,gpr_o_254_sv2v_reg,
  gpr_o_253_sv2v_reg,gpr_o_252_sv2v_reg,gpr_o_251_sv2v_reg,gpr_o_250_sv2v_reg,
  gpr_o_249_sv2v_reg,gpr_o_248_sv2v_reg,gpr_o_247_sv2v_reg,gpr_o_246_sv2v_reg,gpr_o_245_sv2v_reg,
  gpr_o_244_sv2v_reg,gpr_o_243_sv2v_reg,gpr_o_242_sv2v_reg,gpr_o_241_sv2v_reg,
  gpr_o_240_sv2v_reg,gpr_o_239_sv2v_reg,gpr_o_238_sv2v_reg,gpr_o_237_sv2v_reg,
  gpr_o_236_sv2v_reg,gpr_o_235_sv2v_reg,gpr_o_234_sv2v_reg,gpr_o_233_sv2v_reg,
  gpr_o_232_sv2v_reg,gpr_o_231_sv2v_reg,gpr_o_230_sv2v_reg,gpr_o_229_sv2v_reg,
  gpr_o_228_sv2v_reg,gpr_o_227_sv2v_reg,gpr_o_226_sv2v_reg,gpr_o_225_sv2v_reg,gpr_o_224_sv2v_reg,
  gpr_o_223_sv2v_reg,gpr_o_222_sv2v_reg,gpr_o_221_sv2v_reg,gpr_o_220_sv2v_reg,
  gpr_o_219_sv2v_reg,gpr_o_218_sv2v_reg,gpr_o_217_sv2v_reg,gpr_o_216_sv2v_reg,
  gpr_o_215_sv2v_reg,gpr_o_214_sv2v_reg,gpr_o_213_sv2v_reg,gpr_o_212_sv2v_reg,
  gpr_o_211_sv2v_reg,gpr_o_210_sv2v_reg,gpr_o_209_sv2v_reg,gpr_o_208_sv2v_reg,
  gpr_o_207_sv2v_reg,gpr_o_206_sv2v_reg,gpr_o_205_sv2v_reg,gpr_o_204_sv2v_reg,gpr_o_203_sv2v_reg,
  gpr_o_202_sv2v_reg,gpr_o_201_sv2v_reg,gpr_o_200_sv2v_reg,gpr_o_199_sv2v_reg,
  gpr_o_198_sv2v_reg,gpr_o_197_sv2v_reg,gpr_o_196_sv2v_reg,gpr_o_195_sv2v_reg,
  gpr_o_194_sv2v_reg,gpr_o_193_sv2v_reg,gpr_o_192_sv2v_reg,gpr_o_191_sv2v_reg,
  gpr_o_190_sv2v_reg,gpr_o_189_sv2v_reg,gpr_o_188_sv2v_reg,gpr_o_187_sv2v_reg,
  gpr_o_186_sv2v_reg,gpr_o_185_sv2v_reg,gpr_o_184_sv2v_reg,gpr_o_183_sv2v_reg,gpr_o_182_sv2v_reg,
  gpr_o_181_sv2v_reg,gpr_o_180_sv2v_reg,gpr_o_179_sv2v_reg,gpr_o_178_sv2v_reg,
  gpr_o_177_sv2v_reg,gpr_o_176_sv2v_reg,gpr_o_175_sv2v_reg,gpr_o_174_sv2v_reg,
  gpr_o_173_sv2v_reg,gpr_o_172_sv2v_reg,gpr_o_171_sv2v_reg,gpr_o_170_sv2v_reg,
  gpr_o_169_sv2v_reg,gpr_o_168_sv2v_reg,gpr_o_167_sv2v_reg,gpr_o_166_sv2v_reg,gpr_o_165_sv2v_reg,
  gpr_o_164_sv2v_reg,gpr_o_163_sv2v_reg,gpr_o_162_sv2v_reg,gpr_o_161_sv2v_reg,
  gpr_o_160_sv2v_reg,gpr_o_159_sv2v_reg,gpr_o_158_sv2v_reg,gpr_o_157_sv2v_reg,
  gpr_o_156_sv2v_reg,gpr_o_155_sv2v_reg,gpr_o_154_sv2v_reg,gpr_o_153_sv2v_reg,
  gpr_o_152_sv2v_reg,gpr_o_151_sv2v_reg,gpr_o_150_sv2v_reg,gpr_o_149_sv2v_reg,
  gpr_o_148_sv2v_reg,gpr_o_147_sv2v_reg,gpr_o_146_sv2v_reg,gpr_o_145_sv2v_reg,gpr_o_144_sv2v_reg,
  gpr_o_143_sv2v_reg,gpr_o_142_sv2v_reg,gpr_o_141_sv2v_reg,gpr_o_140_sv2v_reg,
  gpr_o_139_sv2v_reg,gpr_o_138_sv2v_reg,gpr_o_137_sv2v_reg,gpr_o_136_sv2v_reg,
  gpr_o_135_sv2v_reg,gpr_o_134_sv2v_reg,gpr_o_133_sv2v_reg,gpr_o_132_sv2v_reg,
  gpr_o_131_sv2v_reg,gpr_o_130_sv2v_reg,gpr_o_129_sv2v_reg,gpr_o_128_sv2v_reg,
  gpr_o_127_sv2v_reg,gpr_o_126_sv2v_reg,gpr_o_125_sv2v_reg,gpr_o_124_sv2v_reg,gpr_o_123_sv2v_reg,
  gpr_o_122_sv2v_reg,gpr_o_121_sv2v_reg,gpr_o_120_sv2v_reg,gpr_o_119_sv2v_reg,
  gpr_o_118_sv2v_reg,gpr_o_117_sv2v_reg,gpr_o_116_sv2v_reg,gpr_o_115_sv2v_reg,
  gpr_o_114_sv2v_reg,gpr_o_113_sv2v_reg,gpr_o_112_sv2v_reg,gpr_o_111_sv2v_reg,
  gpr_o_110_sv2v_reg,gpr_o_109_sv2v_reg,gpr_o_108_sv2v_reg,gpr_o_107_sv2v_reg,
  gpr_o_106_sv2v_reg,gpr_o_105_sv2v_reg,gpr_o_104_sv2v_reg,gpr_o_103_sv2v_reg,gpr_o_102_sv2v_reg,
  gpr_o_101_sv2v_reg,gpr_o_100_sv2v_reg,gpr_o_99_sv2v_reg,gpr_o_98_sv2v_reg,
  gpr_o_97_sv2v_reg,gpr_o_96_sv2v_reg,gpr_o_95_sv2v_reg,gpr_o_94_sv2v_reg,
  gpr_o_93_sv2v_reg,gpr_o_92_sv2v_reg,gpr_o_91_sv2v_reg,gpr_o_90_sv2v_reg,gpr_o_89_sv2v_reg,
  gpr_o_88_sv2v_reg,gpr_o_87_sv2v_reg,gpr_o_86_sv2v_reg,gpr_o_85_sv2v_reg,
  gpr_o_84_sv2v_reg,gpr_o_83_sv2v_reg,gpr_o_82_sv2v_reg,gpr_o_81_sv2v_reg,gpr_o_80_sv2v_reg,
  gpr_o_79_sv2v_reg,gpr_o_78_sv2v_reg,gpr_o_77_sv2v_reg,gpr_o_76_sv2v_reg,
  gpr_o_75_sv2v_reg,gpr_o_74_sv2v_reg,gpr_o_73_sv2v_reg,gpr_o_72_sv2v_reg,gpr_o_71_sv2v_reg,
  gpr_o_70_sv2v_reg,gpr_o_69_sv2v_reg,gpr_o_68_sv2v_reg,gpr_o_67_sv2v_reg,
  gpr_o_66_sv2v_reg,gpr_o_65_sv2v_reg,gpr_o_64_sv2v_reg,gpr_o_63_sv2v_reg,gpr_o_62_sv2v_reg,
  gpr_o_61_sv2v_reg,gpr_o_60_sv2v_reg,gpr_o_59_sv2v_reg,gpr_o_58_sv2v_reg,
  gpr_o_57_sv2v_reg,gpr_o_56_sv2v_reg,gpr_o_55_sv2v_reg,gpr_o_54_sv2v_reg,
  gpr_o_53_sv2v_reg,gpr_o_52_sv2v_reg,gpr_o_51_sv2v_reg,gpr_o_50_sv2v_reg,gpr_o_49_sv2v_reg,
  gpr_o_48_sv2v_reg,gpr_o_47_sv2v_reg,gpr_o_46_sv2v_reg,gpr_o_45_sv2v_reg,
  gpr_o_44_sv2v_reg,gpr_o_43_sv2v_reg,gpr_o_42_sv2v_reg,gpr_o_41_sv2v_reg,gpr_o_40_sv2v_reg,
  gpr_o_39_sv2v_reg,gpr_o_38_sv2v_reg,gpr_o_37_sv2v_reg,gpr_o_36_sv2v_reg,
  gpr_o_35_sv2v_reg,gpr_o_34_sv2v_reg,gpr_o_33_sv2v_reg,gpr_o_32_sv2v_reg,gpr_o_31_sv2v_reg,
  gpr_o_30_sv2v_reg,gpr_o_29_sv2v_reg,gpr_o_28_sv2v_reg,gpr_o_27_sv2v_reg,
  gpr_o_26_sv2v_reg,gpr_o_25_sv2v_reg,gpr_o_24_sv2v_reg,gpr_o_23_sv2v_reg,gpr_o_22_sv2v_reg,
  gpr_o_21_sv2v_reg,gpr_o_20_sv2v_reg,gpr_o_19_sv2v_reg,gpr_o_18_sv2v_reg,
  gpr_o_17_sv2v_reg,gpr_o_16_sv2v_reg,gpr_o_15_sv2v_reg,gpr_o_14_sv2v_reg,
  gpr_o_13_sv2v_reg,gpr_o_12_sv2v_reg,gpr_o_11_sv2v_reg,gpr_o_10_sv2v_reg,gpr_o_9_sv2v_reg,
  gpr_o_8_sv2v_reg,gpr_o_7_sv2v_reg,gpr_o_6_sv2v_reg,gpr_o_5_sv2v_reg,gpr_o_4_sv2v_reg,
  gpr_o_3_sv2v_reg,gpr_o_2_sv2v_reg,gpr_o_1_sv2v_reg,gpr_o_0_sv2v_reg,
  nc_data_o_63_sv2v_reg,nc_data_o_62_sv2v_reg,nc_data_o_61_sv2v_reg,nc_data_o_60_sv2v_reg,
  nc_data_o_59_sv2v_reg,nc_data_o_58_sv2v_reg,nc_data_o_57_sv2v_reg,
  nc_data_o_56_sv2v_reg,nc_data_o_55_sv2v_reg,nc_data_o_54_sv2v_reg,nc_data_o_53_sv2v_reg,
  nc_data_o_52_sv2v_reg,nc_data_o_51_sv2v_reg,nc_data_o_50_sv2v_reg,nc_data_o_49_sv2v_reg,
  nc_data_o_48_sv2v_reg,nc_data_o_47_sv2v_reg,nc_data_o_46_sv2v_reg,
  nc_data_o_45_sv2v_reg,nc_data_o_44_sv2v_reg,nc_data_o_43_sv2v_reg,nc_data_o_42_sv2v_reg,
  nc_data_o_41_sv2v_reg,nc_data_o_40_sv2v_reg,nc_data_o_39_sv2v_reg,nc_data_o_38_sv2v_reg,
  nc_data_o_37_sv2v_reg,nc_data_o_36_sv2v_reg,nc_data_o_35_sv2v_reg,
  nc_data_o_34_sv2v_reg,nc_data_o_33_sv2v_reg,nc_data_o_32_sv2v_reg,nc_data_o_31_sv2v_reg,
  nc_data_o_30_sv2v_reg,nc_data_o_29_sv2v_reg,nc_data_o_28_sv2v_reg,nc_data_o_27_sv2v_reg,
  nc_data_o_26_sv2v_reg,nc_data_o_25_sv2v_reg,nc_data_o_24_sv2v_reg,
  nc_data_o_23_sv2v_reg,nc_data_o_22_sv2v_reg,nc_data_o_21_sv2v_reg,nc_data_o_20_sv2v_reg,
  nc_data_o_19_sv2v_reg,nc_data_o_18_sv2v_reg,nc_data_o_17_sv2v_reg,
  nc_data_o_16_sv2v_reg,nc_data_o_15_sv2v_reg,nc_data_o_14_sv2v_reg,nc_data_o_13_sv2v_reg,
  nc_data_o_12_sv2v_reg,nc_data_o_11_sv2v_reg,nc_data_o_10_sv2v_reg,nc_data_o_9_sv2v_reg,
  nc_data_o_8_sv2v_reg,nc_data_o_7_sv2v_reg,nc_data_o_6_sv2v_reg,nc_data_o_5_sv2v_reg,
  nc_data_o_4_sv2v_reg,nc_data_o_3_sv2v_reg,nc_data_o_2_sv2v_reg,
  nc_data_o_1_sv2v_reg,nc_data_o_0_sv2v_reg;
  assign coh_state_o[2] = coh_state_o_2_sv2v_reg;
  assign coh_state_o[1] = coh_state_o_1_sv2v_reg;
  assign coh_state_o[0] = coh_state_o_0_sv2v_reg;
  assign mshr_o[121] = mshr_o_121_sv2v_reg;
  assign mshr_o[120] = mshr_o_120_sv2v_reg;
  assign mshr_o[119] = mshr_o_119_sv2v_reg;
  assign mshr_o[118] = mshr_o_118_sv2v_reg;
  assign mshr_o[117] = mshr_o_117_sv2v_reg;
  assign mshr_o[116] = mshr_o_116_sv2v_reg;
  assign mshr_o[115] = mshr_o_115_sv2v_reg;
  assign mshr_o[114] = mshr_o_114_sv2v_reg;
  assign mshr_o[113] = mshr_o_113_sv2v_reg;
  assign mshr_o[112] = mshr_o_112_sv2v_reg;
  assign mshr_o[111] = mshr_o_111_sv2v_reg;
  assign mshr_o[110] = mshr_o_110_sv2v_reg;
  assign mshr_o[109] = mshr_o_109_sv2v_reg;
  assign mshr_o[108] = mshr_o_108_sv2v_reg;
  assign mshr_o[107] = mshr_o_107_sv2v_reg;
  assign mshr_o[106] = mshr_o_106_sv2v_reg;
  assign mshr_o[105] = mshr_o_105_sv2v_reg;
  assign mshr_o[104] = mshr_o_104_sv2v_reg;
  assign mshr_o[103] = mshr_o_103_sv2v_reg;
  assign mshr_o[102] = mshr_o_102_sv2v_reg;
  assign mshr_o[101] = mshr_o_101_sv2v_reg;
  assign mshr_o[100] = mshr_o_100_sv2v_reg;
  assign mshr_o[99] = mshr_o_99_sv2v_reg;
  assign mshr_o[98] = mshr_o_98_sv2v_reg;
  assign mshr_o[97] = mshr_o_97_sv2v_reg;
  assign mshr_o[96] = mshr_o_96_sv2v_reg;
  assign mshr_o[95] = mshr_o_95_sv2v_reg;
  assign mshr_o[94] = mshr_o_94_sv2v_reg;
  assign mshr_o[93] = mshr_o_93_sv2v_reg;
  assign mshr_o[92] = mshr_o_92_sv2v_reg;
  assign mshr_o[91] = mshr_o_91_sv2v_reg;
  assign mshr_o[90] = mshr_o_90_sv2v_reg;
  assign mshr_o[89] = mshr_o_89_sv2v_reg;
  assign mshr_o[88] = mshr_o_88_sv2v_reg;
  assign mshr_o[87] = mshr_o_87_sv2v_reg;
  assign mshr_o[86] = mshr_o_86_sv2v_reg;
  assign mshr_o[85] = mshr_o_85_sv2v_reg;
  assign mshr_o[84] = mshr_o_84_sv2v_reg;
  assign mshr_o[83] = mshr_o_83_sv2v_reg;
  assign mshr_o[82] = mshr_o_82_sv2v_reg;
  assign mshr_o[81] = mshr_o_81_sv2v_reg;
  assign mshr_o[80] = mshr_o_80_sv2v_reg;
  assign mshr_o[79] = mshr_o_79_sv2v_reg;
  assign mshr_o[78] = mshr_o_78_sv2v_reg;
  assign mshr_o[77] = mshr_o_77_sv2v_reg;
  assign mshr_o[76] = mshr_o_76_sv2v_reg;
  assign mshr_o[75] = mshr_o_75_sv2v_reg;
  assign mshr_o[74] = mshr_o_74_sv2v_reg;
  assign mshr_o[73] = mshr_o_73_sv2v_reg;
  assign mshr_o[72] = mshr_o_72_sv2v_reg;
  assign mshr_o[71] = mshr_o_71_sv2v_reg;
  assign mshr_o[70] = mshr_o_70_sv2v_reg;
  assign mshr_o[69] = mshr_o_69_sv2v_reg;
  assign mshr_o[68] = mshr_o_68_sv2v_reg;
  assign mshr_o[67] = mshr_o_67_sv2v_reg;
  assign mshr_o[66] = mshr_o_66_sv2v_reg;
  assign mshr_o[65] = mshr_o_65_sv2v_reg;
  assign mshr_o[64] = mshr_o_64_sv2v_reg;
  assign mshr_o[63] = mshr_o_63_sv2v_reg;
  assign mshr_o[62] = mshr_o_62_sv2v_reg;
  assign mshr_o[61] = mshr_o_61_sv2v_reg;
  assign mshr_o[60] = mshr_o_60_sv2v_reg;
  assign mshr_o[59] = mshr_o_59_sv2v_reg;
  assign mshr_o[58] = mshr_o_58_sv2v_reg;
  assign mshr_o[57] = mshr_o_57_sv2v_reg;
  assign mshr_o[56] = mshr_o_56_sv2v_reg;
  assign mshr_o[55] = mshr_o_55_sv2v_reg;
  assign mshr_o[54] = mshr_o_54_sv2v_reg;
  assign mshr_o[53] = mshr_o_53_sv2v_reg;
  assign mshr_o[52] = mshr_o_52_sv2v_reg;
  assign mshr_o[51] = mshr_o_51_sv2v_reg;
  assign mshr_o[50] = mshr_o_50_sv2v_reg;
  assign mshr_o[49] = mshr_o_49_sv2v_reg;
  assign mshr_o[48] = mshr_o_48_sv2v_reg;
  assign mshr_o[47] = mshr_o_47_sv2v_reg;
  assign mshr_o[46] = mshr_o_46_sv2v_reg;
  assign mshr_o[45] = mshr_o_45_sv2v_reg;
  assign mshr_o[44] = mshr_o_44_sv2v_reg;
  assign mshr_o[43] = mshr_o_43_sv2v_reg;
  assign mshr_o[42] = mshr_o_42_sv2v_reg;
  assign mshr_o[41] = mshr_o_41_sv2v_reg;
  assign mshr_o[40] = mshr_o_40_sv2v_reg;
  assign mshr_o[39] = mshr_o_39_sv2v_reg;
  assign mshr_o[38] = mshr_o_38_sv2v_reg;
  assign mshr_o[37] = mshr_o_37_sv2v_reg;
  assign mshr_o[36] = mshr_o_36_sv2v_reg;
  assign mshr_o[35] = mshr_o_35_sv2v_reg;
  assign mshr_o[34] = mshr_o_34_sv2v_reg;
  assign mshr_o[33] = mshr_o_33_sv2v_reg;
  assign mshr_o[32] = mshr_o_32_sv2v_reg;
  assign mshr_o[31] = mshr_o_31_sv2v_reg;
  assign mshr_o[30] = mshr_o_30_sv2v_reg;
  assign mshr_o[29] = mshr_o_29_sv2v_reg;
  assign mshr_o[28] = mshr_o_28_sv2v_reg;
  assign mshr_o[27] = mshr_o_27_sv2v_reg;
  assign mshr_o[26] = mshr_o_26_sv2v_reg;
  assign mshr_o[25] = mshr_o_25_sv2v_reg;
  assign mshr_o[24] = mshr_o_24_sv2v_reg;
  assign mshr_o[23] = mshr_o_23_sv2v_reg;
  assign mshr_o[22] = mshr_o_22_sv2v_reg;
  assign mshr_o[21] = mshr_o_21_sv2v_reg;
  assign mshr_o[20] = mshr_o_20_sv2v_reg;
  assign mshr_o[19] = mshr_o_19_sv2v_reg;
  assign mshr_o[18] = mshr_o_18_sv2v_reg;
  assign mshr_o[17] = mshr_o_17_sv2v_reg;
  assign mshr_o[16] = mshr_o_16_sv2v_reg;
  assign mshr_o[15] = mshr_o_15_sv2v_reg;
  assign mshr_o[14] = mshr_o_14_sv2v_reg;
  assign mshr_o[13] = mshr_o_13_sv2v_reg;
  assign mshr_o[12] = mshr_o_12_sv2v_reg;
  assign mshr_o[11] = mshr_o_11_sv2v_reg;
  assign mshr_o[10] = mshr_o_10_sv2v_reg;
  assign mshr_o[9] = mshr_o_9_sv2v_reg;
  assign mshr_o[8] = mshr_o_8_sv2v_reg;
  assign mshr_o[7] = mshr_o_7_sv2v_reg;
  assign mshr_o[6] = mshr_o_6_sv2v_reg;
  assign mshr_o[5] = mshr_o_5_sv2v_reg;
  assign mshr_o[4] = mshr_o_4_sv2v_reg;
  assign mshr_o[3] = mshr_o_3_sv2v_reg;
  assign mshr_o[2] = mshr_o_2_sv2v_reg;
  assign mshr_o[1] = mshr_o_1_sv2v_reg;
  assign mshr_o[0] = mshr_o_0_sv2v_reg;
  assign gpr_o[383] = gpr_o_383_sv2v_reg;
  assign gpr_o[382] = gpr_o_382_sv2v_reg;
  assign gpr_o[381] = gpr_o_381_sv2v_reg;
  assign gpr_o[380] = gpr_o_380_sv2v_reg;
  assign gpr_o[379] = gpr_o_379_sv2v_reg;
  assign gpr_o[378] = gpr_o_378_sv2v_reg;
  assign gpr_o[377] = gpr_o_377_sv2v_reg;
  assign gpr_o[376] = gpr_o_376_sv2v_reg;
  assign gpr_o[375] = gpr_o_375_sv2v_reg;
  assign gpr_o[374] = gpr_o_374_sv2v_reg;
  assign gpr_o[373] = gpr_o_373_sv2v_reg;
  assign gpr_o[372] = gpr_o_372_sv2v_reg;
  assign gpr_o[371] = gpr_o_371_sv2v_reg;
  assign gpr_o[370] = gpr_o_370_sv2v_reg;
  assign gpr_o[369] = gpr_o_369_sv2v_reg;
  assign gpr_o[368] = gpr_o_368_sv2v_reg;
  assign gpr_o[367] = gpr_o_367_sv2v_reg;
  assign gpr_o[366] = gpr_o_366_sv2v_reg;
  assign gpr_o[365] = gpr_o_365_sv2v_reg;
  assign gpr_o[364] = gpr_o_364_sv2v_reg;
  assign gpr_o[363] = gpr_o_363_sv2v_reg;
  assign gpr_o[362] = gpr_o_362_sv2v_reg;
  assign gpr_o[361] = gpr_o_361_sv2v_reg;
  assign gpr_o[360] = gpr_o_360_sv2v_reg;
  assign gpr_o[359] = gpr_o_359_sv2v_reg;
  assign gpr_o[358] = gpr_o_358_sv2v_reg;
  assign gpr_o[357] = gpr_o_357_sv2v_reg;
  assign gpr_o[356] = gpr_o_356_sv2v_reg;
  assign gpr_o[355] = gpr_o_355_sv2v_reg;
  assign gpr_o[354] = gpr_o_354_sv2v_reg;
  assign gpr_o[353] = gpr_o_353_sv2v_reg;
  assign gpr_o[352] = gpr_o_352_sv2v_reg;
  assign gpr_o[351] = gpr_o_351_sv2v_reg;
  assign gpr_o[350] = gpr_o_350_sv2v_reg;
  assign gpr_o[349] = gpr_o_349_sv2v_reg;
  assign gpr_o[348] = gpr_o_348_sv2v_reg;
  assign gpr_o[347] = gpr_o_347_sv2v_reg;
  assign gpr_o[346] = gpr_o_346_sv2v_reg;
  assign gpr_o[345] = gpr_o_345_sv2v_reg;
  assign gpr_o[344] = gpr_o_344_sv2v_reg;
  assign gpr_o[343] = gpr_o_343_sv2v_reg;
  assign gpr_o[342] = gpr_o_342_sv2v_reg;
  assign gpr_o[341] = gpr_o_341_sv2v_reg;
  assign gpr_o[340] = gpr_o_340_sv2v_reg;
  assign gpr_o[339] = gpr_o_339_sv2v_reg;
  assign gpr_o[338] = gpr_o_338_sv2v_reg;
  assign gpr_o[337] = gpr_o_337_sv2v_reg;
  assign gpr_o[336] = gpr_o_336_sv2v_reg;
  assign gpr_o[335] = gpr_o_335_sv2v_reg;
  assign gpr_o[334] = gpr_o_334_sv2v_reg;
  assign gpr_o[333] = gpr_o_333_sv2v_reg;
  assign gpr_o[332] = gpr_o_332_sv2v_reg;
  assign gpr_o[331] = gpr_o_331_sv2v_reg;
  assign gpr_o[330] = gpr_o_330_sv2v_reg;
  assign gpr_o[329] = gpr_o_329_sv2v_reg;
  assign gpr_o[328] = gpr_o_328_sv2v_reg;
  assign gpr_o[327] = gpr_o_327_sv2v_reg;
  assign gpr_o[326] = gpr_o_326_sv2v_reg;
  assign gpr_o[325] = gpr_o_325_sv2v_reg;
  assign gpr_o[324] = gpr_o_324_sv2v_reg;
  assign gpr_o[323] = gpr_o_323_sv2v_reg;
  assign gpr_o[322] = gpr_o_322_sv2v_reg;
  assign gpr_o[321] = gpr_o_321_sv2v_reg;
  assign gpr_o[320] = gpr_o_320_sv2v_reg;
  assign gpr_o[319] = gpr_o_319_sv2v_reg;
  assign gpr_o[318] = gpr_o_318_sv2v_reg;
  assign gpr_o[317] = gpr_o_317_sv2v_reg;
  assign gpr_o[316] = gpr_o_316_sv2v_reg;
  assign gpr_o[315] = gpr_o_315_sv2v_reg;
  assign gpr_o[314] = gpr_o_314_sv2v_reg;
  assign gpr_o[313] = gpr_o_313_sv2v_reg;
  assign gpr_o[312] = gpr_o_312_sv2v_reg;
  assign gpr_o[311] = gpr_o_311_sv2v_reg;
  assign gpr_o[310] = gpr_o_310_sv2v_reg;
  assign gpr_o[309] = gpr_o_309_sv2v_reg;
  assign gpr_o[308] = gpr_o_308_sv2v_reg;
  assign gpr_o[307] = gpr_o_307_sv2v_reg;
  assign gpr_o[306] = gpr_o_306_sv2v_reg;
  assign gpr_o[305] = gpr_o_305_sv2v_reg;
  assign gpr_o[304] = gpr_o_304_sv2v_reg;
  assign gpr_o[303] = gpr_o_303_sv2v_reg;
  assign gpr_o[302] = gpr_o_302_sv2v_reg;
  assign gpr_o[301] = gpr_o_301_sv2v_reg;
  assign gpr_o[300] = gpr_o_300_sv2v_reg;
  assign gpr_o[299] = gpr_o_299_sv2v_reg;
  assign gpr_o[298] = gpr_o_298_sv2v_reg;
  assign gpr_o[297] = gpr_o_297_sv2v_reg;
  assign gpr_o[296] = gpr_o_296_sv2v_reg;
  assign gpr_o[295] = gpr_o_295_sv2v_reg;
  assign gpr_o[294] = gpr_o_294_sv2v_reg;
  assign gpr_o[293] = gpr_o_293_sv2v_reg;
  assign gpr_o[292] = gpr_o_292_sv2v_reg;
  assign gpr_o[291] = gpr_o_291_sv2v_reg;
  assign gpr_o[290] = gpr_o_290_sv2v_reg;
  assign gpr_o[289] = gpr_o_289_sv2v_reg;
  assign gpr_o[288] = gpr_o_288_sv2v_reg;
  assign gpr_o[287] = gpr_o_287_sv2v_reg;
  assign gpr_o[286] = gpr_o_286_sv2v_reg;
  assign gpr_o[285] = gpr_o_285_sv2v_reg;
  assign gpr_o[284] = gpr_o_284_sv2v_reg;
  assign gpr_o[283] = gpr_o_283_sv2v_reg;
  assign gpr_o[282] = gpr_o_282_sv2v_reg;
  assign gpr_o[281] = gpr_o_281_sv2v_reg;
  assign gpr_o[280] = gpr_o_280_sv2v_reg;
  assign gpr_o[279] = gpr_o_279_sv2v_reg;
  assign gpr_o[278] = gpr_o_278_sv2v_reg;
  assign gpr_o[277] = gpr_o_277_sv2v_reg;
  assign gpr_o[276] = gpr_o_276_sv2v_reg;
  assign gpr_o[275] = gpr_o_275_sv2v_reg;
  assign gpr_o[274] = gpr_o_274_sv2v_reg;
  assign gpr_o[273] = gpr_o_273_sv2v_reg;
  assign gpr_o[272] = gpr_o_272_sv2v_reg;
  assign gpr_o[271] = gpr_o_271_sv2v_reg;
  assign gpr_o[270] = gpr_o_270_sv2v_reg;
  assign gpr_o[269] = gpr_o_269_sv2v_reg;
  assign gpr_o[268] = gpr_o_268_sv2v_reg;
  assign gpr_o[267] = gpr_o_267_sv2v_reg;
  assign gpr_o[266] = gpr_o_266_sv2v_reg;
  assign gpr_o[265] = gpr_o_265_sv2v_reg;
  assign gpr_o[264] = gpr_o_264_sv2v_reg;
  assign gpr_o[263] = gpr_o_263_sv2v_reg;
  assign gpr_o[262] = gpr_o_262_sv2v_reg;
  assign gpr_o[261] = gpr_o_261_sv2v_reg;
  assign gpr_o[260] = gpr_o_260_sv2v_reg;
  assign gpr_o[259] = gpr_o_259_sv2v_reg;
  assign gpr_o[258] = gpr_o_258_sv2v_reg;
  assign gpr_o[257] = gpr_o_257_sv2v_reg;
  assign gpr_o[256] = gpr_o_256_sv2v_reg;
  assign gpr_o[255] = gpr_o_255_sv2v_reg;
  assign gpr_o[254] = gpr_o_254_sv2v_reg;
  assign gpr_o[253] = gpr_o_253_sv2v_reg;
  assign gpr_o[252] = gpr_o_252_sv2v_reg;
  assign gpr_o[251] = gpr_o_251_sv2v_reg;
  assign gpr_o[250] = gpr_o_250_sv2v_reg;
  assign gpr_o[249] = gpr_o_249_sv2v_reg;
  assign gpr_o[248] = gpr_o_248_sv2v_reg;
  assign gpr_o[247] = gpr_o_247_sv2v_reg;
  assign gpr_o[246] = gpr_o_246_sv2v_reg;
  assign gpr_o[245] = gpr_o_245_sv2v_reg;
  assign gpr_o[244] = gpr_o_244_sv2v_reg;
  assign gpr_o[243] = gpr_o_243_sv2v_reg;
  assign gpr_o[242] = gpr_o_242_sv2v_reg;
  assign gpr_o[241] = gpr_o_241_sv2v_reg;
  assign gpr_o[240] = gpr_o_240_sv2v_reg;
  assign gpr_o[239] = gpr_o_239_sv2v_reg;
  assign gpr_o[238] = gpr_o_238_sv2v_reg;
  assign gpr_o[237] = gpr_o_237_sv2v_reg;
  assign gpr_o[236] = gpr_o_236_sv2v_reg;
  assign gpr_o[235] = gpr_o_235_sv2v_reg;
  assign gpr_o[234] = gpr_o_234_sv2v_reg;
  assign gpr_o[233] = gpr_o_233_sv2v_reg;
  assign gpr_o[232] = gpr_o_232_sv2v_reg;
  assign gpr_o[231] = gpr_o_231_sv2v_reg;
  assign gpr_o[230] = gpr_o_230_sv2v_reg;
  assign gpr_o[229] = gpr_o_229_sv2v_reg;
  assign gpr_o[228] = gpr_o_228_sv2v_reg;
  assign gpr_o[227] = gpr_o_227_sv2v_reg;
  assign gpr_o[226] = gpr_o_226_sv2v_reg;
  assign gpr_o[225] = gpr_o_225_sv2v_reg;
  assign gpr_o[224] = gpr_o_224_sv2v_reg;
  assign gpr_o[223] = gpr_o_223_sv2v_reg;
  assign gpr_o[222] = gpr_o_222_sv2v_reg;
  assign gpr_o[221] = gpr_o_221_sv2v_reg;
  assign gpr_o[220] = gpr_o_220_sv2v_reg;
  assign gpr_o[219] = gpr_o_219_sv2v_reg;
  assign gpr_o[218] = gpr_o_218_sv2v_reg;
  assign gpr_o[217] = gpr_o_217_sv2v_reg;
  assign gpr_o[216] = gpr_o_216_sv2v_reg;
  assign gpr_o[215] = gpr_o_215_sv2v_reg;
  assign gpr_o[214] = gpr_o_214_sv2v_reg;
  assign gpr_o[213] = gpr_o_213_sv2v_reg;
  assign gpr_o[212] = gpr_o_212_sv2v_reg;
  assign gpr_o[211] = gpr_o_211_sv2v_reg;
  assign gpr_o[210] = gpr_o_210_sv2v_reg;
  assign gpr_o[209] = gpr_o_209_sv2v_reg;
  assign gpr_o[208] = gpr_o_208_sv2v_reg;
  assign gpr_o[207] = gpr_o_207_sv2v_reg;
  assign gpr_o[206] = gpr_o_206_sv2v_reg;
  assign gpr_o[205] = gpr_o_205_sv2v_reg;
  assign gpr_o[204] = gpr_o_204_sv2v_reg;
  assign gpr_o[203] = gpr_o_203_sv2v_reg;
  assign gpr_o[202] = gpr_o_202_sv2v_reg;
  assign gpr_o[201] = gpr_o_201_sv2v_reg;
  assign gpr_o[200] = gpr_o_200_sv2v_reg;
  assign gpr_o[199] = gpr_o_199_sv2v_reg;
  assign gpr_o[198] = gpr_o_198_sv2v_reg;
  assign gpr_o[197] = gpr_o_197_sv2v_reg;
  assign gpr_o[196] = gpr_o_196_sv2v_reg;
  assign gpr_o[195] = gpr_o_195_sv2v_reg;
  assign gpr_o[194] = gpr_o_194_sv2v_reg;
  assign gpr_o[193] = gpr_o_193_sv2v_reg;
  assign gpr_o[192] = gpr_o_192_sv2v_reg;
  assign gpr_o[191] = gpr_o_191_sv2v_reg;
  assign gpr_o[190] = gpr_o_190_sv2v_reg;
  assign gpr_o[189] = gpr_o_189_sv2v_reg;
  assign gpr_o[188] = gpr_o_188_sv2v_reg;
  assign gpr_o[187] = gpr_o_187_sv2v_reg;
  assign gpr_o[186] = gpr_o_186_sv2v_reg;
  assign gpr_o[185] = gpr_o_185_sv2v_reg;
  assign gpr_o[184] = gpr_o_184_sv2v_reg;
  assign gpr_o[183] = gpr_o_183_sv2v_reg;
  assign gpr_o[182] = gpr_o_182_sv2v_reg;
  assign gpr_o[181] = gpr_o_181_sv2v_reg;
  assign gpr_o[180] = gpr_o_180_sv2v_reg;
  assign gpr_o[179] = gpr_o_179_sv2v_reg;
  assign gpr_o[178] = gpr_o_178_sv2v_reg;
  assign gpr_o[177] = gpr_o_177_sv2v_reg;
  assign gpr_o[176] = gpr_o_176_sv2v_reg;
  assign gpr_o[175] = gpr_o_175_sv2v_reg;
  assign gpr_o[174] = gpr_o_174_sv2v_reg;
  assign gpr_o[173] = gpr_o_173_sv2v_reg;
  assign gpr_o[172] = gpr_o_172_sv2v_reg;
  assign gpr_o[171] = gpr_o_171_sv2v_reg;
  assign gpr_o[170] = gpr_o_170_sv2v_reg;
  assign gpr_o[169] = gpr_o_169_sv2v_reg;
  assign gpr_o[168] = gpr_o_168_sv2v_reg;
  assign gpr_o[167] = gpr_o_167_sv2v_reg;
  assign gpr_o[166] = gpr_o_166_sv2v_reg;
  assign gpr_o[165] = gpr_o_165_sv2v_reg;
  assign gpr_o[164] = gpr_o_164_sv2v_reg;
  assign gpr_o[163] = gpr_o_163_sv2v_reg;
  assign gpr_o[162] = gpr_o_162_sv2v_reg;
  assign gpr_o[161] = gpr_o_161_sv2v_reg;
  assign gpr_o[160] = gpr_o_160_sv2v_reg;
  assign gpr_o[159] = gpr_o_159_sv2v_reg;
  assign gpr_o[158] = gpr_o_158_sv2v_reg;
  assign gpr_o[157] = gpr_o_157_sv2v_reg;
  assign gpr_o[156] = gpr_o_156_sv2v_reg;
  assign gpr_o[155] = gpr_o_155_sv2v_reg;
  assign gpr_o[154] = gpr_o_154_sv2v_reg;
  assign gpr_o[153] = gpr_o_153_sv2v_reg;
  assign gpr_o[152] = gpr_o_152_sv2v_reg;
  assign gpr_o[151] = gpr_o_151_sv2v_reg;
  assign gpr_o[150] = gpr_o_150_sv2v_reg;
  assign gpr_o[149] = gpr_o_149_sv2v_reg;
  assign gpr_o[148] = gpr_o_148_sv2v_reg;
  assign gpr_o[147] = gpr_o_147_sv2v_reg;
  assign gpr_o[146] = gpr_o_146_sv2v_reg;
  assign gpr_o[145] = gpr_o_145_sv2v_reg;
  assign gpr_o[144] = gpr_o_144_sv2v_reg;
  assign gpr_o[143] = gpr_o_143_sv2v_reg;
  assign gpr_o[142] = gpr_o_142_sv2v_reg;
  assign gpr_o[141] = gpr_o_141_sv2v_reg;
  assign gpr_o[140] = gpr_o_140_sv2v_reg;
  assign gpr_o[139] = gpr_o_139_sv2v_reg;
  assign gpr_o[138] = gpr_o_138_sv2v_reg;
  assign gpr_o[137] = gpr_o_137_sv2v_reg;
  assign gpr_o[136] = gpr_o_136_sv2v_reg;
  assign gpr_o[135] = gpr_o_135_sv2v_reg;
  assign gpr_o[134] = gpr_o_134_sv2v_reg;
  assign gpr_o[133] = gpr_o_133_sv2v_reg;
  assign gpr_o[132] = gpr_o_132_sv2v_reg;
  assign gpr_o[131] = gpr_o_131_sv2v_reg;
  assign gpr_o[130] = gpr_o_130_sv2v_reg;
  assign gpr_o[129] = gpr_o_129_sv2v_reg;
  assign gpr_o[128] = gpr_o_128_sv2v_reg;
  assign gpr_o[127] = gpr_o_127_sv2v_reg;
  assign gpr_o[126] = gpr_o_126_sv2v_reg;
  assign gpr_o[125] = gpr_o_125_sv2v_reg;
  assign gpr_o[124] = gpr_o_124_sv2v_reg;
  assign gpr_o[123] = gpr_o_123_sv2v_reg;
  assign gpr_o[122] = gpr_o_122_sv2v_reg;
  assign gpr_o[121] = gpr_o_121_sv2v_reg;
  assign gpr_o[120] = gpr_o_120_sv2v_reg;
  assign gpr_o[119] = gpr_o_119_sv2v_reg;
  assign gpr_o[118] = gpr_o_118_sv2v_reg;
  assign gpr_o[117] = gpr_o_117_sv2v_reg;
  assign gpr_o[116] = gpr_o_116_sv2v_reg;
  assign gpr_o[115] = gpr_o_115_sv2v_reg;
  assign gpr_o[114] = gpr_o_114_sv2v_reg;
  assign gpr_o[113] = gpr_o_113_sv2v_reg;
  assign gpr_o[112] = gpr_o_112_sv2v_reg;
  assign gpr_o[111] = gpr_o_111_sv2v_reg;
  assign gpr_o[110] = gpr_o_110_sv2v_reg;
  assign gpr_o[109] = gpr_o_109_sv2v_reg;
  assign gpr_o[108] = gpr_o_108_sv2v_reg;
  assign gpr_o[107] = gpr_o_107_sv2v_reg;
  assign gpr_o[106] = gpr_o_106_sv2v_reg;
  assign gpr_o[105] = gpr_o_105_sv2v_reg;
  assign gpr_o[104] = gpr_o_104_sv2v_reg;
  assign gpr_o[103] = gpr_o_103_sv2v_reg;
  assign gpr_o[102] = gpr_o_102_sv2v_reg;
  assign gpr_o[101] = gpr_o_101_sv2v_reg;
  assign gpr_o[100] = gpr_o_100_sv2v_reg;
  assign gpr_o[99] = gpr_o_99_sv2v_reg;
  assign gpr_o[98] = gpr_o_98_sv2v_reg;
  assign gpr_o[97] = gpr_o_97_sv2v_reg;
  assign gpr_o[96] = gpr_o_96_sv2v_reg;
  assign gpr_o[95] = gpr_o_95_sv2v_reg;
  assign gpr_o[94] = gpr_o_94_sv2v_reg;
  assign gpr_o[93] = gpr_o_93_sv2v_reg;
  assign gpr_o[92] = gpr_o_92_sv2v_reg;
  assign gpr_o[91] = gpr_o_91_sv2v_reg;
  assign gpr_o[90] = gpr_o_90_sv2v_reg;
  assign gpr_o[89] = gpr_o_89_sv2v_reg;
  assign gpr_o[88] = gpr_o_88_sv2v_reg;
  assign gpr_o[87] = gpr_o_87_sv2v_reg;
  assign gpr_o[86] = gpr_o_86_sv2v_reg;
  assign gpr_o[85] = gpr_o_85_sv2v_reg;
  assign gpr_o[84] = gpr_o_84_sv2v_reg;
  assign gpr_o[83] = gpr_o_83_sv2v_reg;
  assign gpr_o[82] = gpr_o_82_sv2v_reg;
  assign gpr_o[81] = gpr_o_81_sv2v_reg;
  assign gpr_o[80] = gpr_o_80_sv2v_reg;
  assign gpr_o[79] = gpr_o_79_sv2v_reg;
  assign gpr_o[78] = gpr_o_78_sv2v_reg;
  assign gpr_o[77] = gpr_o_77_sv2v_reg;
  assign gpr_o[76] = gpr_o_76_sv2v_reg;
  assign gpr_o[75] = gpr_o_75_sv2v_reg;
  assign gpr_o[74] = gpr_o_74_sv2v_reg;
  assign gpr_o[73] = gpr_o_73_sv2v_reg;
  assign gpr_o[72] = gpr_o_72_sv2v_reg;
  assign gpr_o[71] = gpr_o_71_sv2v_reg;
  assign gpr_o[70] = gpr_o_70_sv2v_reg;
  assign gpr_o[69] = gpr_o_69_sv2v_reg;
  assign gpr_o[68] = gpr_o_68_sv2v_reg;
  assign gpr_o[67] = gpr_o_67_sv2v_reg;
  assign gpr_o[66] = gpr_o_66_sv2v_reg;
  assign gpr_o[65] = gpr_o_65_sv2v_reg;
  assign gpr_o[64] = gpr_o_64_sv2v_reg;
  assign gpr_o[63] = gpr_o_63_sv2v_reg;
  assign gpr_o[62] = gpr_o_62_sv2v_reg;
  assign gpr_o[61] = gpr_o_61_sv2v_reg;
  assign gpr_o[60] = gpr_o_60_sv2v_reg;
  assign gpr_o[59] = gpr_o_59_sv2v_reg;
  assign gpr_o[58] = gpr_o_58_sv2v_reg;
  assign gpr_o[57] = gpr_o_57_sv2v_reg;
  assign gpr_o[56] = gpr_o_56_sv2v_reg;
  assign gpr_o[55] = gpr_o_55_sv2v_reg;
  assign gpr_o[54] = gpr_o_54_sv2v_reg;
  assign gpr_o[53] = gpr_o_53_sv2v_reg;
  assign gpr_o[52] = gpr_o_52_sv2v_reg;
  assign gpr_o[51] = gpr_o_51_sv2v_reg;
  assign gpr_o[50] = gpr_o_50_sv2v_reg;
  assign gpr_o[49] = gpr_o_49_sv2v_reg;
  assign gpr_o[48] = gpr_o_48_sv2v_reg;
  assign gpr_o[47] = gpr_o_47_sv2v_reg;
  assign gpr_o[46] = gpr_o_46_sv2v_reg;
  assign gpr_o[45] = gpr_o_45_sv2v_reg;
  assign gpr_o[44] = gpr_o_44_sv2v_reg;
  assign gpr_o[43] = gpr_o_43_sv2v_reg;
  assign gpr_o[42] = gpr_o_42_sv2v_reg;
  assign gpr_o[41] = gpr_o_41_sv2v_reg;
  assign gpr_o[40] = gpr_o_40_sv2v_reg;
  assign gpr_o[39] = gpr_o_39_sv2v_reg;
  assign gpr_o[38] = gpr_o_38_sv2v_reg;
  assign gpr_o[37] = gpr_o_37_sv2v_reg;
  assign gpr_o[36] = gpr_o_36_sv2v_reg;
  assign gpr_o[35] = gpr_o_35_sv2v_reg;
  assign gpr_o[34] = gpr_o_34_sv2v_reg;
  assign gpr_o[33] = gpr_o_33_sv2v_reg;
  assign gpr_o[32] = gpr_o_32_sv2v_reg;
  assign gpr_o[31] = gpr_o_31_sv2v_reg;
  assign gpr_o[30] = gpr_o_30_sv2v_reg;
  assign gpr_o[29] = gpr_o_29_sv2v_reg;
  assign gpr_o[28] = gpr_o_28_sv2v_reg;
  assign gpr_o[27] = gpr_o_27_sv2v_reg;
  assign gpr_o[26] = gpr_o_26_sv2v_reg;
  assign gpr_o[25] = gpr_o_25_sv2v_reg;
  assign gpr_o[24] = gpr_o_24_sv2v_reg;
  assign gpr_o[23] = gpr_o_23_sv2v_reg;
  assign gpr_o[22] = gpr_o_22_sv2v_reg;
  assign gpr_o[21] = gpr_o_21_sv2v_reg;
  assign gpr_o[20] = gpr_o_20_sv2v_reg;
  assign gpr_o[19] = gpr_o_19_sv2v_reg;
  assign gpr_o[18] = gpr_o_18_sv2v_reg;
  assign gpr_o[17] = gpr_o_17_sv2v_reg;
  assign gpr_o[16] = gpr_o_16_sv2v_reg;
  assign gpr_o[15] = gpr_o_15_sv2v_reg;
  assign gpr_o[14] = gpr_o_14_sv2v_reg;
  assign gpr_o[13] = gpr_o_13_sv2v_reg;
  assign gpr_o[12] = gpr_o_12_sv2v_reg;
  assign gpr_o[11] = gpr_o_11_sv2v_reg;
  assign gpr_o[10] = gpr_o_10_sv2v_reg;
  assign gpr_o[9] = gpr_o_9_sv2v_reg;
  assign gpr_o[8] = gpr_o_8_sv2v_reg;
  assign gpr_o[7] = gpr_o_7_sv2v_reg;
  assign gpr_o[6] = gpr_o_6_sv2v_reg;
  assign gpr_o[5] = gpr_o_5_sv2v_reg;
  assign gpr_o[4] = gpr_o_4_sv2v_reg;
  assign gpr_o[3] = gpr_o_3_sv2v_reg;
  assign gpr_o[2] = gpr_o_2_sv2v_reg;
  assign gpr_o[1] = gpr_o_1_sv2v_reg;
  assign gpr_o[0] = gpr_o_0_sv2v_reg;
  assign nc_data_o[63] = nc_data_o_63_sv2v_reg;
  assign nc_data_o[62] = nc_data_o_62_sv2v_reg;
  assign nc_data_o[61] = nc_data_o_61_sv2v_reg;
  assign nc_data_o[60] = nc_data_o_60_sv2v_reg;
  assign nc_data_o[59] = nc_data_o_59_sv2v_reg;
  assign nc_data_o[58] = nc_data_o_58_sv2v_reg;
  assign nc_data_o[57] = nc_data_o_57_sv2v_reg;
  assign nc_data_o[56] = nc_data_o_56_sv2v_reg;
  assign nc_data_o[55] = nc_data_o_55_sv2v_reg;
  assign nc_data_o[54] = nc_data_o_54_sv2v_reg;
  assign nc_data_o[53] = nc_data_o_53_sv2v_reg;
  assign nc_data_o[52] = nc_data_o_52_sv2v_reg;
  assign nc_data_o[51] = nc_data_o_51_sv2v_reg;
  assign nc_data_o[50] = nc_data_o_50_sv2v_reg;
  assign nc_data_o[49] = nc_data_o_49_sv2v_reg;
  assign nc_data_o[48] = nc_data_o_48_sv2v_reg;
  assign nc_data_o[47] = nc_data_o_47_sv2v_reg;
  assign nc_data_o[46] = nc_data_o_46_sv2v_reg;
  assign nc_data_o[45] = nc_data_o_45_sv2v_reg;
  assign nc_data_o[44] = nc_data_o_44_sv2v_reg;
  assign nc_data_o[43] = nc_data_o_43_sv2v_reg;
  assign nc_data_o[42] = nc_data_o_42_sv2v_reg;
  assign nc_data_o[41] = nc_data_o_41_sv2v_reg;
  assign nc_data_o[40] = nc_data_o_40_sv2v_reg;
  assign nc_data_o[39] = nc_data_o_39_sv2v_reg;
  assign nc_data_o[38] = nc_data_o_38_sv2v_reg;
  assign nc_data_o[37] = nc_data_o_37_sv2v_reg;
  assign nc_data_o[36] = nc_data_o_36_sv2v_reg;
  assign nc_data_o[35] = nc_data_o_35_sv2v_reg;
  assign nc_data_o[34] = nc_data_o_34_sv2v_reg;
  assign nc_data_o[33] = nc_data_o_33_sv2v_reg;
  assign nc_data_o[32] = nc_data_o_32_sv2v_reg;
  assign nc_data_o[31] = nc_data_o_31_sv2v_reg;
  assign nc_data_o[30] = nc_data_o_30_sv2v_reg;
  assign nc_data_o[29] = nc_data_o_29_sv2v_reg;
  assign nc_data_o[28] = nc_data_o_28_sv2v_reg;
  assign nc_data_o[27] = nc_data_o_27_sv2v_reg;
  assign nc_data_o[26] = nc_data_o_26_sv2v_reg;
  assign nc_data_o[25] = nc_data_o_25_sv2v_reg;
  assign nc_data_o[24] = nc_data_o_24_sv2v_reg;
  assign nc_data_o[23] = nc_data_o_23_sv2v_reg;
  assign nc_data_o[22] = nc_data_o_22_sv2v_reg;
  assign nc_data_o[21] = nc_data_o_21_sv2v_reg;
  assign nc_data_o[20] = nc_data_o_20_sv2v_reg;
  assign nc_data_o[19] = nc_data_o_19_sv2v_reg;
  assign nc_data_o[18] = nc_data_o_18_sv2v_reg;
  assign nc_data_o[17] = nc_data_o_17_sv2v_reg;
  assign nc_data_o[16] = nc_data_o_16_sv2v_reg;
  assign nc_data_o[15] = nc_data_o_15_sv2v_reg;
  assign nc_data_o[14] = nc_data_o_14_sv2v_reg;
  assign nc_data_o[13] = nc_data_o_13_sv2v_reg;
  assign nc_data_o[12] = nc_data_o_12_sv2v_reg;
  assign nc_data_o[11] = nc_data_o_11_sv2v_reg;
  assign nc_data_o[10] = nc_data_o_10_sv2v_reg;
  assign nc_data_o[9] = nc_data_o_9_sv2v_reg;
  assign nc_data_o[8] = nc_data_o_8_sv2v_reg;
  assign nc_data_o[7] = nc_data_o_7_sv2v_reg;
  assign nc_data_o[6] = nc_data_o_6_sv2v_reg;
  assign nc_data_o[5] = nc_data_o_5_sv2v_reg;
  assign nc_data_o[4] = nc_data_o_4_sv2v_reg;
  assign nc_data_o[3] = nc_data_o_3_sv2v_reg;
  assign nc_data_o[2] = nc_data_o_2_sv2v_reg;
  assign nc_data_o[1] = nc_data_o_1_sv2v_reg;
  assign nc_data_o[0] = nc_data_o_0_sv2v_reg;
  assign N1438 = N1436 & N1437;
  assign N1439 = decoded_inst_i[125] | N1437;
  assign N1441 = N1436 | decoded_inst_i[124];
  assign N1443 = decoded_inst_i[125] & decoded_inst_i[124];
  assign N1447 = N1445 & N1446;
  assign N1448 = decoded_inst_i[123] | N1446;
  assign N1450 = N1445 | decoded_inst_i[122];
  assign N1452 = decoded_inst_i[123] & decoded_inst_i[122];
  assign N1458 = N1456 & N1457;
  assign N1459 = decoded_inst_i[121] | N1457;
  assign N1461 = N1456 | decoded_inst_i[120];
  assign N1463 = decoded_inst_i[121] & decoded_inst_i[120];
  assign N1467 = N1465 & N1466;
  assign N1468 = decoded_inst_i[119] | N1466;
  assign N1470 = N1465 | decoded_inst_i[118];
  assign N1472 = decoded_inst_i[119] & decoded_inst_i[118];

  always @(posedge clk_i) begin
    if(N2119) begin
      coh_state_o_2_sv2v_reg <= N2122;
    end 
  end


  always @(posedge clk_i) begin
    if(N2119) begin
      coh_state_o_1_sv2v_reg <= N2121;
    end 
  end


  always @(posedge clk_i) begin
    if(N2119) begin
      coh_state_o_0_sv2v_reg <= N2120;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_121_sv2v_reg <= N1661;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_120_sv2v_reg <= N1660;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_119_sv2v_reg <= N1659;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_118_sv2v_reg <= N1658;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_117_sv2v_reg <= N1657;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_116_sv2v_reg <= N1656;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_115_sv2v_reg <= N1655;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_114_sv2v_reg <= N1654;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_113_sv2v_reg <= N1653;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_112_sv2v_reg <= N1652;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_111_sv2v_reg <= N1651;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_110_sv2v_reg <= N1650;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_109_sv2v_reg <= N1649;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_108_sv2v_reg <= N1648;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_107_sv2v_reg <= N1647;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_106_sv2v_reg <= N1646;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_105_sv2v_reg <= N1645;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_104_sv2v_reg <= N1644;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_103_sv2v_reg <= N1643;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_102_sv2v_reg <= N1642;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_101_sv2v_reg <= N1641;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_100_sv2v_reg <= N1640;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_99_sv2v_reg <= N1639;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_98_sv2v_reg <= N1638;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_97_sv2v_reg <= N1637;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_96_sv2v_reg <= N1636;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_95_sv2v_reg <= N1635;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_94_sv2v_reg <= N1634;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_93_sv2v_reg <= N1633;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_92_sv2v_reg <= N1632;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_91_sv2v_reg <= N1631;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_90_sv2v_reg <= N1630;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_89_sv2v_reg <= N1629;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_88_sv2v_reg <= N1628;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_87_sv2v_reg <= N1627;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_86_sv2v_reg <= N1626;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_85_sv2v_reg <= N1625;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_84_sv2v_reg <= N1624;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_83_sv2v_reg <= N1623;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_82_sv2v_reg <= N1622;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_81_sv2v_reg <= N1621;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_80_sv2v_reg <= N1620;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_79_sv2v_reg <= N1619;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_78_sv2v_reg <= N1618;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_77_sv2v_reg <= N1617;
    end 
  end


  always @(posedge clk_i) begin
    if(N1615) begin
      mshr_o_76_sv2v_reg <= N1616;
    end 
  end


  always @(posedge clk_i) begin
    if(N1611) begin
      mshr_o_75_sv2v_reg <= N1614;
    end 
  end


  always @(posedge clk_i) begin
    if(N1611) begin
      mshr_o_74_sv2v_reg <= N1613;
    end 
  end


  always @(posedge clk_i) begin
    if(N1611) begin
      mshr_o_73_sv2v_reg <= N1612;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_72_sv2v_reg <= N1610;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_71_sv2v_reg <= N1609;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_70_sv2v_reg <= N1608;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_69_sv2v_reg <= N1607;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_68_sv2v_reg <= N1606;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_67_sv2v_reg <= N1605;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_66_sv2v_reg <= N1604;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_65_sv2v_reg <= N1603;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_64_sv2v_reg <= N1602;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_63_sv2v_reg <= N1601;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_62_sv2v_reg <= N1600;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_61_sv2v_reg <= N1599;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_60_sv2v_reg <= N1598;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_59_sv2v_reg <= N1597;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_58_sv2v_reg <= N1596;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_57_sv2v_reg <= N1595;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_56_sv2v_reg <= N1594;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_55_sv2v_reg <= N1593;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_54_sv2v_reg <= N1592;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_53_sv2v_reg <= N1591;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_52_sv2v_reg <= N1590;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_51_sv2v_reg <= N1589;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_50_sv2v_reg <= N1588;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_49_sv2v_reg <= N1587;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_48_sv2v_reg <= N1586;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_47_sv2v_reg <= N1585;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_46_sv2v_reg <= N1584;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_45_sv2v_reg <= N1583;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_44_sv2v_reg <= N1582;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_43_sv2v_reg <= N1581;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_42_sv2v_reg <= N1580;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_41_sv2v_reg <= N1579;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_40_sv2v_reg <= N1578;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_39_sv2v_reg <= N1577;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_38_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_37_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_36_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_35_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_34_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1576) begin
      mshr_o_33_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1572) begin
      mshr_o_32_sv2v_reg <= N1575;
    end 
  end


  always @(posedge clk_i) begin
    if(N1572) begin
      mshr_o_31_sv2v_reg <= N1574;
    end 
  end


  always @(posedge clk_i) begin
    if(N1572) begin
      mshr_o_30_sv2v_reg <= N1573;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_29_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_28_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_27_sv2v_reg <= 1'b0;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_26_sv2v_reg <= N1571;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_25_sv2v_reg <= N1570;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_24_sv2v_reg <= N1569;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_23_sv2v_reg <= N1568;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_22_sv2v_reg <= N1567;
    end 
  end


  always @(posedge clk_i) begin
    if(N1565) begin
      mshr_o_21_sv2v_reg <= N1566;
    end 
  end


  always @(posedge clk_i) begin
    if(N1561) begin
      mshr_o_20_sv2v_reg <= N1564;
    end 
  end


  always @(posedge clk_i) begin
    if(N1561) begin
      mshr_o_19_sv2v_reg <= N1563;
    end 
  end


  always @(posedge clk_i) begin
    if(N1561) begin
      mshr_o_18_sv2v_reg <= N1562;
    end 
  end


  always @(posedge clk_i) begin
    if(N1559) begin
      mshr_o_17_sv2v_reg <= N1560;
    end 
  end


  always @(posedge clk_i) begin
    if(N1557) begin
      mshr_o_16_sv2v_reg <= N1558;
    end 
  end


  always @(posedge clk_i) begin
    if(N1555) begin
      mshr_o_15_sv2v_reg <= N1556;
    end 
  end


  always @(posedge clk_i) begin
    if(N1553) begin
      mshr_o_14_sv2v_reg <= N1554;
    end 
  end


  always @(posedge clk_i) begin
    if(N1551) begin
      mshr_o_13_sv2v_reg <= N1552;
    end 
  end


  always @(posedge clk_i) begin
    if(N1549) begin
      mshr_o_12_sv2v_reg <= N1550;
    end 
  end


  always @(posedge clk_i) begin
    if(N1547) begin
      mshr_o_11_sv2v_reg <= N1548;
    end 
  end


  always @(posedge clk_i) begin
    if(N1545) begin
      mshr_o_10_sv2v_reg <= N1546;
    end 
  end


  always @(posedge clk_i) begin
    if(N1543) begin
      mshr_o_9_sv2v_reg <= N1544;
    end 
  end


  always @(posedge clk_i) begin
    if(N1541) begin
      mshr_o_8_sv2v_reg <= N1542;
    end 
  end


  always @(posedge clk_i) begin
    if(N1539) begin
      mshr_o_7_sv2v_reg <= N1540;
    end 
  end


  always @(posedge clk_i) begin
    if(N1537) begin
      mshr_o_6_sv2v_reg <= N1538;
    end 
  end


  always @(posedge clk_i) begin
    if(N1535) begin
      mshr_o_5_sv2v_reg <= N1536;
    end 
  end


  always @(posedge clk_i) begin
    if(N1533) begin
      mshr_o_4_sv2v_reg <= N1534;
    end 
  end


  always @(posedge clk_i) begin
    if(N1531) begin
      mshr_o_3_sv2v_reg <= N1532;
    end 
  end


  always @(posedge clk_i) begin
    if(N1529) begin
      mshr_o_2_sv2v_reg <= N1530;
    end 
  end


  always @(posedge clk_i) begin
    if(N1526) begin
      mshr_o_1_sv2v_reg <= N1528;
    end 
  end


  always @(posedge clk_i) begin
    if(N1526) begin
      mshr_o_0_sv2v_reg <= N1527;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_383_sv2v_reg <= N2053;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_382_sv2v_reg <= N2052;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_381_sv2v_reg <= N2051;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_380_sv2v_reg <= N2050;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_379_sv2v_reg <= N2049;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_378_sv2v_reg <= N2048;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_377_sv2v_reg <= N2047;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_376_sv2v_reg <= N2046;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_375_sv2v_reg <= N2045;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_374_sv2v_reg <= N2044;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_373_sv2v_reg <= N2043;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_372_sv2v_reg <= N2042;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_371_sv2v_reg <= N2041;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_370_sv2v_reg <= N2040;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_369_sv2v_reg <= N2039;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_368_sv2v_reg <= N2038;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_367_sv2v_reg <= N2037;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_366_sv2v_reg <= N2036;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_365_sv2v_reg <= N2035;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_364_sv2v_reg <= N2034;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_363_sv2v_reg <= N2033;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_362_sv2v_reg <= N2032;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_361_sv2v_reg <= N2031;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_360_sv2v_reg <= N2030;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_359_sv2v_reg <= N2029;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_358_sv2v_reg <= N2028;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_357_sv2v_reg <= N2027;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_356_sv2v_reg <= N2026;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_355_sv2v_reg <= N2025;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_354_sv2v_reg <= N2024;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_353_sv2v_reg <= N2023;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_352_sv2v_reg <= N2022;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_351_sv2v_reg <= N2021;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_350_sv2v_reg <= N2020;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_349_sv2v_reg <= N2019;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_348_sv2v_reg <= N2018;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_347_sv2v_reg <= N2017;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_346_sv2v_reg <= N2016;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_345_sv2v_reg <= N2015;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_344_sv2v_reg <= N2014;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_343_sv2v_reg <= N2013;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_342_sv2v_reg <= N2012;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_341_sv2v_reg <= N2011;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_340_sv2v_reg <= N2010;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_339_sv2v_reg <= N2009;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_338_sv2v_reg <= N2008;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_337_sv2v_reg <= N2007;
    end 
  end


  always @(posedge clk_i) begin
    if(N2005) begin
      gpr_o_336_sv2v_reg <= N2006;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_335_sv2v_reg <= N2004;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_334_sv2v_reg <= N2003;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_333_sv2v_reg <= N2002;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_332_sv2v_reg <= N2001;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_331_sv2v_reg <= N2000;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_330_sv2v_reg <= N1999;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_329_sv2v_reg <= N1998;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_328_sv2v_reg <= N1997;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_327_sv2v_reg <= N1996;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_326_sv2v_reg <= N1995;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_325_sv2v_reg <= N1994;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_324_sv2v_reg <= N1993;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_323_sv2v_reg <= N1992;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_322_sv2v_reg <= N1991;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_321_sv2v_reg <= N1990;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_320_sv2v_reg <= N1989;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_319_sv2v_reg <= N1988;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_318_sv2v_reg <= N1987;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_317_sv2v_reg <= N1986;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_316_sv2v_reg <= N1985;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_315_sv2v_reg <= N1984;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_314_sv2v_reg <= N1983;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_313_sv2v_reg <= N1982;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_312_sv2v_reg <= N1981;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_311_sv2v_reg <= N1980;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_310_sv2v_reg <= N1979;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_309_sv2v_reg <= N1978;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_308_sv2v_reg <= N1977;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_307_sv2v_reg <= N1976;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_306_sv2v_reg <= N1975;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_305_sv2v_reg <= N1974;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_304_sv2v_reg <= N1973;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_303_sv2v_reg <= N1972;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_302_sv2v_reg <= N1971;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_301_sv2v_reg <= N1970;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_300_sv2v_reg <= N1969;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_299_sv2v_reg <= N1968;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_298_sv2v_reg <= N1967;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_297_sv2v_reg <= N1966;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_296_sv2v_reg <= N1965;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_295_sv2v_reg <= N1964;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_294_sv2v_reg <= N1963;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_293_sv2v_reg <= N1962;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_292_sv2v_reg <= N1961;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_291_sv2v_reg <= N1960;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_290_sv2v_reg <= N1959;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_289_sv2v_reg <= N1958;
    end 
  end


  always @(posedge clk_i) begin
    if(N1956) begin
      gpr_o_288_sv2v_reg <= N1957;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_287_sv2v_reg <= N1955;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_286_sv2v_reg <= N1954;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_285_sv2v_reg <= N1953;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_284_sv2v_reg <= N1952;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_283_sv2v_reg <= N1951;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_282_sv2v_reg <= N1950;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_281_sv2v_reg <= N1949;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_280_sv2v_reg <= N1948;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_279_sv2v_reg <= N1947;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_278_sv2v_reg <= N1946;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_277_sv2v_reg <= N1945;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_276_sv2v_reg <= N1944;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_275_sv2v_reg <= N1943;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_274_sv2v_reg <= N1942;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_273_sv2v_reg <= N1941;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_272_sv2v_reg <= N1940;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_271_sv2v_reg <= N1939;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_270_sv2v_reg <= N1938;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_269_sv2v_reg <= N1937;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_268_sv2v_reg <= N1936;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_267_sv2v_reg <= N1935;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_266_sv2v_reg <= N1934;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_265_sv2v_reg <= N1933;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_264_sv2v_reg <= N1932;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_263_sv2v_reg <= N1931;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_262_sv2v_reg <= N1930;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_261_sv2v_reg <= N1929;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_260_sv2v_reg <= N1928;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_259_sv2v_reg <= N1927;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_258_sv2v_reg <= N1926;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_257_sv2v_reg <= N1925;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_256_sv2v_reg <= N1924;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_255_sv2v_reg <= N1923;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_254_sv2v_reg <= N1922;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_253_sv2v_reg <= N1921;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_252_sv2v_reg <= N1920;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_251_sv2v_reg <= N1919;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_250_sv2v_reg <= N1918;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_249_sv2v_reg <= N1917;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_248_sv2v_reg <= N1916;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_247_sv2v_reg <= N1915;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_246_sv2v_reg <= N1914;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_245_sv2v_reg <= N1913;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_244_sv2v_reg <= N1912;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_243_sv2v_reg <= N1911;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_242_sv2v_reg <= N1910;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_241_sv2v_reg <= N1909;
    end 
  end


  always @(posedge clk_i) begin
    if(N1907) begin
      gpr_o_240_sv2v_reg <= N1908;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_239_sv2v_reg <= N1906;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_238_sv2v_reg <= N1905;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_237_sv2v_reg <= N1904;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_236_sv2v_reg <= N1903;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_235_sv2v_reg <= N1902;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_234_sv2v_reg <= N1901;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_233_sv2v_reg <= N1900;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_232_sv2v_reg <= N1899;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_231_sv2v_reg <= N1898;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_230_sv2v_reg <= N1897;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_229_sv2v_reg <= N1896;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_228_sv2v_reg <= N1895;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_227_sv2v_reg <= N1894;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_226_sv2v_reg <= N1893;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_225_sv2v_reg <= N1892;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_224_sv2v_reg <= N1891;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_223_sv2v_reg <= N1890;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_222_sv2v_reg <= N1889;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_221_sv2v_reg <= N1888;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_220_sv2v_reg <= N1887;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_219_sv2v_reg <= N1886;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_218_sv2v_reg <= N1885;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_217_sv2v_reg <= N1884;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_216_sv2v_reg <= N1883;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_215_sv2v_reg <= N1882;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_214_sv2v_reg <= N1881;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_213_sv2v_reg <= N1880;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_212_sv2v_reg <= N1879;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_211_sv2v_reg <= N1878;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_210_sv2v_reg <= N1877;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_209_sv2v_reg <= N1876;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_208_sv2v_reg <= N1875;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_207_sv2v_reg <= N1874;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_206_sv2v_reg <= N1873;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_205_sv2v_reg <= N1872;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_204_sv2v_reg <= N1871;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_203_sv2v_reg <= N1870;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_202_sv2v_reg <= N1869;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_201_sv2v_reg <= N1868;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_200_sv2v_reg <= N1867;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_199_sv2v_reg <= N1866;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_198_sv2v_reg <= N1865;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_197_sv2v_reg <= N1864;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_196_sv2v_reg <= N1863;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_195_sv2v_reg <= N1862;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_194_sv2v_reg <= N1861;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_193_sv2v_reg <= N1860;
    end 
  end


  always @(posedge clk_i) begin
    if(N1858) begin
      gpr_o_192_sv2v_reg <= N1859;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_191_sv2v_reg <= N1857;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_190_sv2v_reg <= N1856;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_189_sv2v_reg <= N1855;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_188_sv2v_reg <= N1854;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_187_sv2v_reg <= N1853;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_186_sv2v_reg <= N1852;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_185_sv2v_reg <= N1851;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_184_sv2v_reg <= N1850;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_183_sv2v_reg <= N1849;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_182_sv2v_reg <= N1848;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_181_sv2v_reg <= N1847;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_180_sv2v_reg <= N1846;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_179_sv2v_reg <= N1845;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_178_sv2v_reg <= N1844;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_177_sv2v_reg <= N1843;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_176_sv2v_reg <= N1842;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_175_sv2v_reg <= N1841;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_174_sv2v_reg <= N1840;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_173_sv2v_reg <= N1839;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_172_sv2v_reg <= N1838;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_171_sv2v_reg <= N1837;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_170_sv2v_reg <= N1836;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_169_sv2v_reg <= N1835;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_168_sv2v_reg <= N1834;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_167_sv2v_reg <= N1833;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_166_sv2v_reg <= N1832;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_165_sv2v_reg <= N1831;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_164_sv2v_reg <= N1830;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_163_sv2v_reg <= N1829;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_162_sv2v_reg <= N1828;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_161_sv2v_reg <= N1827;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_160_sv2v_reg <= N1826;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_159_sv2v_reg <= N1825;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_158_sv2v_reg <= N1824;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_157_sv2v_reg <= N1823;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_156_sv2v_reg <= N1822;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_155_sv2v_reg <= N1821;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_154_sv2v_reg <= N1820;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_153_sv2v_reg <= N1819;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_152_sv2v_reg <= N1818;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_151_sv2v_reg <= N1817;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_150_sv2v_reg <= N1816;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_149_sv2v_reg <= N1815;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_148_sv2v_reg <= N1814;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_147_sv2v_reg <= N1813;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_146_sv2v_reg <= N1812;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_145_sv2v_reg <= N1811;
    end 
  end


  always @(posedge clk_i) begin
    if(N1809) begin
      gpr_o_144_sv2v_reg <= N1810;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_143_sv2v_reg <= N1808;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_142_sv2v_reg <= N1807;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_141_sv2v_reg <= N1806;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_140_sv2v_reg <= N1805;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_139_sv2v_reg <= N1804;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_138_sv2v_reg <= N1803;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_137_sv2v_reg <= N1802;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_136_sv2v_reg <= N1801;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_135_sv2v_reg <= N1800;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_134_sv2v_reg <= N1799;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_133_sv2v_reg <= N1798;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_132_sv2v_reg <= N1797;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_131_sv2v_reg <= N1796;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_130_sv2v_reg <= N1795;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_129_sv2v_reg <= N1794;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_128_sv2v_reg <= N1793;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_127_sv2v_reg <= N1792;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_126_sv2v_reg <= N1791;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_125_sv2v_reg <= N1790;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_124_sv2v_reg <= N1789;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_123_sv2v_reg <= N1788;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_122_sv2v_reg <= N1787;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_121_sv2v_reg <= N1786;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_120_sv2v_reg <= N1785;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_119_sv2v_reg <= N1784;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_118_sv2v_reg <= N1783;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_117_sv2v_reg <= N1782;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_116_sv2v_reg <= N1781;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_115_sv2v_reg <= N1780;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_114_sv2v_reg <= N1779;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_113_sv2v_reg <= N1778;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_112_sv2v_reg <= N1777;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_111_sv2v_reg <= N1776;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_110_sv2v_reg <= N1775;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_109_sv2v_reg <= N1774;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_108_sv2v_reg <= N1773;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_107_sv2v_reg <= N1772;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_106_sv2v_reg <= N1771;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_105_sv2v_reg <= N1770;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_104_sv2v_reg <= N1769;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_103_sv2v_reg <= N1768;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_102_sv2v_reg <= N1767;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_101_sv2v_reg <= N1766;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_100_sv2v_reg <= N1765;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_99_sv2v_reg <= N1764;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_98_sv2v_reg <= N1763;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_97_sv2v_reg <= N1762;
    end 
  end


  always @(posedge clk_i) begin
    if(N1760) begin
      gpr_o_96_sv2v_reg <= N1761;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_95_sv2v_reg <= N1759;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_94_sv2v_reg <= N1758;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_93_sv2v_reg <= N1757;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_92_sv2v_reg <= N1756;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_91_sv2v_reg <= N1755;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_90_sv2v_reg <= N1754;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_89_sv2v_reg <= N1753;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_88_sv2v_reg <= N1752;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_87_sv2v_reg <= N1751;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_86_sv2v_reg <= N1750;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_85_sv2v_reg <= N1749;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_84_sv2v_reg <= N1748;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_83_sv2v_reg <= N1747;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_82_sv2v_reg <= N1746;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_81_sv2v_reg <= N1745;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_80_sv2v_reg <= N1744;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_79_sv2v_reg <= N1743;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_78_sv2v_reg <= N1742;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_77_sv2v_reg <= N1741;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_76_sv2v_reg <= N1740;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_75_sv2v_reg <= N1739;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_74_sv2v_reg <= N1738;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_73_sv2v_reg <= N1737;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_72_sv2v_reg <= N1736;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_71_sv2v_reg <= N1735;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_70_sv2v_reg <= N1734;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_69_sv2v_reg <= N1733;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_68_sv2v_reg <= N1732;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_67_sv2v_reg <= N1731;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_66_sv2v_reg <= N1730;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_65_sv2v_reg <= N1729;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_64_sv2v_reg <= N1728;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_63_sv2v_reg <= N1727;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_62_sv2v_reg <= N1726;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_61_sv2v_reg <= N1725;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_60_sv2v_reg <= N1724;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_59_sv2v_reg <= N1723;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_58_sv2v_reg <= N1722;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_57_sv2v_reg <= N1721;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_56_sv2v_reg <= N1720;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_55_sv2v_reg <= N1719;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_54_sv2v_reg <= N1718;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_53_sv2v_reg <= N1717;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_52_sv2v_reg <= N1716;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_51_sv2v_reg <= N1715;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_50_sv2v_reg <= N1714;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_49_sv2v_reg <= N1713;
    end 
  end


  always @(posedge clk_i) begin
    if(N1711) begin
      gpr_o_48_sv2v_reg <= N1712;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_47_sv2v_reg <= N1710;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_46_sv2v_reg <= N1709;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_45_sv2v_reg <= N1708;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_44_sv2v_reg <= N1707;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_43_sv2v_reg <= N1706;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_42_sv2v_reg <= N1705;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_41_sv2v_reg <= N1704;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_40_sv2v_reg <= N1703;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_39_sv2v_reg <= N1702;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_38_sv2v_reg <= N1701;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_37_sv2v_reg <= N1700;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_36_sv2v_reg <= N1699;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_35_sv2v_reg <= N1698;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_34_sv2v_reg <= N1697;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_33_sv2v_reg <= N1696;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_32_sv2v_reg <= N1695;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_31_sv2v_reg <= N1694;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_30_sv2v_reg <= N1693;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_29_sv2v_reg <= N1692;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_28_sv2v_reg <= N1691;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_27_sv2v_reg <= N1690;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_26_sv2v_reg <= N1689;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_25_sv2v_reg <= N1688;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_24_sv2v_reg <= N1687;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_23_sv2v_reg <= N1686;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_22_sv2v_reg <= N1685;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_21_sv2v_reg <= N1684;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_20_sv2v_reg <= N1683;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_19_sv2v_reg <= N1682;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_18_sv2v_reg <= N1681;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_17_sv2v_reg <= N1680;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_16_sv2v_reg <= N1679;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_15_sv2v_reg <= N1678;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_14_sv2v_reg <= N1677;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_13_sv2v_reg <= N1676;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_12_sv2v_reg <= N1675;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_11_sv2v_reg <= N1674;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_10_sv2v_reg <= N1673;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_9_sv2v_reg <= N1672;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_8_sv2v_reg <= N1671;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_7_sv2v_reg <= N1670;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_6_sv2v_reg <= N1669;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_5_sv2v_reg <= N1668;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_4_sv2v_reg <= N1667;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_3_sv2v_reg <= N1666;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_2_sv2v_reg <= N1665;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_1_sv2v_reg <= N1664;
    end 
  end


  always @(posedge clk_i) begin
    if(N1662) begin
      gpr_o_0_sv2v_reg <= N1663;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_63_sv2v_reg <= N2118;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_62_sv2v_reg <= N2117;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_61_sv2v_reg <= N2116;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_60_sv2v_reg <= N2115;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_59_sv2v_reg <= N2114;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_58_sv2v_reg <= N2113;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_57_sv2v_reg <= N2112;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_56_sv2v_reg <= N2111;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_55_sv2v_reg <= N2110;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_54_sv2v_reg <= N2109;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_53_sv2v_reg <= N2108;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_52_sv2v_reg <= N2107;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_51_sv2v_reg <= N2106;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_50_sv2v_reg <= N2105;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_49_sv2v_reg <= N2104;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_48_sv2v_reg <= N2103;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_47_sv2v_reg <= N2102;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_46_sv2v_reg <= N2101;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_45_sv2v_reg <= N2100;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_44_sv2v_reg <= N2099;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_43_sv2v_reg <= N2098;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_42_sv2v_reg <= N2097;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_41_sv2v_reg <= N2096;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_40_sv2v_reg <= N2095;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_39_sv2v_reg <= N2094;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_38_sv2v_reg <= N2093;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_37_sv2v_reg <= N2092;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_36_sv2v_reg <= N2091;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_35_sv2v_reg <= N2090;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_34_sv2v_reg <= N2089;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_33_sv2v_reg <= N2088;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_32_sv2v_reg <= N2087;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_31_sv2v_reg <= N2086;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_30_sv2v_reg <= N2085;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_29_sv2v_reg <= N2084;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_28_sv2v_reg <= N2083;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_27_sv2v_reg <= N2082;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_26_sv2v_reg <= N2081;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_25_sv2v_reg <= N2080;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_24_sv2v_reg <= N2079;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_23_sv2v_reg <= N2078;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_22_sv2v_reg <= N2077;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_21_sv2v_reg <= N2076;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_20_sv2v_reg <= N2075;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_19_sv2v_reg <= N2074;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_18_sv2v_reg <= N2073;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_17_sv2v_reg <= N2072;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_16_sv2v_reg <= N2071;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_15_sv2v_reg <= N2070;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_14_sv2v_reg <= N2069;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_13_sv2v_reg <= N2068;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_12_sv2v_reg <= N2067;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_11_sv2v_reg <= N2066;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_10_sv2v_reg <= N2065;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_9_sv2v_reg <= N2064;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_8_sv2v_reg <= N2063;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_7_sv2v_reg <= N2062;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_6_sv2v_reg <= N2061;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_5_sv2v_reg <= N2060;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_4_sv2v_reg <= N2059;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_3_sv2v_reg <= N2058;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_2_sv2v_reg <= N2057;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_1_sv2v_reg <= N2056;
    end 
  end


  always @(posedge clk_i) begin
    if(N2054) begin
      nc_data_o_0_sv2v_reg <= N2055;
    end 
  end

  assign N2123 = ~decoded_inst_i[188];
  assign N2124 = decoded_inst_i[187] | N2123;
  assign N2125 = ~N2124;
  assign N2126 = ~decoded_inst_i[200];
  assign N2127 = decoded_inst_i[202] | decoded_inst_i[203];
  assign N2128 = decoded_inst_i[201] | N2127;
  assign N2129 = N2126 | N2128;
  assign N2130 = decoded_inst_i[199] | N2129;
  assign N2131 = ~N2130;
  assign N2132 = decoded_inst_i[200] | N2128;
  assign N2133 = decoded_inst_i[199] | N2132;
  assign N2134 = ~N2133;
  assign N2135 = ~lce_req_i[11];
  assign N2136 = N2135 | lce_req_i[12];
  assign N2137 = lce_req_i[10] | N2136;
  assign N2138 = ~N2137;
  assign N2139 = ~lce_req_i[10];
  assign N2140 = N2139 | N2136;
  assign N2141 = ~N2140;
  assign N2142 = ~decoded_inst_i[205];
  assign N2143 = decoded_inst_i[206] | decoded_inst_i[207];
  assign N2144 = N2142 | N2143;
  assign N2145 = decoded_inst_i[204] | N2144;
  assign N2146 = ~N2145;
  assign { N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143 } = (N0)? dir_tag_i : 
                                                                                                                                                                                      (N1)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N0 = N141;
  assign N1 = N142;
  assign { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } = (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N3)? { N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N139;
  assign N3 = N140;
  assign { N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203 } = (N4)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N5)? { N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171 } : 1'b0;
  assign N4 = N137;
  assign N5 = N138;
  assign { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235 } = (N6)? mov_src_i : 
                                                                                                                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N206, N205, N204, N203 } : 1'b0;
  assign N6 = N135;
  assign N7 = N136;
  assign gpr_n[47:0] = (N8)? alu_res_i : 
                       (N9)? { N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235 } : 1'b0;
  assign N8 = N133;
  assign N9 = N134;
  assign { N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293 } = (N10)? dir_tag_i : 
                                                                                                                                                                                      (N11)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N10 = N291;
  assign N11 = N292;
  assign { N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321 } = (N12)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N13)? { N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N12 = N289;
  assign N13 = N290;
  assign { N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353 } = (N14)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N15)? { N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321 } : 1'b0;
  assign N14 = N287;
  assign N15 = N288;
  assign { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385 } = (N16)? mov_src_i : 
                                                                                                                                                                                                                                                                                                              (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N356, N355, N354, N353 } : 1'b0;
  assign N16 = N285;
  assign N17 = N286;
  assign gpr_n[95:48] = (N18)? alu_res_i : 
                        (N19)? { N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385 } : 1'b0;
  assign N18 = N283;
  assign N19 = N284;
  assign { N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443 } = (N20)? dir_tag_i : 
                                                                                                                                                                                      (N21)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N20 = N441;
  assign N21 = N442;
  assign { N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471 } = (N22)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N23)? { N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = N439;
  assign N23 = N440;
  assign { N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503 } = (N24)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N25)? { N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471 } : 1'b0;
  assign N24 = N437;
  assign N25 = N438;
  assign { N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } = (N26)? mov_src_i : 
                                                                                                                                                                                                                                                                                                              (N27)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N506, N505, N504, N503 } : 1'b0;
  assign N26 = N435;
  assign N27 = N436;
  assign gpr_n[143:96] = (N28)? alu_res_i : 
                         (N29)? { N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535 } : 1'b0;
  assign N28 = N433;
  assign N29 = N434;
  assign { N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593 } = (N30)? dir_tag_i : 
                                                                                                                                                                                      (N31)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N30 = N591;
  assign N31 = N592;
  assign { N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621 } = (N32)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N33)? { N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N32 = N589;
  assign N33 = N590;
  assign { N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653 } = (N34)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N35)? { N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621 } : 1'b0;
  assign N34 = N587;
  assign N35 = N588;
  assign { N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685 } = (N36)? mov_src_i : 
                                                                                                                                                                                                                                                                                                              (N37)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N656, N655, N654, N653 } : 1'b0;
  assign N36 = N585;
  assign N37 = N586;
  assign gpr_n[191:144] = (N38)? alu_res_i : 
                          (N39)? { N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685 } : 1'b0;
  assign N38 = N583;
  assign N39 = N584;
  assign { N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743 } = (N40)? dir_tag_i : 
                                                                                                                                                                                      (N41)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N40 = N741;
  assign N41 = N742;
  assign { N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771 } = (N42)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N43)? { N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N42 = N739;
  assign N43 = N740;
  assign { N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803 } = (N44)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N45)? { N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771 } : 1'b0;
  assign N44 = N737;
  assign N45 = N738;
  assign { N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835 } = (N46)? mov_src_i : 
                                                                                                                                                                                                                                                                                                              (N47)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N806, N805, N804, N803 } : 1'b0;
  assign N46 = N735;
  assign N47 = N736;
  assign gpr_n[239:192] = (N48)? alu_res_i : 
                          (N49)? { N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835 } : 1'b0;
  assign N48 = N733;
  assign N49 = N734;
  assign { N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893 } = (N50)? dir_tag_i : 
                                                                                                                                                                                      (N51)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N50 = N891;
  assign N51 = N892;
  assign { N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921 } = (N52)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                              (N53)? { N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N52 = N889;
  assign N53 = N890;
  assign { N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953 } = (N54)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                              (N55)? { N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921 } : 1'b0;
  assign N54 = N887;
  assign N55 = N888;
  assign { N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985 } = (N56)? mov_src_i : 
                                                                                                                                                                                                                                                                                                                                               (N57)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N956, N955, N954, N953 } : 1'b0;
  assign N56 = N885;
  assign N57 = N886;
  assign gpr_n[287:240] = (N58)? alu_res_i : 
                          (N59)? { N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985 } : 1'b0;
  assign N58 = N883;
  assign N59 = N884;
  assign { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043 } = (N60)? dir_tag_i : 
                                                                                                                                                                                                                  (N61)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N60 = N1041;
  assign N61 = N1042;
  assign { N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071 } = (N62)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                                                              (N63)? { N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N62 = N1039;
  assign N63 = N1040;
  assign { N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103 } = (N64)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                                                              (N65)? { N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071 } : 1'b0;
  assign N64 = N1037;
  assign N65 = N1038;
  assign { N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135 } = (N66)? mov_src_i : 
                                                                                                                                                                                                                                                                                                                                                              (N67)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1106, N1105, N1104, N1103 } : 1'b0;
  assign N66 = N1035;
  assign N67 = N1036;
  assign gpr_n[335:288] = (N68)? alu_res_i : 
                          (N69)? { N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135 } : 1'b0;
  assign N68 = N1033;
  assign N69 = N1034;
  assign { N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193 } = (N70)? dir_tag_i : 
                                                                                                                                                                                                                  (N71)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N70 = N1191;
  assign N71 = N1192;
  assign { N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221 } = (N72)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mem_resp_type_i } : 
                                                                                                                                                                                                                                              (N73)? { N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N72 = N1189;
  assign N73 = N1190;
  assign { N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253 } = (N74)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, lce_resp_type_i } : 
                                                                                                                                                                                                                                              (N75)? { N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221 } : 1'b0;
  assign N74 = N1187;
  assign N75 = N1188;
  assign { N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285 } = (N76)? mov_src_i : 
                                                                                                                                                                                                                                                                                                                                                              (N77)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N1256, N1255, N1254, N1253 } : 1'b0;
  assign N76 = N1185;
  assign N77 = N1186;
  assign gpr_n[383:336] = (N78)? alu_res_i : 
                          (N79)? { N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285 } : 1'b0;
  assign N78 = N1183;
  assign N79 = N1184;
  assign { N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336 } = (N80)? { lce_req_i[9:4], lce_req_i[52:13] } : 
                                                                                                                                                                                                                                                                                                                                                (N81)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N80 = N1335;
  assign N81 = decoded_inst_i[128];
  assign { N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382 } = (N82)? { N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336 } : 
                                                                                                                                                                                                                                                                                                                                                (N83)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N82 = N1334;
  assign N83 = decoded_inst_i[129];
  assign { N1432, N1431, N1430 } = (N84)? lce_req_i[56:54] : 
                                   (N85)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N84 = N1429;
  assign N85 = decoded_inst_i[126];
  assign { N1435, N1434, N1433 } = (N86)? { N1432, N1431, N1430 } : 
                                   (N87)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N86 = N1428;
  assign N87 = decoded_inst_i[127];
  assign N1444 = (N88)? lce_req_i[10] : 
                 (N89)? 1'b0 : 
                 (N90)? decoded_inst_i[135] : 
                 (N91)? 1'b0 : 1'b0;
  assign N88 = N1438;
  assign N89 = N1440;
  assign N90 = N1442;
  assign N91 = N1443;
  assign { N1455, N1454, N1453 } = (N92)? { uc_req, lce_req_i[54:53] } : 
                                   (N93)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N94)? { decoded_inst_i[135:135], 1'b0, 1'b0 } : 
                                   (N95)? { 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N92 = N1447;
  assign N93 = N1449;
  assign N94 = N1451;
  assign N95 = N1452;
  assign N1464 = (N96)? lce_req_i[53] : 
                 (N97)? 1'b0 : 
                 (N98)? decoded_inst_i[135] : 
                 (N99)? 1'b0 : 1'b0;
  assign N96 = N1458;
  assign N97 = N1460;
  assign N98 = N1462;
  assign N99 = N1463;
  assign N1473 = (N100)? lce_req_i[57] : 
                 (N101)? 1'b0 : 
                 (N102)? decoded_inst_i[135] : 
                 (N103)? 1'b0 : 1'b0;
  assign N100 = N1467;
  assign N101 = N1469;
  assign N102 = N1471;
  assign N103 = N1472;
  assign N1475 = (N104)? null_wb_flag_i : 
                 (N105)? decoded_inst_i[135] : 1'b0;
  assign N104 = N1474;
  assign N105 = decoded_inst_i[107];
  assign N1477 = (N106)? gad_transfer_flag_i : 
                 (N107)? decoded_inst_i[135] : 1'b0;
  assign N106 = N1476;
  assign N107 = decoded_inst_i[111];
  assign N1479 = (N108)? pending_o_i : 
                 (N109)? decoded_inst_i[135] : 1'b0;
  assign N108 = N1478;
  assign N109 = decoded_inst_i[117];
  assign N1481 = (N110)? gad_replacement_flag_i : 
                 (N111)? decoded_inst_i[135] : 1'b0;
  assign N110 = N1480;
  assign N111 = decoded_inst_i[110];
  assign N1483 = (N112)? gad_upgrade_flag_i : 
                 (N113)? decoded_inst_i[135] : 1'b0;
  assign N112 = N1482;
  assign N113 = decoded_inst_i[109];
  assign N1485 = (N114)? gad_invalidate_flag_i : 
                 (N115)? decoded_inst_i[135] : 1'b0;
  assign N114 = N1484;
  assign N115 = decoded_inst_i[108];
  assign N1487 = (N116)? gad_cached_flag_i : 
                 (N117)? decoded_inst_i[135] : 1'b0;
  assign N116 = N1486;
  assign N117 = decoded_inst_i[115];
  assign N1489 = (N118)? gad_cached_exclusive_flag_i : 
                 (N119)? decoded_inst_i[135] : 1'b0;
  assign N118 = N1488;
  assign N119 = decoded_inst_i[114];
  assign N1491 = (N120)? gad_cached_owned_flag_i : 
                 (N121)? decoded_inst_i[135] : 1'b0;
  assign N120 = N1490;
  assign N121 = decoded_inst_i[113];
  assign N1493 = (N122)? gad_cached_dirty_flag_i : 
                 (N123)? decoded_inst_i[135] : 1'b0;
  assign N122 = N1492;
  assign N123 = decoded_inst_i[112];
  assign N1495 = (N124)? dir_lru_cached_excl_i : 
                 (N125)? decoded_inst_i[135] : 1'b0;
  assign N124 = N1494;
  assign N125 = decoded_inst_i[116];
  assign N1497 = (N126)? decoded_inst_i[5] : 
                 (N127)? decoded_inst_i[135] : 1'b0;
  assign N126 = N1496;
  assign N127 = decoded_inst_i[106];
  assign { mshr_n_lce_id__5_, mshr_n_lce_id__4_, mshr_n_lce_id__3_, mshr_n_lce_id__2_, mshr_n_lce_id__1_, mshr_n_lce_id__0_, mshr_n_paddr__39_, mshr_n_paddr__38_, mshr_n_paddr__37_, mshr_n_paddr__36_, mshr_n_paddr__35_, mshr_n_paddr__34_, mshr_n_paddr__33_, mshr_n_paddr__32_, mshr_n_paddr__31_, mshr_n_paddr__30_, mshr_n_paddr__29_, mshr_n_paddr__28_, mshr_n_paddr__27_, mshr_n_paddr__26_, mshr_n_paddr__25_, mshr_n_paddr__24_, mshr_n_paddr__23_, mshr_n_paddr__22_, mshr_n_paddr__21_, mshr_n_paddr__20_, mshr_n_paddr__19_, mshr_n_paddr__18_, mshr_n_paddr__17_, mshr_n_paddr__16_, mshr_n_paddr__15_, mshr_n_paddr__14_, mshr_n_paddr__13_, mshr_n_paddr__12_, mshr_n_paddr__11_, mshr_n_paddr__10_, mshr_n_paddr__9_, mshr_n_paddr__8_, mshr_n_paddr__7_, mshr_n_paddr__6_, mshr_n_paddr__5_, mshr_n_paddr__4_, mshr_n_paddr__3_, mshr_n_paddr__2_, mshr_n_paddr__1_, mshr_n_paddr__0_, mshr_n_way_id__2_, mshr_n_way_id__1_, mshr_n_way_id__0_, mshr_n_lru_paddr__39_, mshr_n_lru_paddr__38_, mshr_n_lru_paddr__37_, mshr_n_lru_paddr__36_, mshr_n_lru_paddr__35_, mshr_n_lru_paddr__34_, mshr_n_lru_paddr__33_, mshr_n_lru_paddr__32_, mshr_n_lru_paddr__31_, mshr_n_lru_paddr__30_, mshr_n_lru_paddr__29_, mshr_n_lru_paddr__28_, mshr_n_lru_paddr__27_, mshr_n_lru_paddr__26_, mshr_n_lru_paddr__25_, mshr_n_lru_paddr__24_, mshr_n_lru_paddr__23_, mshr_n_lru_paddr__22_, mshr_n_lru_paddr__21_, mshr_n_lru_paddr__20_, mshr_n_lru_paddr__19_, mshr_n_lru_paddr__18_, mshr_n_lru_paddr__17_, mshr_n_lru_paddr__16_, mshr_n_lru_paddr__15_, mshr_n_lru_paddr__14_, mshr_n_lru_paddr__13_, mshr_n_lru_paddr__12_, mshr_n_lru_paddr__11_, mshr_n_lru_paddr__10_, mshr_n_lru_paddr__9_, mshr_n_lru_paddr__8_, mshr_n_lru_paddr__7_, mshr_n_lru_paddr__6_, mshr_n_lru_way_id__2_, mshr_n_lru_way_id__1_, mshr_n_lru_way_id__0_, mshr_n_tr_lce_id__2_, mshr_n_tr_lce_id__1_, mshr_n_tr_lce_id__0_, mshr_n_tr_way_id__2_, mshr_n_tr_way_id__1_, mshr_n_tr_way_id__0_, mshr_n_next_coh_state__2_, mshr_n_next_coh_state__1_, mshr_n_next_coh_state__0_, mshr_n_flags__15_, mshr_n_flags__14_, mshr_n_flags__13_, mshr_n_flags__12_, mshr_n_flags__11_, mshr_n_flags__10_, mshr_n_flags__9_, mshr_n_flags__8_, mshr_n_flags__7_, mshr_n_flags__6_, mshr_n_flags__5_, mshr_n_flags__4_, mshr_n_flags__3_, mshr_n_flags__2_, mshr_n_flags__1_, mshr_n_flags__0_, mshr_n_uc_req_size__1_, mshr_n_uc_req_size__0_ } = (N128)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, coh_state_o, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 (N1333)? { N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, gad_req_addr_way_i, dir_lru_tag_i, mshr_o[87:82], N1435, N1434, N1433, gad_transfer_lce_i, gad_transfer_lce_way_i, decoded_inst_i[137:135], N1497, N1475, N1485, N1483, N1481, N1477, N1493, N1491, N1489, N1487, N1495, N1479, N1473, N1464, N1455, N1444, N1454, N1453 } : 1'b0;
  assign N128 = decoded_inst_i[10];
  assign N1500 = (N129)? 1'b1 : 
                 (N130)? decoded_inst_i[31] : 1'b0;
  assign N129 = dir_lru_v_i;
  assign N130 = N1499;
  assign { N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502 } = (N128)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                               (N1333)? { decoded_inst_i[24:23], dir_lru_v_i, decoded_inst_i[22:21], N1501, decoded_inst_i[41:32], N1500, decoded_inst_i[30:26], decoded_inst_i[17:17] } : 1'b0;
  assign { N1615, N1611, N1576, N1572, N1565, N1561, N1559, N1557, N1555, N1553, N1551, N1549, N1547, N1545, N1543, N1541, N1539, N1537, N1535, N1533, N1531, N1529, N1526 } = (N131)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                               (N132)? { N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502 } : 1'b0;
  assign N131 = reset_i;
  assign N132 = N1498;
  assign { N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1614, N1613, N1612, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1575, N1574, N1573, N1571, N1570, N1569, N1568, N1567, N1566, N1564, N1563, N1562, N1560, N1558, N1556, N1554, N1552, N1550, N1548, N1546, N1544, N1542, N1540, N1538, N1536, N1534, N1532, N1530, N1528, N1527 } = (N131)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (N132)? { mshr_n_lce_id__5_, mshr_n_lce_id__4_, mshr_n_lce_id__3_, mshr_n_lce_id__2_, mshr_n_lce_id__1_, mshr_n_lce_id__0_, mshr_n_paddr__39_, mshr_n_paddr__38_, mshr_n_paddr__37_, mshr_n_paddr__36_, mshr_n_paddr__35_, mshr_n_paddr__34_, mshr_n_paddr__33_, mshr_n_paddr__32_, mshr_n_paddr__31_, mshr_n_paddr__30_, mshr_n_paddr__29_, mshr_n_paddr__28_, mshr_n_paddr__27_, mshr_n_paddr__26_, mshr_n_paddr__25_, mshr_n_paddr__24_, mshr_n_paddr__23_, mshr_n_paddr__22_, mshr_n_paddr__21_, mshr_n_paddr__20_, mshr_n_paddr__19_, mshr_n_paddr__18_, mshr_n_paddr__17_, mshr_n_paddr__16_, mshr_n_paddr__15_, mshr_n_paddr__14_, mshr_n_paddr__13_, mshr_n_paddr__12_, mshr_n_paddr__11_, mshr_n_paddr__10_, mshr_n_paddr__9_, mshr_n_paddr__8_, mshr_n_paddr__7_, mshr_n_paddr__6_, mshr_n_paddr__5_, mshr_n_paddr__4_, mshr_n_paddr__3_, mshr_n_paddr__2_, mshr_n_paddr__1_, mshr_n_paddr__0_, mshr_n_way_id__2_, mshr_n_way_id__1_, mshr_n_way_id__0_, mshr_n_lru_paddr__39_, mshr_n_lru_paddr__38_, mshr_n_lru_paddr__37_, mshr_n_lru_paddr__36_, mshr_n_lru_paddr__35_, mshr_n_lru_paddr__34_, mshr_n_lru_paddr__33_, mshr_n_lru_paddr__32_, mshr_n_lru_paddr__31_, mshr_n_lru_paddr__30_, mshr_n_lru_paddr__29_, mshr_n_lru_paddr__28_, mshr_n_lru_paddr__27_, mshr_n_lru_paddr__26_, mshr_n_lru_paddr__25_, mshr_n_lru_paddr__24_, mshr_n_lru_paddr__23_, mshr_n_lru_paddr__22_, mshr_n_lru_paddr__21_, mshr_n_lru_paddr__20_, mshr_n_lru_paddr__19_, mshr_n_lru_paddr__18_, mshr_n_lru_paddr__17_, mshr_n_lru_paddr__16_, mshr_n_lru_paddr__15_, mshr_n_lru_paddr__14_, mshr_n_lru_paddr__13_, mshr_n_lru_paddr__12_, mshr_n_lru_paddr__11_, mshr_n_lru_paddr__10_, mshr_n_lru_paddr__9_, mshr_n_lru_paddr__8_, mshr_n_lru_paddr__7_, mshr_n_lru_paddr__6_, mshr_n_lru_way_id__2_, mshr_n_lru_way_id__1_, mshr_n_lru_way_id__0_, mshr_n_tr_lce_id__2_, mshr_n_tr_lce_id__1_, mshr_n_tr_lce_id__0_, mshr_n_tr_way_id__2_, mshr_n_tr_way_id__1_, mshr_n_tr_way_id__0_, mshr_n_next_coh_state__2_, mshr_n_next_coh_state__1_, mshr_n_next_coh_state__0_, mshr_n_flags__15_, mshr_n_flags__14_, mshr_n_flags__13_, mshr_n_flags__12_, mshr_n_flags__11_, mshr_n_flags__10_, mshr_n_flags__9_, mshr_n_flags__8_, mshr_n_flags__7_, mshr_n_flags__6_, mshr_n_flags__5_, mshr_n_flags__4_, mshr_n_flags__3_, mshr_n_flags__2_, mshr_n_flags__1_, mshr_n_flags__0_, mshr_n_uc_req_size__1_, mshr_n_uc_req_size__0_ } : 1'b0;
  assign { N2005, N1956, N1907, N1858, N1809, N1760, N1711, N1662 } = (N131)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                      (N132)? decoded_inst_i[49:42] : 1'b0;
  assign { N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663 } = (N131)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N132)? gpr_n : 1'b0;
  assign N2054 = (N131)? 1'b1 : 
                 (N132)? decoded_inst_i[18] : 1'b0;
  assign { N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055 } = (N131)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N132)? lce_req_i[118:55] : 1'b0;
  assign N2119 = (N131)? 1'b1 : 
                 (N132)? N1525 : 1'b0;
  assign { N2122, N2121, N2120 } = (N131)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N132)? mov_src_i[2:0] : 1'b0;
  assign uc_req = N2138 | N2141;
  assign N133 = decoded_inst_i[50] & decoded_inst_i[42];
  assign N134 = ~N133;
  assign N135 = decoded_inst_i[51] & decoded_inst_i[42];
  assign N136 = ~N135;
  assign N137 = decoded_inst_i[20] & decoded_inst_i[42];
  assign N138 = ~N137;
  assign N139 = decoded_inst_i[19] & decoded_inst_i[42];
  assign N140 = ~N139;
  assign N141 = N2147 & decoded_inst_i[42];
  assign N2147 = decoded_inst_i[85] & N2146;
  assign N142 = ~N141;
  assign N283 = decoded_inst_i[50] & decoded_inst_i[43];
  assign N284 = ~N283;
  assign N285 = decoded_inst_i[51] & decoded_inst_i[43];
  assign N286 = ~N285;
  assign N287 = decoded_inst_i[20] & decoded_inst_i[43];
  assign N288 = ~N287;
  assign N289 = decoded_inst_i[19] & decoded_inst_i[43];
  assign N290 = ~N289;
  assign N291 = N2148 & decoded_inst_i[43];
  assign N2148 = decoded_inst_i[85] & N2146;
  assign N292 = ~N291;
  assign N433 = decoded_inst_i[50] & decoded_inst_i[44];
  assign N434 = ~N433;
  assign N435 = decoded_inst_i[51] & decoded_inst_i[44];
  assign N436 = ~N435;
  assign N437 = decoded_inst_i[20] & decoded_inst_i[44];
  assign N438 = ~N437;
  assign N439 = decoded_inst_i[19] & decoded_inst_i[44];
  assign N440 = ~N439;
  assign N441 = N2149 & decoded_inst_i[44];
  assign N2149 = decoded_inst_i[85] & N2146;
  assign N442 = ~N441;
  assign N583 = decoded_inst_i[50] & decoded_inst_i[45];
  assign N584 = ~N583;
  assign N585 = decoded_inst_i[51] & decoded_inst_i[45];
  assign N586 = ~N585;
  assign N587 = decoded_inst_i[20] & decoded_inst_i[45];
  assign N588 = ~N587;
  assign N589 = decoded_inst_i[19] & decoded_inst_i[45];
  assign N590 = ~N589;
  assign N591 = N2150 & decoded_inst_i[45];
  assign N2150 = decoded_inst_i[85] & N2146;
  assign N592 = ~N591;
  assign N733 = decoded_inst_i[50] & decoded_inst_i[46];
  assign N734 = ~N733;
  assign N735 = decoded_inst_i[51] & decoded_inst_i[46];
  assign N736 = ~N735;
  assign N737 = decoded_inst_i[20] & decoded_inst_i[46];
  assign N738 = ~N737;
  assign N739 = decoded_inst_i[19] & decoded_inst_i[46];
  assign N740 = ~N739;
  assign N741 = N2151 & decoded_inst_i[46];
  assign N2151 = decoded_inst_i[85] & N2146;
  assign N742 = ~N741;
  assign N883 = decoded_inst_i[50] & decoded_inst_i[47];
  assign N884 = ~N883;
  assign N885 = decoded_inst_i[51] & decoded_inst_i[47];
  assign N886 = ~N885;
  assign N887 = decoded_inst_i[20] & decoded_inst_i[47];
  assign N888 = ~N887;
  assign N889 = decoded_inst_i[19] & decoded_inst_i[47];
  assign N890 = ~N889;
  assign N891 = N2152 & decoded_inst_i[47];
  assign N2152 = decoded_inst_i[85] & N2146;
  assign N892 = ~N891;
  assign N1033 = decoded_inst_i[50] & decoded_inst_i[48];
  assign N1034 = ~N1033;
  assign N1035 = decoded_inst_i[51] & decoded_inst_i[48];
  assign N1036 = ~N1035;
  assign N1037 = decoded_inst_i[20] & decoded_inst_i[48];
  assign N1038 = ~N1037;
  assign N1039 = decoded_inst_i[19] & decoded_inst_i[48];
  assign N1040 = ~N1039;
  assign N1041 = N2153 & decoded_inst_i[48];
  assign N2153 = decoded_inst_i[85] & N2146;
  assign N1042 = ~N1041;
  assign N1183 = decoded_inst_i[50] & decoded_inst_i[49];
  assign N1184 = ~N1183;
  assign N1185 = decoded_inst_i[51] & decoded_inst_i[49];
  assign N1186 = ~N1185;
  assign N1187 = decoded_inst_i[20] & decoded_inst_i[49];
  assign N1188 = ~N1187;
  assign N1189 = decoded_inst_i[19] & decoded_inst_i[49];
  assign N1190 = ~N1189;
  assign N1191 = N2154 & decoded_inst_i[49];
  assign N2154 = decoded_inst_i[85] & N2146;
  assign N1192 = ~N1191;
  assign N1333 = ~decoded_inst_i[10];
  assign N1334 = ~decoded_inst_i[129];
  assign N1335 = ~decoded_inst_i[128];
  assign N1428 = ~decoded_inst_i[127];
  assign N1429 = ~decoded_inst_i[126];
  assign N1436 = ~decoded_inst_i[125];
  assign N1437 = ~decoded_inst_i[124];
  assign N1440 = ~N1439;
  assign N1442 = ~N1441;
  assign N1445 = ~decoded_inst_i[123];
  assign N1446 = ~decoded_inst_i[122];
  assign N1449 = ~N1448;
  assign N1451 = ~N1450;
  assign N1456 = ~decoded_inst_i[121];
  assign N1457 = ~decoded_inst_i[120];
  assign N1460 = ~N1459;
  assign N1462 = ~N1461;
  assign N1465 = ~decoded_inst_i[119];
  assign N1466 = ~decoded_inst_i[118];
  assign N1469 = ~N1468;
  assign N1471 = ~N1470;
  assign N1474 = ~decoded_inst_i[107];
  assign N1476 = ~decoded_inst_i[111];
  assign N1478 = ~decoded_inst_i[117];
  assign N1480 = ~decoded_inst_i[110];
  assign N1482 = ~decoded_inst_i[109];
  assign N1484 = ~decoded_inst_i[108];
  assign N1486 = ~decoded_inst_i[115];
  assign N1488 = ~decoded_inst_i[114];
  assign N1490 = ~decoded_inst_i[113];
  assign N1492 = ~decoded_inst_i[112];
  assign N1494 = ~decoded_inst_i[116];
  assign N1496 = ~decoded_inst_i[106];
  assign N1498 = ~reset_i;
  assign N1499 = ~dir_lru_v_i;
  assign N1501 = N2155 & N2134;
  assign N2155 = decoded_inst_i[51] & N2125;
  assign N1525 = N2156 & N2131;
  assign N2156 = decoded_inst_i[51] & N2125;

endmodule