module bsg_mem_1r1w_synth_width_p76_els_p4_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [1:0] w_addr_i;
  input [75:0] w_data_i;
  input [1:0] r_addr_i;
  output [75:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [75:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20;
  reg [303:0] mem;
  assign r_data_o[75] = (N8)? mem[75] : 
                        (N10)? mem[151] : 
                        (N9)? mem[227] : 
                        (N11)? mem[303] : 1'b0;
  assign r_data_o[74] = (N8)? mem[74] : 
                        (N10)? mem[150] : 
                        (N9)? mem[226] : 
                        (N11)? mem[302] : 1'b0;
  assign r_data_o[73] = (N8)? mem[73] : 
                        (N10)? mem[149] : 
                        (N9)? mem[225] : 
                        (N11)? mem[301] : 1'b0;
  assign r_data_o[72] = (N8)? mem[72] : 
                        (N10)? mem[148] : 
                        (N9)? mem[224] : 
                        (N11)? mem[300] : 1'b0;
  assign r_data_o[71] = (N8)? mem[71] : 
                        (N10)? mem[147] : 
                        (N9)? mem[223] : 
                        (N11)? mem[299] : 1'b0;
  assign r_data_o[70] = (N8)? mem[70] : 
                        (N10)? mem[146] : 
                        (N9)? mem[222] : 
                        (N11)? mem[298] : 1'b0;
  assign r_data_o[69] = (N8)? mem[69] : 
                        (N10)? mem[145] : 
                        (N9)? mem[221] : 
                        (N11)? mem[297] : 1'b0;
  assign r_data_o[68] = (N8)? mem[68] : 
                        (N10)? mem[144] : 
                        (N9)? mem[220] : 
                        (N11)? mem[296] : 1'b0;
  assign r_data_o[67] = (N8)? mem[67] : 
                        (N10)? mem[143] : 
                        (N9)? mem[219] : 
                        (N11)? mem[295] : 1'b0;
  assign r_data_o[66] = (N8)? mem[66] : 
                        (N10)? mem[142] : 
                        (N9)? mem[218] : 
                        (N11)? mem[294] : 1'b0;
  assign r_data_o[65] = (N8)? mem[65] : 
                        (N10)? mem[141] : 
                        (N9)? mem[217] : 
                        (N11)? mem[293] : 1'b0;
  assign r_data_o[64] = (N8)? mem[64] : 
                        (N10)? mem[140] : 
                        (N9)? mem[216] : 
                        (N11)? mem[292] : 1'b0;
  assign r_data_o[63] = (N8)? mem[63] : 
                        (N10)? mem[139] : 
                        (N9)? mem[215] : 
                        (N11)? mem[291] : 1'b0;
  assign r_data_o[62] = (N8)? mem[62] : 
                        (N10)? mem[138] : 
                        (N9)? mem[214] : 
                        (N11)? mem[290] : 1'b0;
  assign r_data_o[61] = (N8)? mem[61] : 
                        (N10)? mem[137] : 
                        (N9)? mem[213] : 
                        (N11)? mem[289] : 1'b0;
  assign r_data_o[60] = (N8)? mem[60] : 
                        (N10)? mem[136] : 
                        (N9)? mem[212] : 
                        (N11)? mem[288] : 1'b0;
  assign r_data_o[59] = (N8)? mem[59] : 
                        (N10)? mem[135] : 
                        (N9)? mem[211] : 
                        (N11)? mem[287] : 1'b0;
  assign r_data_o[58] = (N8)? mem[58] : 
                        (N10)? mem[134] : 
                        (N9)? mem[210] : 
                        (N11)? mem[286] : 1'b0;
  assign r_data_o[57] = (N8)? mem[57] : 
                        (N10)? mem[133] : 
                        (N9)? mem[209] : 
                        (N11)? mem[285] : 1'b0;
  assign r_data_o[56] = (N8)? mem[56] : 
                        (N10)? mem[132] : 
                        (N9)? mem[208] : 
                        (N11)? mem[284] : 1'b0;
  assign r_data_o[55] = (N8)? mem[55] : 
                        (N10)? mem[131] : 
                        (N9)? mem[207] : 
                        (N11)? mem[283] : 1'b0;
  assign r_data_o[54] = (N8)? mem[54] : 
                        (N10)? mem[130] : 
                        (N9)? mem[206] : 
                        (N11)? mem[282] : 1'b0;
  assign r_data_o[53] = (N8)? mem[53] : 
                        (N10)? mem[129] : 
                        (N9)? mem[205] : 
                        (N11)? mem[281] : 1'b0;
  assign r_data_o[52] = (N8)? mem[52] : 
                        (N10)? mem[128] : 
                        (N9)? mem[204] : 
                        (N11)? mem[280] : 1'b0;
  assign r_data_o[51] = (N8)? mem[51] : 
                        (N10)? mem[127] : 
                        (N9)? mem[203] : 
                        (N11)? mem[279] : 1'b0;
  assign r_data_o[50] = (N8)? mem[50] : 
                        (N10)? mem[126] : 
                        (N9)? mem[202] : 
                        (N11)? mem[278] : 1'b0;
  assign r_data_o[49] = (N8)? mem[49] : 
                        (N10)? mem[125] : 
                        (N9)? mem[201] : 
                        (N11)? mem[277] : 1'b0;
  assign r_data_o[48] = (N8)? mem[48] : 
                        (N10)? mem[124] : 
                        (N9)? mem[200] : 
                        (N11)? mem[276] : 1'b0;
  assign r_data_o[47] = (N8)? mem[47] : 
                        (N10)? mem[123] : 
                        (N9)? mem[199] : 
                        (N11)? mem[275] : 1'b0;
  assign r_data_o[46] = (N8)? mem[46] : 
                        (N10)? mem[122] : 
                        (N9)? mem[198] : 
                        (N11)? mem[274] : 1'b0;
  assign r_data_o[45] = (N8)? mem[45] : 
                        (N10)? mem[121] : 
                        (N9)? mem[197] : 
                        (N11)? mem[273] : 1'b0;
  assign r_data_o[44] = (N8)? mem[44] : 
                        (N10)? mem[120] : 
                        (N9)? mem[196] : 
                        (N11)? mem[272] : 1'b0;
  assign r_data_o[43] = (N8)? mem[43] : 
                        (N10)? mem[119] : 
                        (N9)? mem[195] : 
                        (N11)? mem[271] : 1'b0;
  assign r_data_o[42] = (N8)? mem[42] : 
                        (N10)? mem[118] : 
                        (N9)? mem[194] : 
                        (N11)? mem[270] : 1'b0;
  assign r_data_o[41] = (N8)? mem[41] : 
                        (N10)? mem[117] : 
                        (N9)? mem[193] : 
                        (N11)? mem[269] : 1'b0;
  assign r_data_o[40] = (N8)? mem[40] : 
                        (N10)? mem[116] : 
                        (N9)? mem[192] : 
                        (N11)? mem[268] : 1'b0;
  assign r_data_o[39] = (N8)? mem[39] : 
                        (N10)? mem[115] : 
                        (N9)? mem[191] : 
                        (N11)? mem[267] : 1'b0;
  assign r_data_o[38] = (N8)? mem[38] : 
                        (N10)? mem[114] : 
                        (N9)? mem[190] : 
                        (N11)? mem[266] : 1'b0;
  assign r_data_o[37] = (N8)? mem[37] : 
                        (N10)? mem[113] : 
                        (N9)? mem[189] : 
                        (N11)? mem[265] : 1'b0;
  assign r_data_o[36] = (N8)? mem[36] : 
                        (N10)? mem[112] : 
                        (N9)? mem[188] : 
                        (N11)? mem[264] : 1'b0;
  assign r_data_o[35] = (N8)? mem[35] : 
                        (N10)? mem[111] : 
                        (N9)? mem[187] : 
                        (N11)? mem[263] : 1'b0;
  assign r_data_o[34] = (N8)? mem[34] : 
                        (N10)? mem[110] : 
                        (N9)? mem[186] : 
                        (N11)? mem[262] : 1'b0;
  assign r_data_o[33] = (N8)? mem[33] : 
                        (N10)? mem[109] : 
                        (N9)? mem[185] : 
                        (N11)? mem[261] : 1'b0;
  assign r_data_o[32] = (N8)? mem[32] : 
                        (N10)? mem[108] : 
                        (N9)? mem[184] : 
                        (N11)? mem[260] : 1'b0;
  assign r_data_o[31] = (N8)? mem[31] : 
                        (N10)? mem[107] : 
                        (N9)? mem[183] : 
                        (N11)? mem[259] : 1'b0;
  assign r_data_o[30] = (N8)? mem[30] : 
                        (N10)? mem[106] : 
                        (N9)? mem[182] : 
                        (N11)? mem[258] : 1'b0;
  assign r_data_o[29] = (N8)? mem[29] : 
                        (N10)? mem[105] : 
                        (N9)? mem[181] : 
                        (N11)? mem[257] : 1'b0;
  assign r_data_o[28] = (N8)? mem[28] : 
                        (N10)? mem[104] : 
                        (N9)? mem[180] : 
                        (N11)? mem[256] : 1'b0;
  assign r_data_o[27] = (N8)? mem[27] : 
                        (N10)? mem[103] : 
                        (N9)? mem[179] : 
                        (N11)? mem[255] : 1'b0;
  assign r_data_o[26] = (N8)? mem[26] : 
                        (N10)? mem[102] : 
                        (N9)? mem[178] : 
                        (N11)? mem[254] : 1'b0;
  assign r_data_o[25] = (N8)? mem[25] : 
                        (N10)? mem[101] : 
                        (N9)? mem[177] : 
                        (N11)? mem[253] : 1'b0;
  assign r_data_o[24] = (N8)? mem[24] : 
                        (N10)? mem[100] : 
                        (N9)? mem[176] : 
                        (N11)? mem[252] : 1'b0;
  assign r_data_o[23] = (N8)? mem[23] : 
                        (N10)? mem[99] : 
                        (N9)? mem[175] : 
                        (N11)? mem[251] : 1'b0;
  assign r_data_o[22] = (N8)? mem[22] : 
                        (N10)? mem[98] : 
                        (N9)? mem[174] : 
                        (N11)? mem[250] : 1'b0;
  assign r_data_o[21] = (N8)? mem[21] : 
                        (N10)? mem[97] : 
                        (N9)? mem[173] : 
                        (N11)? mem[249] : 1'b0;
  assign r_data_o[20] = (N8)? mem[20] : 
                        (N10)? mem[96] : 
                        (N9)? mem[172] : 
                        (N11)? mem[248] : 1'b0;
  assign r_data_o[19] = (N8)? mem[19] : 
                        (N10)? mem[95] : 
                        (N9)? mem[171] : 
                        (N11)? mem[247] : 1'b0;
  assign r_data_o[18] = (N8)? mem[18] : 
                        (N10)? mem[94] : 
                        (N9)? mem[170] : 
                        (N11)? mem[246] : 1'b0;
  assign r_data_o[17] = (N8)? mem[17] : 
                        (N10)? mem[93] : 
                        (N9)? mem[169] : 
                        (N11)? mem[245] : 1'b0;
  assign r_data_o[16] = (N8)? mem[16] : 
                        (N10)? mem[92] : 
                        (N9)? mem[168] : 
                        (N11)? mem[244] : 1'b0;
  assign r_data_o[15] = (N8)? mem[15] : 
                        (N10)? mem[91] : 
                        (N9)? mem[167] : 
                        (N11)? mem[243] : 1'b0;
  assign r_data_o[14] = (N8)? mem[14] : 
                        (N10)? mem[90] : 
                        (N9)? mem[166] : 
                        (N11)? mem[242] : 1'b0;
  assign r_data_o[13] = (N8)? mem[13] : 
                        (N10)? mem[89] : 
                        (N9)? mem[165] : 
                        (N11)? mem[241] : 1'b0;
  assign r_data_o[12] = (N8)? mem[12] : 
                        (N10)? mem[88] : 
                        (N9)? mem[164] : 
                        (N11)? mem[240] : 1'b0;
  assign r_data_o[11] = (N8)? mem[11] : 
                        (N10)? mem[87] : 
                        (N9)? mem[163] : 
                        (N11)? mem[239] : 1'b0;
  assign r_data_o[10] = (N8)? mem[10] : 
                        (N10)? mem[86] : 
                        (N9)? mem[162] : 
                        (N11)? mem[238] : 1'b0;
  assign r_data_o[9] = (N8)? mem[9] : 
                       (N10)? mem[85] : 
                       (N9)? mem[161] : 
                       (N11)? mem[237] : 1'b0;
  assign r_data_o[8] = (N8)? mem[8] : 
                       (N10)? mem[84] : 
                       (N9)? mem[160] : 
                       (N11)? mem[236] : 1'b0;
  assign r_data_o[7] = (N8)? mem[7] : 
                       (N10)? mem[83] : 
                       (N9)? mem[159] : 
                       (N11)? mem[235] : 1'b0;
  assign r_data_o[6] = (N8)? mem[6] : 
                       (N10)? mem[82] : 
                       (N9)? mem[158] : 
                       (N11)? mem[234] : 1'b0;
  assign r_data_o[5] = (N8)? mem[5] : 
                       (N10)? mem[81] : 
                       (N9)? mem[157] : 
                       (N11)? mem[233] : 1'b0;
  assign r_data_o[4] = (N8)? mem[4] : 
                       (N10)? mem[80] : 
                       (N9)? mem[156] : 
                       (N11)? mem[232] : 1'b0;
  assign r_data_o[3] = (N8)? mem[3] : 
                       (N10)? mem[79] : 
                       (N9)? mem[155] : 
                       (N11)? mem[231] : 1'b0;
  assign r_data_o[2] = (N8)? mem[2] : 
                       (N10)? mem[78] : 
                       (N9)? mem[154] : 
                       (N11)? mem[230] : 1'b0;
  assign r_data_o[1] = (N8)? mem[1] : 
                       (N10)? mem[77] : 
                       (N9)? mem[153] : 
                       (N11)? mem[229] : 1'b0;
  assign r_data_o[0] = (N8)? mem[0] : 
                       (N10)? mem[76] : 
                       (N9)? mem[152] : 
                       (N11)? mem[228] : 1'b0;

  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[303] <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[302] <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[301] <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[300] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[299] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[298] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[297] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[296] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[295] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[294] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[293] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[292] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[291] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[290] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[289] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[288] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[287] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[286] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[285] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[284] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[283] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[282] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[281] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[280] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[279] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[278] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[277] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[276] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[275] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[274] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[273] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[272] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[271] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[270] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[269] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[268] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[267] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[266] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[265] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[264] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[263] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[262] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[261] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[260] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[259] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[258] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[257] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[256] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[255] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[254] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[253] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[252] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[251] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[250] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[249] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[248] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[247] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[246] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[245] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[244] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[243] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[242] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[241] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[240] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[239] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[238] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[237] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[236] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[235] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[234] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[233] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[232] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[231] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[230] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[229] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N20) begin
      mem[228] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[227] <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[226] <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[225] <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[224] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[223] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[222] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[221] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[220] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[219] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[218] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[217] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[216] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[215] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[214] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[213] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[212] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[211] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[210] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[209] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[208] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[207] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[206] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[205] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[204] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[203] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[202] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[201] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[200] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[199] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[198] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[197] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[196] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[195] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[194] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[193] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[192] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[191] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[190] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[189] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[188] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[187] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[186] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[185] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[184] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[183] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[182] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[181] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[180] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[179] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[178] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[177] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[176] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[175] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[174] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[173] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[172] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[171] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[170] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[169] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[168] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[167] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[166] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[165] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[164] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[163] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[162] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[161] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[160] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[159] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[158] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[157] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[156] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[155] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[154] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[153] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N19) begin
      mem[152] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[151] <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[150] <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[149] <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[148] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[147] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[146] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[145] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[144] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[143] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[142] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[141] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[140] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[139] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[138] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[137] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[136] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[135] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[134] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[133] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[132] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[131] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[130] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[129] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[128] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[127] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[126] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[125] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[124] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[123] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[122] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[121] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[120] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[119] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[118] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[117] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[116] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[115] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[114] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[113] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[112] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[111] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[110] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[109] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[108] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[107] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[106] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[105] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[104] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[103] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[102] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[101] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[100] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[99] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[98] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[97] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[96] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[95] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[94] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[93] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[92] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[91] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[90] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[89] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[88] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[87] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[86] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[85] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[84] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[83] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[82] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[81] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[80] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[79] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[78] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[77] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N18) begin
      mem[76] <= w_data_i[0];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[75] <= w_data_i[75];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[74] <= w_data_i[74];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[73] <= w_data_i[73];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[72] <= w_data_i[72];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[71] <= w_data_i[71];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[70] <= w_data_i[70];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[69] <= w_data_i[69];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[68] <= w_data_i[68];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[67] <= w_data_i[67];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[66] <= w_data_i[66];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[65] <= w_data_i[65];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[64] <= w_data_i[64];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[63] <= w_data_i[63];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[62] <= w_data_i[62];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[61] <= w_data_i[61];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[60] <= w_data_i[60];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[59] <= w_data_i[59];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[58] <= w_data_i[58];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[57] <= w_data_i[57];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[56] <= w_data_i[56];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[55] <= w_data_i[55];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[54] <= w_data_i[54];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[53] <= w_data_i[53];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[52] <= w_data_i[52];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[51] <= w_data_i[51];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[50] <= w_data_i[50];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[49] <= w_data_i[49];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[48] <= w_data_i[48];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[47] <= w_data_i[47];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[46] <= w_data_i[46];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[45] <= w_data_i[45];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[44] <= w_data_i[44];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[43] <= w_data_i[43];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[42] <= w_data_i[42];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[41] <= w_data_i[41];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[40] <= w_data_i[40];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[39] <= w_data_i[39];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[38] <= w_data_i[38];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[37] <= w_data_i[37];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[36] <= w_data_i[36];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[35] <= w_data_i[35];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[34] <= w_data_i[34];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[33] <= w_data_i[33];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[32] <= w_data_i[32];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[31] <= w_data_i[31];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[30] <= w_data_i[30];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[29] <= w_data_i[29];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[28] <= w_data_i[28];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[27] <= w_data_i[27];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[26] <= w_data_i[26];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[25] <= w_data_i[25];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[24] <= w_data_i[24];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[23] <= w_data_i[23];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[22] <= w_data_i[22];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[21] <= w_data_i[21];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[20] <= w_data_i[20];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[19] <= w_data_i[19];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[18] <= w_data_i[18];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[17] <= w_data_i[17];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[16] <= w_data_i[16];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[15] <= w_data_i[15];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[14] <= w_data_i[14];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[13] <= w_data_i[13];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[12] <= w_data_i[12];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[11] <= w_data_i[11];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[10] <= w_data_i[10];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[9] <= w_data_i[9];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[8] <= w_data_i[8];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[7] <= w_data_i[7];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[6] <= w_data_i[6];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[5] <= w_data_i[5];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[4] <= w_data_i[4];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[3] <= w_data_i[3];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[2] <= w_data_i[2];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[1] <= w_data_i[1];
    end 
  end


  always @(posedge w_clk_i) begin
    if(N17) begin
      mem[0] <= w_data_i[0];
    end 
  end

  assign N16 = w_addr_i[0] & w_addr_i[1];
  assign N15 = N0 & w_addr_i[1];
  assign N0 = ~w_addr_i[0];
  assign N14 = w_addr_i[0] & N1;
  assign N1 = ~w_addr_i[1];
  assign N13 = N2 & N3;
  assign N2 = ~w_addr_i[0];
  assign N3 = ~w_addr_i[1];
  assign { N20, N19, N18, N17 } = (N4)? { N16, N15, N14, N13 } : 
                                  (N5)? { 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N4 = w_v_i;
  assign N5 = N12;
  assign N6 = ~r_addr_i[0];
  assign N7 = ~r_addr_i[1];
  assign N8 = N6 & N7;
  assign N9 = N6 & r_addr_i[1];
  assign N10 = r_addr_i[0] & N7;
  assign N11 = r_addr_i[0] & r_addr_i[1];
  assign N12 = ~w_v_i;

endmodule