module btb_NR_ENTRIES64
(
  clk_i,
  rst_ni,
  flush_i,
  debug_mode_i,
  vpc_i,
  btb_update_i,
  btb_prediction_o
);

  input [63:0] vpc_i;
  input [129:0] btb_update_i;
  output [64:0] btb_prediction_o;
  input clk_i;
  input rst_ni;
  input flush_i;
  input debug_mode_i;
  wire [64:0] btb_prediction_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520;
  reg [4159:0] btb_q;
  assign btb_prediction_o[64] = (N141)? btb_q[64] : 
                                (N143)? btb_q[129] : 
                                (N145)? btb_q[194] : 
                                (N147)? btb_q[259] : 
                                (N149)? btb_q[324] : 
                                (N151)? btb_q[389] : 
                                (N153)? btb_q[454] : 
                                (N155)? btb_q[519] : 
                                (N157)? btb_q[584] : 
                                (N159)? btb_q[649] : 
                                (N161)? btb_q[714] : 
                                (N163)? btb_q[779] : 
                                (N165)? btb_q[844] : 
                                (N167)? btb_q[909] : 
                                (N169)? btb_q[974] : 
                                (N171)? btb_q[1039] : 
                                (N173)? btb_q[1104] : 
                                (N175)? btb_q[1169] : 
                                (N177)? btb_q[1234] : 
                                (N179)? btb_q[1299] : 
                                (N181)? btb_q[1364] : 
                                (N183)? btb_q[1429] : 
                                (N185)? btb_q[1494] : 
                                (N187)? btb_q[1559] : 
                                (N189)? btb_q[1624] : 
                                (N191)? btb_q[1689] : 
                                (N193)? btb_q[1754] : 
                                (N195)? btb_q[1819] : 
                                (N197)? btb_q[1884] : 
                                (N199)? btb_q[1949] : 
                                (N201)? btb_q[2014] : 
                                (N203)? btb_q[2079] : 
                                (N142)? btb_q[2144] : 
                                (N144)? btb_q[2209] : 
                                (N146)? btb_q[2274] : 
                                (N148)? btb_q[2339] : 
                                (N150)? btb_q[2404] : 
                                (N152)? btb_q[2469] : 
                                (N154)? btb_q[2534] : 
                                (N156)? btb_q[2599] : 
                                (N158)? btb_q[2664] : 
                                (N160)? btb_q[2729] : 
                                (N162)? btb_q[2794] : 
                                (N164)? btb_q[2859] : 
                                (N166)? btb_q[2924] : 
                                (N168)? btb_q[2989] : 
                                (N170)? btb_q[3054] : 
                                (N172)? btb_q[3119] : 
                                (N174)? btb_q[3184] : 
                                (N176)? btb_q[3249] : 
                                (N178)? btb_q[3314] : 
                                (N180)? btb_q[3379] : 
                                (N182)? btb_q[3444] : 
                                (N184)? btb_q[3509] : 
                                (N186)? btb_q[3574] : 
                                (N188)? btb_q[3639] : 
                                (N190)? btb_q[3704] : 
                                (N192)? btb_q[3769] : 
                                (N194)? btb_q[3834] : 
                                (N196)? btb_q[3899] : 
                                (N198)? btb_q[3964] : 
                                (N200)? btb_q[4029] : 
                                (N202)? btb_q[4094] : 
                                (N204)? btb_q[4159] : 1'b0;
  assign btb_prediction_o[63] = (N141)? btb_q[63] : 
                                (N143)? btb_q[128] : 
                                (N145)? btb_q[193] : 
                                (N147)? btb_q[258] : 
                                (N149)? btb_q[323] : 
                                (N151)? btb_q[388] : 
                                (N153)? btb_q[453] : 
                                (N155)? btb_q[518] : 
                                (N157)? btb_q[583] : 
                                (N159)? btb_q[648] : 
                                (N161)? btb_q[713] : 
                                (N163)? btb_q[778] : 
                                (N165)? btb_q[843] : 
                                (N167)? btb_q[908] : 
                                (N169)? btb_q[973] : 
                                (N171)? btb_q[1038] : 
                                (N173)? btb_q[1103] : 
                                (N175)? btb_q[1168] : 
                                (N177)? btb_q[1233] : 
                                (N179)? btb_q[1298] : 
                                (N181)? btb_q[1363] : 
                                (N183)? btb_q[1428] : 
                                (N185)? btb_q[1493] : 
                                (N187)? btb_q[1558] : 
                                (N189)? btb_q[1623] : 
                                (N191)? btb_q[1688] : 
                                (N193)? btb_q[1753] : 
                                (N195)? btb_q[1818] : 
                                (N197)? btb_q[1883] : 
                                (N199)? btb_q[1948] : 
                                (N201)? btb_q[2013] : 
                                (N203)? btb_q[2078] : 
                                (N142)? btb_q[2143] : 
                                (N144)? btb_q[2208] : 
                                (N146)? btb_q[2273] : 
                                (N148)? btb_q[2338] : 
                                (N150)? btb_q[2403] : 
                                (N152)? btb_q[2468] : 
                                (N154)? btb_q[2533] : 
                                (N156)? btb_q[2598] : 
                                (N158)? btb_q[2663] : 
                                (N160)? btb_q[2728] : 
                                (N162)? btb_q[2793] : 
                                (N164)? btb_q[2858] : 
                                (N166)? btb_q[2923] : 
                                (N168)? btb_q[2988] : 
                                (N170)? btb_q[3053] : 
                                (N172)? btb_q[3118] : 
                                (N174)? btb_q[3183] : 
                                (N176)? btb_q[3248] : 
                                (N178)? btb_q[3313] : 
                                (N180)? btb_q[3378] : 
                                (N182)? btb_q[3443] : 
                                (N184)? btb_q[3508] : 
                                (N186)? btb_q[3573] : 
                                (N188)? btb_q[3638] : 
                                (N190)? btb_q[3703] : 
                                (N192)? btb_q[3768] : 
                                (N194)? btb_q[3833] : 
                                (N196)? btb_q[3898] : 
                                (N198)? btb_q[3963] : 
                                (N200)? btb_q[4028] : 
                                (N202)? btb_q[4093] : 
                                (N204)? btb_q[4158] : 1'b0;
  assign btb_prediction_o[62] = (N141)? btb_q[62] : 
                                (N143)? btb_q[127] : 
                                (N145)? btb_q[192] : 
                                (N147)? btb_q[257] : 
                                (N149)? btb_q[322] : 
                                (N151)? btb_q[387] : 
                                (N153)? btb_q[452] : 
                                (N155)? btb_q[517] : 
                                (N157)? btb_q[582] : 
                                (N159)? btb_q[647] : 
                                (N161)? btb_q[712] : 
                                (N163)? btb_q[777] : 
                                (N165)? btb_q[842] : 
                                (N167)? btb_q[907] : 
                                (N169)? btb_q[972] : 
                                (N171)? btb_q[1037] : 
                                (N173)? btb_q[1102] : 
                                (N175)? btb_q[1167] : 
                                (N177)? btb_q[1232] : 
                                (N179)? btb_q[1297] : 
                                (N181)? btb_q[1362] : 
                                (N183)? btb_q[1427] : 
                                (N185)? btb_q[1492] : 
                                (N187)? btb_q[1557] : 
                                (N189)? btb_q[1622] : 
                                (N191)? btb_q[1687] : 
                                (N193)? btb_q[1752] : 
                                (N195)? btb_q[1817] : 
                                (N197)? btb_q[1882] : 
                                (N199)? btb_q[1947] : 
                                (N201)? btb_q[2012] : 
                                (N203)? btb_q[2077] : 
                                (N142)? btb_q[2142] : 
                                (N144)? btb_q[2207] : 
                                (N146)? btb_q[2272] : 
                                (N148)? btb_q[2337] : 
                                (N150)? btb_q[2402] : 
                                (N152)? btb_q[2467] : 
                                (N154)? btb_q[2532] : 
                                (N156)? btb_q[2597] : 
                                (N158)? btb_q[2662] : 
                                (N160)? btb_q[2727] : 
                                (N162)? btb_q[2792] : 
                                (N164)? btb_q[2857] : 
                                (N166)? btb_q[2922] : 
                                (N168)? btb_q[2987] : 
                                (N170)? btb_q[3052] : 
                                (N172)? btb_q[3117] : 
                                (N174)? btb_q[3182] : 
                                (N176)? btb_q[3247] : 
                                (N178)? btb_q[3312] : 
                                (N180)? btb_q[3377] : 
                                (N182)? btb_q[3442] : 
                                (N184)? btb_q[3507] : 
                                (N186)? btb_q[3572] : 
                                (N188)? btb_q[3637] : 
                                (N190)? btb_q[3702] : 
                                (N192)? btb_q[3767] : 
                                (N194)? btb_q[3832] : 
                                (N196)? btb_q[3897] : 
                                (N198)? btb_q[3962] : 
                                (N200)? btb_q[4027] : 
                                (N202)? btb_q[4092] : 
                                (N204)? btb_q[4157] : 1'b0;
  assign btb_prediction_o[61] = (N141)? btb_q[61] : 
                                (N143)? btb_q[126] : 
                                (N145)? btb_q[191] : 
                                (N147)? btb_q[256] : 
                                (N149)? btb_q[321] : 
                                (N151)? btb_q[386] : 
                                (N153)? btb_q[451] : 
                                (N155)? btb_q[516] : 
                                (N157)? btb_q[581] : 
                                (N159)? btb_q[646] : 
                                (N161)? btb_q[711] : 
                                (N163)? btb_q[776] : 
                                (N165)? btb_q[841] : 
                                (N167)? btb_q[906] : 
                                (N169)? btb_q[971] : 
                                (N171)? btb_q[1036] : 
                                (N173)? btb_q[1101] : 
                                (N175)? btb_q[1166] : 
                                (N177)? btb_q[1231] : 
                                (N179)? btb_q[1296] : 
                                (N181)? btb_q[1361] : 
                                (N183)? btb_q[1426] : 
                                (N185)? btb_q[1491] : 
                                (N187)? btb_q[1556] : 
                                (N189)? btb_q[1621] : 
                                (N191)? btb_q[1686] : 
                                (N193)? btb_q[1751] : 
                                (N195)? btb_q[1816] : 
                                (N197)? btb_q[1881] : 
                                (N199)? btb_q[1946] : 
                                (N201)? btb_q[2011] : 
                                (N203)? btb_q[2076] : 
                                (N142)? btb_q[2141] : 
                                (N144)? btb_q[2206] : 
                                (N146)? btb_q[2271] : 
                                (N148)? btb_q[2336] : 
                                (N150)? btb_q[2401] : 
                                (N152)? btb_q[2466] : 
                                (N154)? btb_q[2531] : 
                                (N156)? btb_q[2596] : 
                                (N158)? btb_q[2661] : 
                                (N160)? btb_q[2726] : 
                                (N162)? btb_q[2791] : 
                                (N164)? btb_q[2856] : 
                                (N166)? btb_q[2921] : 
                                (N168)? btb_q[2986] : 
                                (N170)? btb_q[3051] : 
                                (N172)? btb_q[3116] : 
                                (N174)? btb_q[3181] : 
                                (N176)? btb_q[3246] : 
                                (N178)? btb_q[3311] : 
                                (N180)? btb_q[3376] : 
                                (N182)? btb_q[3441] : 
                                (N184)? btb_q[3506] : 
                                (N186)? btb_q[3571] : 
                                (N188)? btb_q[3636] : 
                                (N190)? btb_q[3701] : 
                                (N192)? btb_q[3766] : 
                                (N194)? btb_q[3831] : 
                                (N196)? btb_q[3896] : 
                                (N198)? btb_q[3961] : 
                                (N200)? btb_q[4026] : 
                                (N202)? btb_q[4091] : 
                                (N204)? btb_q[4156] : 1'b0;
  assign btb_prediction_o[60] = (N141)? btb_q[60] : 
                                (N143)? btb_q[125] : 
                                (N145)? btb_q[190] : 
                                (N147)? btb_q[255] : 
                                (N149)? btb_q[320] : 
                                (N151)? btb_q[385] : 
                                (N153)? btb_q[450] : 
                                (N155)? btb_q[515] : 
                                (N157)? btb_q[580] : 
                                (N159)? btb_q[645] : 
                                (N161)? btb_q[710] : 
                                (N163)? btb_q[775] : 
                                (N165)? btb_q[840] : 
                                (N167)? btb_q[905] : 
                                (N169)? btb_q[970] : 
                                (N171)? btb_q[1035] : 
                                (N173)? btb_q[1100] : 
                                (N175)? btb_q[1165] : 
                                (N177)? btb_q[1230] : 
                                (N179)? btb_q[1295] : 
                                (N181)? btb_q[1360] : 
                                (N183)? btb_q[1425] : 
                                (N185)? btb_q[1490] : 
                                (N187)? btb_q[1555] : 
                                (N189)? btb_q[1620] : 
                                (N191)? btb_q[1685] : 
                                (N193)? btb_q[1750] : 
                                (N195)? btb_q[1815] : 
                                (N197)? btb_q[1880] : 
                                (N199)? btb_q[1945] : 
                                (N201)? btb_q[2010] : 
                                (N203)? btb_q[2075] : 
                                (N142)? btb_q[2140] : 
                                (N144)? btb_q[2205] : 
                                (N146)? btb_q[2270] : 
                                (N148)? btb_q[2335] : 
                                (N150)? btb_q[2400] : 
                                (N152)? btb_q[2465] : 
                                (N154)? btb_q[2530] : 
                                (N156)? btb_q[2595] : 
                                (N158)? btb_q[2660] : 
                                (N160)? btb_q[2725] : 
                                (N162)? btb_q[2790] : 
                                (N164)? btb_q[2855] : 
                                (N166)? btb_q[2920] : 
                                (N168)? btb_q[2985] : 
                                (N170)? btb_q[3050] : 
                                (N172)? btb_q[3115] : 
                                (N174)? btb_q[3180] : 
                                (N176)? btb_q[3245] : 
                                (N178)? btb_q[3310] : 
                                (N180)? btb_q[3375] : 
                                (N182)? btb_q[3440] : 
                                (N184)? btb_q[3505] : 
                                (N186)? btb_q[3570] : 
                                (N188)? btb_q[3635] : 
                                (N190)? btb_q[3700] : 
                                (N192)? btb_q[3765] : 
                                (N194)? btb_q[3830] : 
                                (N196)? btb_q[3895] : 
                                (N198)? btb_q[3960] : 
                                (N200)? btb_q[4025] : 
                                (N202)? btb_q[4090] : 
                                (N204)? btb_q[4155] : 1'b0;
  assign btb_prediction_o[59] = (N141)? btb_q[59] : 
                                (N143)? btb_q[124] : 
                                (N145)? btb_q[189] : 
                                (N147)? btb_q[254] : 
                                (N149)? btb_q[319] : 
                                (N151)? btb_q[384] : 
                                (N153)? btb_q[449] : 
                                (N155)? btb_q[514] : 
                                (N157)? btb_q[579] : 
                                (N159)? btb_q[644] : 
                                (N161)? btb_q[709] : 
                                (N163)? btb_q[774] : 
                                (N165)? btb_q[839] : 
                                (N167)? btb_q[904] : 
                                (N169)? btb_q[969] : 
                                (N171)? btb_q[1034] : 
                                (N173)? btb_q[1099] : 
                                (N175)? btb_q[1164] : 
                                (N177)? btb_q[1229] : 
                                (N179)? btb_q[1294] : 
                                (N181)? btb_q[1359] : 
                                (N183)? btb_q[1424] : 
                                (N185)? btb_q[1489] : 
                                (N187)? btb_q[1554] : 
                                (N189)? btb_q[1619] : 
                                (N191)? btb_q[1684] : 
                                (N193)? btb_q[1749] : 
                                (N195)? btb_q[1814] : 
                                (N197)? btb_q[1879] : 
                                (N199)? btb_q[1944] : 
                                (N201)? btb_q[2009] : 
                                (N203)? btb_q[2074] : 
                                (N142)? btb_q[2139] : 
                                (N144)? btb_q[2204] : 
                                (N146)? btb_q[2269] : 
                                (N148)? btb_q[2334] : 
                                (N150)? btb_q[2399] : 
                                (N152)? btb_q[2464] : 
                                (N154)? btb_q[2529] : 
                                (N156)? btb_q[2594] : 
                                (N158)? btb_q[2659] : 
                                (N160)? btb_q[2724] : 
                                (N162)? btb_q[2789] : 
                                (N164)? btb_q[2854] : 
                                (N166)? btb_q[2919] : 
                                (N168)? btb_q[2984] : 
                                (N170)? btb_q[3049] : 
                                (N172)? btb_q[3114] : 
                                (N174)? btb_q[3179] : 
                                (N176)? btb_q[3244] : 
                                (N178)? btb_q[3309] : 
                                (N180)? btb_q[3374] : 
                                (N182)? btb_q[3439] : 
                                (N184)? btb_q[3504] : 
                                (N186)? btb_q[3569] : 
                                (N188)? btb_q[3634] : 
                                (N190)? btb_q[3699] : 
                                (N192)? btb_q[3764] : 
                                (N194)? btb_q[3829] : 
                                (N196)? btb_q[3894] : 
                                (N198)? btb_q[3959] : 
                                (N200)? btb_q[4024] : 
                                (N202)? btb_q[4089] : 
                                (N204)? btb_q[4154] : 1'b0;
  assign btb_prediction_o[58] = (N141)? btb_q[58] : 
                                (N143)? btb_q[123] : 
                                (N145)? btb_q[188] : 
                                (N147)? btb_q[253] : 
                                (N149)? btb_q[318] : 
                                (N151)? btb_q[383] : 
                                (N153)? btb_q[448] : 
                                (N155)? btb_q[513] : 
                                (N157)? btb_q[578] : 
                                (N159)? btb_q[643] : 
                                (N161)? btb_q[708] : 
                                (N163)? btb_q[773] : 
                                (N165)? btb_q[838] : 
                                (N167)? btb_q[903] : 
                                (N169)? btb_q[968] : 
                                (N171)? btb_q[1033] : 
                                (N173)? btb_q[1098] : 
                                (N175)? btb_q[1163] : 
                                (N177)? btb_q[1228] : 
                                (N179)? btb_q[1293] : 
                                (N181)? btb_q[1358] : 
                                (N183)? btb_q[1423] : 
                                (N185)? btb_q[1488] : 
                                (N187)? btb_q[1553] : 
                                (N189)? btb_q[1618] : 
                                (N191)? btb_q[1683] : 
                                (N193)? btb_q[1748] : 
                                (N195)? btb_q[1813] : 
                                (N197)? btb_q[1878] : 
                                (N199)? btb_q[1943] : 
                                (N201)? btb_q[2008] : 
                                (N203)? btb_q[2073] : 
                                (N142)? btb_q[2138] : 
                                (N144)? btb_q[2203] : 
                                (N146)? btb_q[2268] : 
                                (N148)? btb_q[2333] : 
                                (N150)? btb_q[2398] : 
                                (N152)? btb_q[2463] : 
                                (N154)? btb_q[2528] : 
                                (N156)? btb_q[2593] : 
                                (N158)? btb_q[2658] : 
                                (N160)? btb_q[2723] : 
                                (N162)? btb_q[2788] : 
                                (N164)? btb_q[2853] : 
                                (N166)? btb_q[2918] : 
                                (N168)? btb_q[2983] : 
                                (N170)? btb_q[3048] : 
                                (N172)? btb_q[3113] : 
                                (N174)? btb_q[3178] : 
                                (N176)? btb_q[3243] : 
                                (N178)? btb_q[3308] : 
                                (N180)? btb_q[3373] : 
                                (N182)? btb_q[3438] : 
                                (N184)? btb_q[3503] : 
                                (N186)? btb_q[3568] : 
                                (N188)? btb_q[3633] : 
                                (N190)? btb_q[3698] : 
                                (N192)? btb_q[3763] : 
                                (N194)? btb_q[3828] : 
                                (N196)? btb_q[3893] : 
                                (N198)? btb_q[3958] : 
                                (N200)? btb_q[4023] : 
                                (N202)? btb_q[4088] : 
                                (N204)? btb_q[4153] : 1'b0;
  assign btb_prediction_o[57] = (N141)? btb_q[57] : 
                                (N143)? btb_q[122] : 
                                (N145)? btb_q[187] : 
                                (N147)? btb_q[252] : 
                                (N149)? btb_q[317] : 
                                (N151)? btb_q[382] : 
                                (N153)? btb_q[447] : 
                                (N155)? btb_q[512] : 
                                (N157)? btb_q[577] : 
                                (N159)? btb_q[642] : 
                                (N161)? btb_q[707] : 
                                (N163)? btb_q[772] : 
                                (N165)? btb_q[837] : 
                                (N167)? btb_q[902] : 
                                (N169)? btb_q[967] : 
                                (N171)? btb_q[1032] : 
                                (N173)? btb_q[1097] : 
                                (N175)? btb_q[1162] : 
                                (N177)? btb_q[1227] : 
                                (N179)? btb_q[1292] : 
                                (N181)? btb_q[1357] : 
                                (N183)? btb_q[1422] : 
                                (N185)? btb_q[1487] : 
                                (N187)? btb_q[1552] : 
                                (N189)? btb_q[1617] : 
                                (N191)? btb_q[1682] : 
                                (N193)? btb_q[1747] : 
                                (N195)? btb_q[1812] : 
                                (N197)? btb_q[1877] : 
                                (N199)? btb_q[1942] : 
                                (N201)? btb_q[2007] : 
                                (N203)? btb_q[2072] : 
                                (N142)? btb_q[2137] : 
                                (N144)? btb_q[2202] : 
                                (N146)? btb_q[2267] : 
                                (N148)? btb_q[2332] : 
                                (N150)? btb_q[2397] : 
                                (N152)? btb_q[2462] : 
                                (N154)? btb_q[2527] : 
                                (N156)? btb_q[2592] : 
                                (N158)? btb_q[2657] : 
                                (N160)? btb_q[2722] : 
                                (N162)? btb_q[2787] : 
                                (N164)? btb_q[2852] : 
                                (N166)? btb_q[2917] : 
                                (N168)? btb_q[2982] : 
                                (N170)? btb_q[3047] : 
                                (N172)? btb_q[3112] : 
                                (N174)? btb_q[3177] : 
                                (N176)? btb_q[3242] : 
                                (N178)? btb_q[3307] : 
                                (N180)? btb_q[3372] : 
                                (N182)? btb_q[3437] : 
                                (N184)? btb_q[3502] : 
                                (N186)? btb_q[3567] : 
                                (N188)? btb_q[3632] : 
                                (N190)? btb_q[3697] : 
                                (N192)? btb_q[3762] : 
                                (N194)? btb_q[3827] : 
                                (N196)? btb_q[3892] : 
                                (N198)? btb_q[3957] : 
                                (N200)? btb_q[4022] : 
                                (N202)? btb_q[4087] : 
                                (N204)? btb_q[4152] : 1'b0;
  assign btb_prediction_o[56] = (N141)? btb_q[56] : 
                                (N143)? btb_q[121] : 
                                (N145)? btb_q[186] : 
                                (N147)? btb_q[251] : 
                                (N149)? btb_q[316] : 
                                (N151)? btb_q[381] : 
                                (N153)? btb_q[446] : 
                                (N155)? btb_q[511] : 
                                (N157)? btb_q[576] : 
                                (N159)? btb_q[641] : 
                                (N161)? btb_q[706] : 
                                (N163)? btb_q[771] : 
                                (N165)? btb_q[836] : 
                                (N167)? btb_q[901] : 
                                (N169)? btb_q[966] : 
                                (N171)? btb_q[1031] : 
                                (N173)? btb_q[1096] : 
                                (N175)? btb_q[1161] : 
                                (N177)? btb_q[1226] : 
                                (N179)? btb_q[1291] : 
                                (N181)? btb_q[1356] : 
                                (N183)? btb_q[1421] : 
                                (N185)? btb_q[1486] : 
                                (N187)? btb_q[1551] : 
                                (N189)? btb_q[1616] : 
                                (N191)? btb_q[1681] : 
                                (N193)? btb_q[1746] : 
                                (N195)? btb_q[1811] : 
                                (N197)? btb_q[1876] : 
                                (N199)? btb_q[1941] : 
                                (N201)? btb_q[2006] : 
                                (N203)? btb_q[2071] : 
                                (N142)? btb_q[2136] : 
                                (N144)? btb_q[2201] : 
                                (N146)? btb_q[2266] : 
                                (N148)? btb_q[2331] : 
                                (N150)? btb_q[2396] : 
                                (N152)? btb_q[2461] : 
                                (N154)? btb_q[2526] : 
                                (N156)? btb_q[2591] : 
                                (N158)? btb_q[2656] : 
                                (N160)? btb_q[2721] : 
                                (N162)? btb_q[2786] : 
                                (N164)? btb_q[2851] : 
                                (N166)? btb_q[2916] : 
                                (N168)? btb_q[2981] : 
                                (N170)? btb_q[3046] : 
                                (N172)? btb_q[3111] : 
                                (N174)? btb_q[3176] : 
                                (N176)? btb_q[3241] : 
                                (N178)? btb_q[3306] : 
                                (N180)? btb_q[3371] : 
                                (N182)? btb_q[3436] : 
                                (N184)? btb_q[3501] : 
                                (N186)? btb_q[3566] : 
                                (N188)? btb_q[3631] : 
                                (N190)? btb_q[3696] : 
                                (N192)? btb_q[3761] : 
                                (N194)? btb_q[3826] : 
                                (N196)? btb_q[3891] : 
                                (N198)? btb_q[3956] : 
                                (N200)? btb_q[4021] : 
                                (N202)? btb_q[4086] : 
                                (N204)? btb_q[4151] : 1'b0;
  assign btb_prediction_o[55] = (N141)? btb_q[55] : 
                                (N143)? btb_q[120] : 
                                (N145)? btb_q[185] : 
                                (N147)? btb_q[250] : 
                                (N149)? btb_q[315] : 
                                (N151)? btb_q[380] : 
                                (N153)? btb_q[445] : 
                                (N155)? btb_q[510] : 
                                (N157)? btb_q[575] : 
                                (N159)? btb_q[640] : 
                                (N161)? btb_q[705] : 
                                (N163)? btb_q[770] : 
                                (N165)? btb_q[835] : 
                                (N167)? btb_q[900] : 
                                (N169)? btb_q[965] : 
                                (N171)? btb_q[1030] : 
                                (N173)? btb_q[1095] : 
                                (N175)? btb_q[1160] : 
                                (N177)? btb_q[1225] : 
                                (N179)? btb_q[1290] : 
                                (N181)? btb_q[1355] : 
                                (N183)? btb_q[1420] : 
                                (N185)? btb_q[1485] : 
                                (N187)? btb_q[1550] : 
                                (N189)? btb_q[1615] : 
                                (N191)? btb_q[1680] : 
                                (N193)? btb_q[1745] : 
                                (N195)? btb_q[1810] : 
                                (N197)? btb_q[1875] : 
                                (N199)? btb_q[1940] : 
                                (N201)? btb_q[2005] : 
                                (N203)? btb_q[2070] : 
                                (N142)? btb_q[2135] : 
                                (N144)? btb_q[2200] : 
                                (N146)? btb_q[2265] : 
                                (N148)? btb_q[2330] : 
                                (N150)? btb_q[2395] : 
                                (N152)? btb_q[2460] : 
                                (N154)? btb_q[2525] : 
                                (N156)? btb_q[2590] : 
                                (N158)? btb_q[2655] : 
                                (N160)? btb_q[2720] : 
                                (N162)? btb_q[2785] : 
                                (N164)? btb_q[2850] : 
                                (N166)? btb_q[2915] : 
                                (N168)? btb_q[2980] : 
                                (N170)? btb_q[3045] : 
                                (N172)? btb_q[3110] : 
                                (N174)? btb_q[3175] : 
                                (N176)? btb_q[3240] : 
                                (N178)? btb_q[3305] : 
                                (N180)? btb_q[3370] : 
                                (N182)? btb_q[3435] : 
                                (N184)? btb_q[3500] : 
                                (N186)? btb_q[3565] : 
                                (N188)? btb_q[3630] : 
                                (N190)? btb_q[3695] : 
                                (N192)? btb_q[3760] : 
                                (N194)? btb_q[3825] : 
                                (N196)? btb_q[3890] : 
                                (N198)? btb_q[3955] : 
                                (N200)? btb_q[4020] : 
                                (N202)? btb_q[4085] : 
                                (N204)? btb_q[4150] : 1'b0;
  assign btb_prediction_o[54] = (N141)? btb_q[54] : 
                                (N143)? btb_q[119] : 
                                (N145)? btb_q[184] : 
                                (N147)? btb_q[249] : 
                                (N149)? btb_q[314] : 
                                (N151)? btb_q[379] : 
                                (N153)? btb_q[444] : 
                                (N155)? btb_q[509] : 
                                (N157)? btb_q[574] : 
                                (N159)? btb_q[639] : 
                                (N161)? btb_q[704] : 
                                (N163)? btb_q[769] : 
                                (N165)? btb_q[834] : 
                                (N167)? btb_q[899] : 
                                (N169)? btb_q[964] : 
                                (N171)? btb_q[1029] : 
                                (N173)? btb_q[1094] : 
                                (N175)? btb_q[1159] : 
                                (N177)? btb_q[1224] : 
                                (N179)? btb_q[1289] : 
                                (N181)? btb_q[1354] : 
                                (N183)? btb_q[1419] : 
                                (N185)? btb_q[1484] : 
                                (N187)? btb_q[1549] : 
                                (N189)? btb_q[1614] : 
                                (N191)? btb_q[1679] : 
                                (N193)? btb_q[1744] : 
                                (N195)? btb_q[1809] : 
                                (N197)? btb_q[1874] : 
                                (N199)? btb_q[1939] : 
                                (N201)? btb_q[2004] : 
                                (N203)? btb_q[2069] : 
                                (N142)? btb_q[2134] : 
                                (N144)? btb_q[2199] : 
                                (N146)? btb_q[2264] : 
                                (N148)? btb_q[2329] : 
                                (N150)? btb_q[2394] : 
                                (N152)? btb_q[2459] : 
                                (N154)? btb_q[2524] : 
                                (N156)? btb_q[2589] : 
                                (N158)? btb_q[2654] : 
                                (N160)? btb_q[2719] : 
                                (N162)? btb_q[2784] : 
                                (N164)? btb_q[2849] : 
                                (N166)? btb_q[2914] : 
                                (N168)? btb_q[2979] : 
                                (N170)? btb_q[3044] : 
                                (N172)? btb_q[3109] : 
                                (N174)? btb_q[3174] : 
                                (N176)? btb_q[3239] : 
                                (N178)? btb_q[3304] : 
                                (N180)? btb_q[3369] : 
                                (N182)? btb_q[3434] : 
                                (N184)? btb_q[3499] : 
                                (N186)? btb_q[3564] : 
                                (N188)? btb_q[3629] : 
                                (N190)? btb_q[3694] : 
                                (N192)? btb_q[3759] : 
                                (N194)? btb_q[3824] : 
                                (N196)? btb_q[3889] : 
                                (N198)? btb_q[3954] : 
                                (N200)? btb_q[4019] : 
                                (N202)? btb_q[4084] : 
                                (N204)? btb_q[4149] : 1'b0;
  assign btb_prediction_o[53] = (N141)? btb_q[53] : 
                                (N143)? btb_q[118] : 
                                (N145)? btb_q[183] : 
                                (N147)? btb_q[248] : 
                                (N149)? btb_q[313] : 
                                (N151)? btb_q[378] : 
                                (N153)? btb_q[443] : 
                                (N155)? btb_q[508] : 
                                (N157)? btb_q[573] : 
                                (N159)? btb_q[638] : 
                                (N161)? btb_q[703] : 
                                (N163)? btb_q[768] : 
                                (N165)? btb_q[833] : 
                                (N167)? btb_q[898] : 
                                (N169)? btb_q[963] : 
                                (N171)? btb_q[1028] : 
                                (N173)? btb_q[1093] : 
                                (N175)? btb_q[1158] : 
                                (N177)? btb_q[1223] : 
                                (N179)? btb_q[1288] : 
                                (N181)? btb_q[1353] : 
                                (N183)? btb_q[1418] : 
                                (N185)? btb_q[1483] : 
                                (N187)? btb_q[1548] : 
                                (N189)? btb_q[1613] : 
                                (N191)? btb_q[1678] : 
                                (N193)? btb_q[1743] : 
                                (N195)? btb_q[1808] : 
                                (N197)? btb_q[1873] : 
                                (N199)? btb_q[1938] : 
                                (N201)? btb_q[2003] : 
                                (N203)? btb_q[2068] : 
                                (N142)? btb_q[2133] : 
                                (N144)? btb_q[2198] : 
                                (N146)? btb_q[2263] : 
                                (N148)? btb_q[2328] : 
                                (N150)? btb_q[2393] : 
                                (N152)? btb_q[2458] : 
                                (N154)? btb_q[2523] : 
                                (N156)? btb_q[2588] : 
                                (N158)? btb_q[2653] : 
                                (N160)? btb_q[2718] : 
                                (N162)? btb_q[2783] : 
                                (N164)? btb_q[2848] : 
                                (N166)? btb_q[2913] : 
                                (N168)? btb_q[2978] : 
                                (N170)? btb_q[3043] : 
                                (N172)? btb_q[3108] : 
                                (N174)? btb_q[3173] : 
                                (N176)? btb_q[3238] : 
                                (N178)? btb_q[3303] : 
                                (N180)? btb_q[3368] : 
                                (N182)? btb_q[3433] : 
                                (N184)? btb_q[3498] : 
                                (N186)? btb_q[3563] : 
                                (N188)? btb_q[3628] : 
                                (N190)? btb_q[3693] : 
                                (N192)? btb_q[3758] : 
                                (N194)? btb_q[3823] : 
                                (N196)? btb_q[3888] : 
                                (N198)? btb_q[3953] : 
                                (N200)? btb_q[4018] : 
                                (N202)? btb_q[4083] : 
                                (N204)? btb_q[4148] : 1'b0;
  assign btb_prediction_o[52] = (N141)? btb_q[52] : 
                                (N143)? btb_q[117] : 
                                (N145)? btb_q[182] : 
                                (N147)? btb_q[247] : 
                                (N149)? btb_q[312] : 
                                (N151)? btb_q[377] : 
                                (N153)? btb_q[442] : 
                                (N155)? btb_q[507] : 
                                (N157)? btb_q[572] : 
                                (N159)? btb_q[637] : 
                                (N161)? btb_q[702] : 
                                (N163)? btb_q[767] : 
                                (N165)? btb_q[832] : 
                                (N167)? btb_q[897] : 
                                (N169)? btb_q[962] : 
                                (N171)? btb_q[1027] : 
                                (N173)? btb_q[1092] : 
                                (N175)? btb_q[1157] : 
                                (N177)? btb_q[1222] : 
                                (N179)? btb_q[1287] : 
                                (N181)? btb_q[1352] : 
                                (N183)? btb_q[1417] : 
                                (N185)? btb_q[1482] : 
                                (N187)? btb_q[1547] : 
                                (N189)? btb_q[1612] : 
                                (N191)? btb_q[1677] : 
                                (N193)? btb_q[1742] : 
                                (N195)? btb_q[1807] : 
                                (N197)? btb_q[1872] : 
                                (N199)? btb_q[1937] : 
                                (N201)? btb_q[2002] : 
                                (N203)? btb_q[2067] : 
                                (N142)? btb_q[2132] : 
                                (N144)? btb_q[2197] : 
                                (N146)? btb_q[2262] : 
                                (N148)? btb_q[2327] : 
                                (N150)? btb_q[2392] : 
                                (N152)? btb_q[2457] : 
                                (N154)? btb_q[2522] : 
                                (N156)? btb_q[2587] : 
                                (N158)? btb_q[2652] : 
                                (N160)? btb_q[2717] : 
                                (N162)? btb_q[2782] : 
                                (N164)? btb_q[2847] : 
                                (N166)? btb_q[2912] : 
                                (N168)? btb_q[2977] : 
                                (N170)? btb_q[3042] : 
                                (N172)? btb_q[3107] : 
                                (N174)? btb_q[3172] : 
                                (N176)? btb_q[3237] : 
                                (N178)? btb_q[3302] : 
                                (N180)? btb_q[3367] : 
                                (N182)? btb_q[3432] : 
                                (N184)? btb_q[3497] : 
                                (N186)? btb_q[3562] : 
                                (N188)? btb_q[3627] : 
                                (N190)? btb_q[3692] : 
                                (N192)? btb_q[3757] : 
                                (N194)? btb_q[3822] : 
                                (N196)? btb_q[3887] : 
                                (N198)? btb_q[3952] : 
                                (N200)? btb_q[4017] : 
                                (N202)? btb_q[4082] : 
                                (N204)? btb_q[4147] : 1'b0;
  assign btb_prediction_o[51] = (N141)? btb_q[51] : 
                                (N143)? btb_q[116] : 
                                (N145)? btb_q[181] : 
                                (N147)? btb_q[246] : 
                                (N149)? btb_q[311] : 
                                (N151)? btb_q[376] : 
                                (N153)? btb_q[441] : 
                                (N155)? btb_q[506] : 
                                (N157)? btb_q[571] : 
                                (N159)? btb_q[636] : 
                                (N161)? btb_q[701] : 
                                (N163)? btb_q[766] : 
                                (N165)? btb_q[831] : 
                                (N167)? btb_q[896] : 
                                (N169)? btb_q[961] : 
                                (N171)? btb_q[1026] : 
                                (N173)? btb_q[1091] : 
                                (N175)? btb_q[1156] : 
                                (N177)? btb_q[1221] : 
                                (N179)? btb_q[1286] : 
                                (N181)? btb_q[1351] : 
                                (N183)? btb_q[1416] : 
                                (N185)? btb_q[1481] : 
                                (N187)? btb_q[1546] : 
                                (N189)? btb_q[1611] : 
                                (N191)? btb_q[1676] : 
                                (N193)? btb_q[1741] : 
                                (N195)? btb_q[1806] : 
                                (N197)? btb_q[1871] : 
                                (N199)? btb_q[1936] : 
                                (N201)? btb_q[2001] : 
                                (N203)? btb_q[2066] : 
                                (N142)? btb_q[2131] : 
                                (N144)? btb_q[2196] : 
                                (N146)? btb_q[2261] : 
                                (N148)? btb_q[2326] : 
                                (N150)? btb_q[2391] : 
                                (N152)? btb_q[2456] : 
                                (N154)? btb_q[2521] : 
                                (N156)? btb_q[2586] : 
                                (N158)? btb_q[2651] : 
                                (N160)? btb_q[2716] : 
                                (N162)? btb_q[2781] : 
                                (N164)? btb_q[2846] : 
                                (N166)? btb_q[2911] : 
                                (N168)? btb_q[2976] : 
                                (N170)? btb_q[3041] : 
                                (N172)? btb_q[3106] : 
                                (N174)? btb_q[3171] : 
                                (N176)? btb_q[3236] : 
                                (N178)? btb_q[3301] : 
                                (N180)? btb_q[3366] : 
                                (N182)? btb_q[3431] : 
                                (N184)? btb_q[3496] : 
                                (N186)? btb_q[3561] : 
                                (N188)? btb_q[3626] : 
                                (N190)? btb_q[3691] : 
                                (N192)? btb_q[3756] : 
                                (N194)? btb_q[3821] : 
                                (N196)? btb_q[3886] : 
                                (N198)? btb_q[3951] : 
                                (N200)? btb_q[4016] : 
                                (N202)? btb_q[4081] : 
                                (N204)? btb_q[4146] : 1'b0;
  assign btb_prediction_o[50] = (N141)? btb_q[50] : 
                                (N143)? btb_q[115] : 
                                (N145)? btb_q[180] : 
                                (N147)? btb_q[245] : 
                                (N149)? btb_q[310] : 
                                (N151)? btb_q[375] : 
                                (N153)? btb_q[440] : 
                                (N155)? btb_q[505] : 
                                (N157)? btb_q[570] : 
                                (N159)? btb_q[635] : 
                                (N161)? btb_q[700] : 
                                (N163)? btb_q[765] : 
                                (N165)? btb_q[830] : 
                                (N167)? btb_q[895] : 
                                (N169)? btb_q[960] : 
                                (N171)? btb_q[1025] : 
                                (N173)? btb_q[1090] : 
                                (N175)? btb_q[1155] : 
                                (N177)? btb_q[1220] : 
                                (N179)? btb_q[1285] : 
                                (N181)? btb_q[1350] : 
                                (N183)? btb_q[1415] : 
                                (N185)? btb_q[1480] : 
                                (N187)? btb_q[1545] : 
                                (N189)? btb_q[1610] : 
                                (N191)? btb_q[1675] : 
                                (N193)? btb_q[1740] : 
                                (N195)? btb_q[1805] : 
                                (N197)? btb_q[1870] : 
                                (N199)? btb_q[1935] : 
                                (N201)? btb_q[2000] : 
                                (N203)? btb_q[2065] : 
                                (N142)? btb_q[2130] : 
                                (N144)? btb_q[2195] : 
                                (N146)? btb_q[2260] : 
                                (N148)? btb_q[2325] : 
                                (N150)? btb_q[2390] : 
                                (N152)? btb_q[2455] : 
                                (N154)? btb_q[2520] : 
                                (N156)? btb_q[2585] : 
                                (N158)? btb_q[2650] : 
                                (N160)? btb_q[2715] : 
                                (N162)? btb_q[2780] : 
                                (N164)? btb_q[2845] : 
                                (N166)? btb_q[2910] : 
                                (N168)? btb_q[2975] : 
                                (N170)? btb_q[3040] : 
                                (N172)? btb_q[3105] : 
                                (N174)? btb_q[3170] : 
                                (N176)? btb_q[3235] : 
                                (N178)? btb_q[3300] : 
                                (N180)? btb_q[3365] : 
                                (N182)? btb_q[3430] : 
                                (N184)? btb_q[3495] : 
                                (N186)? btb_q[3560] : 
                                (N188)? btb_q[3625] : 
                                (N190)? btb_q[3690] : 
                                (N192)? btb_q[3755] : 
                                (N194)? btb_q[3820] : 
                                (N196)? btb_q[3885] : 
                                (N198)? btb_q[3950] : 
                                (N200)? btb_q[4015] : 
                                (N202)? btb_q[4080] : 
                                (N204)? btb_q[4145] : 1'b0;
  assign btb_prediction_o[49] = (N141)? btb_q[49] : 
                                (N143)? btb_q[114] : 
                                (N145)? btb_q[179] : 
                                (N147)? btb_q[244] : 
                                (N149)? btb_q[309] : 
                                (N151)? btb_q[374] : 
                                (N153)? btb_q[439] : 
                                (N155)? btb_q[504] : 
                                (N157)? btb_q[569] : 
                                (N159)? btb_q[634] : 
                                (N161)? btb_q[699] : 
                                (N163)? btb_q[764] : 
                                (N165)? btb_q[829] : 
                                (N167)? btb_q[894] : 
                                (N169)? btb_q[959] : 
                                (N171)? btb_q[1024] : 
                                (N173)? btb_q[1089] : 
                                (N175)? btb_q[1154] : 
                                (N177)? btb_q[1219] : 
                                (N179)? btb_q[1284] : 
                                (N181)? btb_q[1349] : 
                                (N183)? btb_q[1414] : 
                                (N185)? btb_q[1479] : 
                                (N187)? btb_q[1544] : 
                                (N189)? btb_q[1609] : 
                                (N191)? btb_q[1674] : 
                                (N193)? btb_q[1739] : 
                                (N195)? btb_q[1804] : 
                                (N197)? btb_q[1869] : 
                                (N199)? btb_q[1934] : 
                                (N201)? btb_q[1999] : 
                                (N203)? btb_q[2064] : 
                                (N142)? btb_q[2129] : 
                                (N144)? btb_q[2194] : 
                                (N146)? btb_q[2259] : 
                                (N148)? btb_q[2324] : 
                                (N150)? btb_q[2389] : 
                                (N152)? btb_q[2454] : 
                                (N154)? btb_q[2519] : 
                                (N156)? btb_q[2584] : 
                                (N158)? btb_q[2649] : 
                                (N160)? btb_q[2714] : 
                                (N162)? btb_q[2779] : 
                                (N164)? btb_q[2844] : 
                                (N166)? btb_q[2909] : 
                                (N168)? btb_q[2974] : 
                                (N170)? btb_q[3039] : 
                                (N172)? btb_q[3104] : 
                                (N174)? btb_q[3169] : 
                                (N176)? btb_q[3234] : 
                                (N178)? btb_q[3299] : 
                                (N180)? btb_q[3364] : 
                                (N182)? btb_q[3429] : 
                                (N184)? btb_q[3494] : 
                                (N186)? btb_q[3559] : 
                                (N188)? btb_q[3624] : 
                                (N190)? btb_q[3689] : 
                                (N192)? btb_q[3754] : 
                                (N194)? btb_q[3819] : 
                                (N196)? btb_q[3884] : 
                                (N198)? btb_q[3949] : 
                                (N200)? btb_q[4014] : 
                                (N202)? btb_q[4079] : 
                                (N204)? btb_q[4144] : 1'b0;
  assign btb_prediction_o[48] = (N141)? btb_q[48] : 
                                (N143)? btb_q[113] : 
                                (N145)? btb_q[178] : 
                                (N147)? btb_q[243] : 
                                (N149)? btb_q[308] : 
                                (N151)? btb_q[373] : 
                                (N153)? btb_q[438] : 
                                (N155)? btb_q[503] : 
                                (N157)? btb_q[568] : 
                                (N159)? btb_q[633] : 
                                (N161)? btb_q[698] : 
                                (N163)? btb_q[763] : 
                                (N165)? btb_q[828] : 
                                (N167)? btb_q[893] : 
                                (N169)? btb_q[958] : 
                                (N171)? btb_q[1023] : 
                                (N173)? btb_q[1088] : 
                                (N175)? btb_q[1153] : 
                                (N177)? btb_q[1218] : 
                                (N179)? btb_q[1283] : 
                                (N181)? btb_q[1348] : 
                                (N183)? btb_q[1413] : 
                                (N185)? btb_q[1478] : 
                                (N187)? btb_q[1543] : 
                                (N189)? btb_q[1608] : 
                                (N191)? btb_q[1673] : 
                                (N193)? btb_q[1738] : 
                                (N195)? btb_q[1803] : 
                                (N197)? btb_q[1868] : 
                                (N199)? btb_q[1933] : 
                                (N201)? btb_q[1998] : 
                                (N203)? btb_q[2063] : 
                                (N142)? btb_q[2128] : 
                                (N144)? btb_q[2193] : 
                                (N146)? btb_q[2258] : 
                                (N148)? btb_q[2323] : 
                                (N150)? btb_q[2388] : 
                                (N152)? btb_q[2453] : 
                                (N154)? btb_q[2518] : 
                                (N156)? btb_q[2583] : 
                                (N158)? btb_q[2648] : 
                                (N160)? btb_q[2713] : 
                                (N162)? btb_q[2778] : 
                                (N164)? btb_q[2843] : 
                                (N166)? btb_q[2908] : 
                                (N168)? btb_q[2973] : 
                                (N170)? btb_q[3038] : 
                                (N172)? btb_q[3103] : 
                                (N174)? btb_q[3168] : 
                                (N176)? btb_q[3233] : 
                                (N178)? btb_q[3298] : 
                                (N180)? btb_q[3363] : 
                                (N182)? btb_q[3428] : 
                                (N184)? btb_q[3493] : 
                                (N186)? btb_q[3558] : 
                                (N188)? btb_q[3623] : 
                                (N190)? btb_q[3688] : 
                                (N192)? btb_q[3753] : 
                                (N194)? btb_q[3818] : 
                                (N196)? btb_q[3883] : 
                                (N198)? btb_q[3948] : 
                                (N200)? btb_q[4013] : 
                                (N202)? btb_q[4078] : 
                                (N204)? btb_q[4143] : 1'b0;
  assign btb_prediction_o[47] = (N141)? btb_q[47] : 
                                (N143)? btb_q[112] : 
                                (N145)? btb_q[177] : 
                                (N147)? btb_q[242] : 
                                (N149)? btb_q[307] : 
                                (N151)? btb_q[372] : 
                                (N153)? btb_q[437] : 
                                (N155)? btb_q[502] : 
                                (N157)? btb_q[567] : 
                                (N159)? btb_q[632] : 
                                (N161)? btb_q[697] : 
                                (N163)? btb_q[762] : 
                                (N165)? btb_q[827] : 
                                (N167)? btb_q[892] : 
                                (N169)? btb_q[957] : 
                                (N171)? btb_q[1022] : 
                                (N173)? btb_q[1087] : 
                                (N175)? btb_q[1152] : 
                                (N177)? btb_q[1217] : 
                                (N179)? btb_q[1282] : 
                                (N181)? btb_q[1347] : 
                                (N183)? btb_q[1412] : 
                                (N185)? btb_q[1477] : 
                                (N187)? btb_q[1542] : 
                                (N189)? btb_q[1607] : 
                                (N191)? btb_q[1672] : 
                                (N193)? btb_q[1737] : 
                                (N195)? btb_q[1802] : 
                                (N197)? btb_q[1867] : 
                                (N199)? btb_q[1932] : 
                                (N201)? btb_q[1997] : 
                                (N203)? btb_q[2062] : 
                                (N142)? btb_q[2127] : 
                                (N144)? btb_q[2192] : 
                                (N146)? btb_q[2257] : 
                                (N148)? btb_q[2322] : 
                                (N150)? btb_q[2387] : 
                                (N152)? btb_q[2452] : 
                                (N154)? btb_q[2517] : 
                                (N156)? btb_q[2582] : 
                                (N158)? btb_q[2647] : 
                                (N160)? btb_q[2712] : 
                                (N162)? btb_q[2777] : 
                                (N164)? btb_q[2842] : 
                                (N166)? btb_q[2907] : 
                                (N168)? btb_q[2972] : 
                                (N170)? btb_q[3037] : 
                                (N172)? btb_q[3102] : 
                                (N174)? btb_q[3167] : 
                                (N176)? btb_q[3232] : 
                                (N178)? btb_q[3297] : 
                                (N180)? btb_q[3362] : 
                                (N182)? btb_q[3427] : 
                                (N184)? btb_q[3492] : 
                                (N186)? btb_q[3557] : 
                                (N188)? btb_q[3622] : 
                                (N190)? btb_q[3687] : 
                                (N192)? btb_q[3752] : 
                                (N194)? btb_q[3817] : 
                                (N196)? btb_q[3882] : 
                                (N198)? btb_q[3947] : 
                                (N200)? btb_q[4012] : 
                                (N202)? btb_q[4077] : 
                                (N204)? btb_q[4142] : 1'b0;
  assign btb_prediction_o[46] = (N141)? btb_q[46] : 
                                (N143)? btb_q[111] : 
                                (N145)? btb_q[176] : 
                                (N147)? btb_q[241] : 
                                (N149)? btb_q[306] : 
                                (N151)? btb_q[371] : 
                                (N153)? btb_q[436] : 
                                (N155)? btb_q[501] : 
                                (N157)? btb_q[566] : 
                                (N159)? btb_q[631] : 
                                (N161)? btb_q[696] : 
                                (N163)? btb_q[761] : 
                                (N165)? btb_q[826] : 
                                (N167)? btb_q[891] : 
                                (N169)? btb_q[956] : 
                                (N171)? btb_q[1021] : 
                                (N173)? btb_q[1086] : 
                                (N175)? btb_q[1151] : 
                                (N177)? btb_q[1216] : 
                                (N179)? btb_q[1281] : 
                                (N181)? btb_q[1346] : 
                                (N183)? btb_q[1411] : 
                                (N185)? btb_q[1476] : 
                                (N187)? btb_q[1541] : 
                                (N189)? btb_q[1606] : 
                                (N191)? btb_q[1671] : 
                                (N193)? btb_q[1736] : 
                                (N195)? btb_q[1801] : 
                                (N197)? btb_q[1866] : 
                                (N199)? btb_q[1931] : 
                                (N201)? btb_q[1996] : 
                                (N203)? btb_q[2061] : 
                                (N142)? btb_q[2126] : 
                                (N144)? btb_q[2191] : 
                                (N146)? btb_q[2256] : 
                                (N148)? btb_q[2321] : 
                                (N150)? btb_q[2386] : 
                                (N152)? btb_q[2451] : 
                                (N154)? btb_q[2516] : 
                                (N156)? btb_q[2581] : 
                                (N158)? btb_q[2646] : 
                                (N160)? btb_q[2711] : 
                                (N162)? btb_q[2776] : 
                                (N164)? btb_q[2841] : 
                                (N166)? btb_q[2906] : 
                                (N168)? btb_q[2971] : 
                                (N170)? btb_q[3036] : 
                                (N172)? btb_q[3101] : 
                                (N174)? btb_q[3166] : 
                                (N176)? btb_q[3231] : 
                                (N178)? btb_q[3296] : 
                                (N180)? btb_q[3361] : 
                                (N182)? btb_q[3426] : 
                                (N184)? btb_q[3491] : 
                                (N186)? btb_q[3556] : 
                                (N188)? btb_q[3621] : 
                                (N190)? btb_q[3686] : 
                                (N192)? btb_q[3751] : 
                                (N194)? btb_q[3816] : 
                                (N196)? btb_q[3881] : 
                                (N198)? btb_q[3946] : 
                                (N200)? btb_q[4011] : 
                                (N202)? btb_q[4076] : 
                                (N204)? btb_q[4141] : 1'b0;
  assign btb_prediction_o[45] = (N141)? btb_q[45] : 
                                (N143)? btb_q[110] : 
                                (N145)? btb_q[175] : 
                                (N147)? btb_q[240] : 
                                (N149)? btb_q[305] : 
                                (N151)? btb_q[370] : 
                                (N153)? btb_q[435] : 
                                (N155)? btb_q[500] : 
                                (N157)? btb_q[565] : 
                                (N159)? btb_q[630] : 
                                (N161)? btb_q[695] : 
                                (N163)? btb_q[760] : 
                                (N165)? btb_q[825] : 
                                (N167)? btb_q[890] : 
                                (N169)? btb_q[955] : 
                                (N171)? btb_q[1020] : 
                                (N173)? btb_q[1085] : 
                                (N175)? btb_q[1150] : 
                                (N177)? btb_q[1215] : 
                                (N179)? btb_q[1280] : 
                                (N181)? btb_q[1345] : 
                                (N183)? btb_q[1410] : 
                                (N185)? btb_q[1475] : 
                                (N187)? btb_q[1540] : 
                                (N189)? btb_q[1605] : 
                                (N191)? btb_q[1670] : 
                                (N193)? btb_q[1735] : 
                                (N195)? btb_q[1800] : 
                                (N197)? btb_q[1865] : 
                                (N199)? btb_q[1930] : 
                                (N201)? btb_q[1995] : 
                                (N203)? btb_q[2060] : 
                                (N142)? btb_q[2125] : 
                                (N144)? btb_q[2190] : 
                                (N146)? btb_q[2255] : 
                                (N148)? btb_q[2320] : 
                                (N150)? btb_q[2385] : 
                                (N152)? btb_q[2450] : 
                                (N154)? btb_q[2515] : 
                                (N156)? btb_q[2580] : 
                                (N158)? btb_q[2645] : 
                                (N160)? btb_q[2710] : 
                                (N162)? btb_q[2775] : 
                                (N164)? btb_q[2840] : 
                                (N166)? btb_q[2905] : 
                                (N168)? btb_q[2970] : 
                                (N170)? btb_q[3035] : 
                                (N172)? btb_q[3100] : 
                                (N174)? btb_q[3165] : 
                                (N176)? btb_q[3230] : 
                                (N178)? btb_q[3295] : 
                                (N180)? btb_q[3360] : 
                                (N182)? btb_q[3425] : 
                                (N184)? btb_q[3490] : 
                                (N186)? btb_q[3555] : 
                                (N188)? btb_q[3620] : 
                                (N190)? btb_q[3685] : 
                                (N192)? btb_q[3750] : 
                                (N194)? btb_q[3815] : 
                                (N196)? btb_q[3880] : 
                                (N198)? btb_q[3945] : 
                                (N200)? btb_q[4010] : 
                                (N202)? btb_q[4075] : 
                                (N204)? btb_q[4140] : 1'b0;
  assign btb_prediction_o[44] = (N141)? btb_q[44] : 
                                (N143)? btb_q[109] : 
                                (N145)? btb_q[174] : 
                                (N147)? btb_q[239] : 
                                (N149)? btb_q[304] : 
                                (N151)? btb_q[369] : 
                                (N153)? btb_q[434] : 
                                (N155)? btb_q[499] : 
                                (N157)? btb_q[564] : 
                                (N159)? btb_q[629] : 
                                (N161)? btb_q[694] : 
                                (N163)? btb_q[759] : 
                                (N165)? btb_q[824] : 
                                (N167)? btb_q[889] : 
                                (N169)? btb_q[954] : 
                                (N171)? btb_q[1019] : 
                                (N173)? btb_q[1084] : 
                                (N175)? btb_q[1149] : 
                                (N177)? btb_q[1214] : 
                                (N179)? btb_q[1279] : 
                                (N181)? btb_q[1344] : 
                                (N183)? btb_q[1409] : 
                                (N185)? btb_q[1474] : 
                                (N187)? btb_q[1539] : 
                                (N189)? btb_q[1604] : 
                                (N191)? btb_q[1669] : 
                                (N193)? btb_q[1734] : 
                                (N195)? btb_q[1799] : 
                                (N197)? btb_q[1864] : 
                                (N199)? btb_q[1929] : 
                                (N201)? btb_q[1994] : 
                                (N203)? btb_q[2059] : 
                                (N142)? btb_q[2124] : 
                                (N144)? btb_q[2189] : 
                                (N146)? btb_q[2254] : 
                                (N148)? btb_q[2319] : 
                                (N150)? btb_q[2384] : 
                                (N152)? btb_q[2449] : 
                                (N154)? btb_q[2514] : 
                                (N156)? btb_q[2579] : 
                                (N158)? btb_q[2644] : 
                                (N160)? btb_q[2709] : 
                                (N162)? btb_q[2774] : 
                                (N164)? btb_q[2839] : 
                                (N166)? btb_q[2904] : 
                                (N168)? btb_q[2969] : 
                                (N170)? btb_q[3034] : 
                                (N172)? btb_q[3099] : 
                                (N174)? btb_q[3164] : 
                                (N176)? btb_q[3229] : 
                                (N178)? btb_q[3294] : 
                                (N180)? btb_q[3359] : 
                                (N182)? btb_q[3424] : 
                                (N184)? btb_q[3489] : 
                                (N186)? btb_q[3554] : 
                                (N188)? btb_q[3619] : 
                                (N190)? btb_q[3684] : 
                                (N192)? btb_q[3749] : 
                                (N194)? btb_q[3814] : 
                                (N196)? btb_q[3879] : 
                                (N198)? btb_q[3944] : 
                                (N200)? btb_q[4009] : 
                                (N202)? btb_q[4074] : 
                                (N204)? btb_q[4139] : 1'b0;
  assign btb_prediction_o[43] = (N141)? btb_q[43] : 
                                (N143)? btb_q[108] : 
                                (N145)? btb_q[173] : 
                                (N147)? btb_q[238] : 
                                (N149)? btb_q[303] : 
                                (N151)? btb_q[368] : 
                                (N153)? btb_q[433] : 
                                (N155)? btb_q[498] : 
                                (N157)? btb_q[563] : 
                                (N159)? btb_q[628] : 
                                (N161)? btb_q[693] : 
                                (N163)? btb_q[758] : 
                                (N165)? btb_q[823] : 
                                (N167)? btb_q[888] : 
                                (N169)? btb_q[953] : 
                                (N171)? btb_q[1018] : 
                                (N173)? btb_q[1083] : 
                                (N175)? btb_q[1148] : 
                                (N177)? btb_q[1213] : 
                                (N179)? btb_q[1278] : 
                                (N181)? btb_q[1343] : 
                                (N183)? btb_q[1408] : 
                                (N185)? btb_q[1473] : 
                                (N187)? btb_q[1538] : 
                                (N189)? btb_q[1603] : 
                                (N191)? btb_q[1668] : 
                                (N193)? btb_q[1733] : 
                                (N195)? btb_q[1798] : 
                                (N197)? btb_q[1863] : 
                                (N199)? btb_q[1928] : 
                                (N201)? btb_q[1993] : 
                                (N203)? btb_q[2058] : 
                                (N142)? btb_q[2123] : 
                                (N144)? btb_q[2188] : 
                                (N146)? btb_q[2253] : 
                                (N148)? btb_q[2318] : 
                                (N150)? btb_q[2383] : 
                                (N152)? btb_q[2448] : 
                                (N154)? btb_q[2513] : 
                                (N156)? btb_q[2578] : 
                                (N158)? btb_q[2643] : 
                                (N160)? btb_q[2708] : 
                                (N162)? btb_q[2773] : 
                                (N164)? btb_q[2838] : 
                                (N166)? btb_q[2903] : 
                                (N168)? btb_q[2968] : 
                                (N170)? btb_q[3033] : 
                                (N172)? btb_q[3098] : 
                                (N174)? btb_q[3163] : 
                                (N176)? btb_q[3228] : 
                                (N178)? btb_q[3293] : 
                                (N180)? btb_q[3358] : 
                                (N182)? btb_q[3423] : 
                                (N184)? btb_q[3488] : 
                                (N186)? btb_q[3553] : 
                                (N188)? btb_q[3618] : 
                                (N190)? btb_q[3683] : 
                                (N192)? btb_q[3748] : 
                                (N194)? btb_q[3813] : 
                                (N196)? btb_q[3878] : 
                                (N198)? btb_q[3943] : 
                                (N200)? btb_q[4008] : 
                                (N202)? btb_q[4073] : 
                                (N204)? btb_q[4138] : 1'b0;
  assign btb_prediction_o[42] = (N141)? btb_q[42] : 
                                (N143)? btb_q[107] : 
                                (N145)? btb_q[172] : 
                                (N147)? btb_q[237] : 
                                (N149)? btb_q[302] : 
                                (N151)? btb_q[367] : 
                                (N153)? btb_q[432] : 
                                (N155)? btb_q[497] : 
                                (N157)? btb_q[562] : 
                                (N159)? btb_q[627] : 
                                (N161)? btb_q[692] : 
                                (N163)? btb_q[757] : 
                                (N165)? btb_q[822] : 
                                (N167)? btb_q[887] : 
                                (N169)? btb_q[952] : 
                                (N171)? btb_q[1017] : 
                                (N173)? btb_q[1082] : 
                                (N175)? btb_q[1147] : 
                                (N177)? btb_q[1212] : 
                                (N179)? btb_q[1277] : 
                                (N181)? btb_q[1342] : 
                                (N183)? btb_q[1407] : 
                                (N185)? btb_q[1472] : 
                                (N187)? btb_q[1537] : 
                                (N189)? btb_q[1602] : 
                                (N191)? btb_q[1667] : 
                                (N193)? btb_q[1732] : 
                                (N195)? btb_q[1797] : 
                                (N197)? btb_q[1862] : 
                                (N199)? btb_q[1927] : 
                                (N201)? btb_q[1992] : 
                                (N203)? btb_q[2057] : 
                                (N142)? btb_q[2122] : 
                                (N144)? btb_q[2187] : 
                                (N146)? btb_q[2252] : 
                                (N148)? btb_q[2317] : 
                                (N150)? btb_q[2382] : 
                                (N152)? btb_q[2447] : 
                                (N154)? btb_q[2512] : 
                                (N156)? btb_q[2577] : 
                                (N158)? btb_q[2642] : 
                                (N160)? btb_q[2707] : 
                                (N162)? btb_q[2772] : 
                                (N164)? btb_q[2837] : 
                                (N166)? btb_q[2902] : 
                                (N168)? btb_q[2967] : 
                                (N170)? btb_q[3032] : 
                                (N172)? btb_q[3097] : 
                                (N174)? btb_q[3162] : 
                                (N176)? btb_q[3227] : 
                                (N178)? btb_q[3292] : 
                                (N180)? btb_q[3357] : 
                                (N182)? btb_q[3422] : 
                                (N184)? btb_q[3487] : 
                                (N186)? btb_q[3552] : 
                                (N188)? btb_q[3617] : 
                                (N190)? btb_q[3682] : 
                                (N192)? btb_q[3747] : 
                                (N194)? btb_q[3812] : 
                                (N196)? btb_q[3877] : 
                                (N198)? btb_q[3942] : 
                                (N200)? btb_q[4007] : 
                                (N202)? btb_q[4072] : 
                                (N204)? btb_q[4137] : 1'b0;
  assign btb_prediction_o[41] = (N141)? btb_q[41] : 
                                (N143)? btb_q[106] : 
                                (N145)? btb_q[171] : 
                                (N147)? btb_q[236] : 
                                (N149)? btb_q[301] : 
                                (N151)? btb_q[366] : 
                                (N153)? btb_q[431] : 
                                (N155)? btb_q[496] : 
                                (N157)? btb_q[561] : 
                                (N159)? btb_q[626] : 
                                (N161)? btb_q[691] : 
                                (N163)? btb_q[756] : 
                                (N165)? btb_q[821] : 
                                (N167)? btb_q[886] : 
                                (N169)? btb_q[951] : 
                                (N171)? btb_q[1016] : 
                                (N173)? btb_q[1081] : 
                                (N175)? btb_q[1146] : 
                                (N177)? btb_q[1211] : 
                                (N179)? btb_q[1276] : 
                                (N181)? btb_q[1341] : 
                                (N183)? btb_q[1406] : 
                                (N185)? btb_q[1471] : 
                                (N187)? btb_q[1536] : 
                                (N189)? btb_q[1601] : 
                                (N191)? btb_q[1666] : 
                                (N193)? btb_q[1731] : 
                                (N195)? btb_q[1796] : 
                                (N197)? btb_q[1861] : 
                                (N199)? btb_q[1926] : 
                                (N201)? btb_q[1991] : 
                                (N203)? btb_q[2056] : 
                                (N142)? btb_q[2121] : 
                                (N144)? btb_q[2186] : 
                                (N146)? btb_q[2251] : 
                                (N148)? btb_q[2316] : 
                                (N150)? btb_q[2381] : 
                                (N152)? btb_q[2446] : 
                                (N154)? btb_q[2511] : 
                                (N156)? btb_q[2576] : 
                                (N158)? btb_q[2641] : 
                                (N160)? btb_q[2706] : 
                                (N162)? btb_q[2771] : 
                                (N164)? btb_q[2836] : 
                                (N166)? btb_q[2901] : 
                                (N168)? btb_q[2966] : 
                                (N170)? btb_q[3031] : 
                                (N172)? btb_q[3096] : 
                                (N174)? btb_q[3161] : 
                                (N176)? btb_q[3226] : 
                                (N178)? btb_q[3291] : 
                                (N180)? btb_q[3356] : 
                                (N182)? btb_q[3421] : 
                                (N184)? btb_q[3486] : 
                                (N186)? btb_q[3551] : 
                                (N188)? btb_q[3616] : 
                                (N190)? btb_q[3681] : 
                                (N192)? btb_q[3746] : 
                                (N194)? btb_q[3811] : 
                                (N196)? btb_q[3876] : 
                                (N198)? btb_q[3941] : 
                                (N200)? btb_q[4006] : 
                                (N202)? btb_q[4071] : 
                                (N204)? btb_q[4136] : 1'b0;
  assign btb_prediction_o[40] = (N141)? btb_q[40] : 
                                (N143)? btb_q[105] : 
                                (N145)? btb_q[170] : 
                                (N147)? btb_q[235] : 
                                (N149)? btb_q[300] : 
                                (N151)? btb_q[365] : 
                                (N153)? btb_q[430] : 
                                (N155)? btb_q[495] : 
                                (N157)? btb_q[560] : 
                                (N159)? btb_q[625] : 
                                (N161)? btb_q[690] : 
                                (N163)? btb_q[755] : 
                                (N165)? btb_q[820] : 
                                (N167)? btb_q[885] : 
                                (N169)? btb_q[950] : 
                                (N171)? btb_q[1015] : 
                                (N173)? btb_q[1080] : 
                                (N175)? btb_q[1145] : 
                                (N177)? btb_q[1210] : 
                                (N179)? btb_q[1275] : 
                                (N181)? btb_q[1340] : 
                                (N183)? btb_q[1405] : 
                                (N185)? btb_q[1470] : 
                                (N187)? btb_q[1535] : 
                                (N189)? btb_q[1600] : 
                                (N191)? btb_q[1665] : 
                                (N193)? btb_q[1730] : 
                                (N195)? btb_q[1795] : 
                                (N197)? btb_q[1860] : 
                                (N199)? btb_q[1925] : 
                                (N201)? btb_q[1990] : 
                                (N203)? btb_q[2055] : 
                                (N142)? btb_q[2120] : 
                                (N144)? btb_q[2185] : 
                                (N146)? btb_q[2250] : 
                                (N148)? btb_q[2315] : 
                                (N150)? btb_q[2380] : 
                                (N152)? btb_q[2445] : 
                                (N154)? btb_q[2510] : 
                                (N156)? btb_q[2575] : 
                                (N158)? btb_q[2640] : 
                                (N160)? btb_q[2705] : 
                                (N162)? btb_q[2770] : 
                                (N164)? btb_q[2835] : 
                                (N166)? btb_q[2900] : 
                                (N168)? btb_q[2965] : 
                                (N170)? btb_q[3030] : 
                                (N172)? btb_q[3095] : 
                                (N174)? btb_q[3160] : 
                                (N176)? btb_q[3225] : 
                                (N178)? btb_q[3290] : 
                                (N180)? btb_q[3355] : 
                                (N182)? btb_q[3420] : 
                                (N184)? btb_q[3485] : 
                                (N186)? btb_q[3550] : 
                                (N188)? btb_q[3615] : 
                                (N190)? btb_q[3680] : 
                                (N192)? btb_q[3745] : 
                                (N194)? btb_q[3810] : 
                                (N196)? btb_q[3875] : 
                                (N198)? btb_q[3940] : 
                                (N200)? btb_q[4005] : 
                                (N202)? btb_q[4070] : 
                                (N204)? btb_q[4135] : 1'b0;
  assign btb_prediction_o[39] = (N141)? btb_q[39] : 
                                (N143)? btb_q[104] : 
                                (N145)? btb_q[169] : 
                                (N147)? btb_q[234] : 
                                (N149)? btb_q[299] : 
                                (N151)? btb_q[364] : 
                                (N153)? btb_q[429] : 
                                (N155)? btb_q[494] : 
                                (N157)? btb_q[559] : 
                                (N159)? btb_q[624] : 
                                (N161)? btb_q[689] : 
                                (N163)? btb_q[754] : 
                                (N165)? btb_q[819] : 
                                (N167)? btb_q[884] : 
                                (N169)? btb_q[949] : 
                                (N171)? btb_q[1014] : 
                                (N173)? btb_q[1079] : 
                                (N175)? btb_q[1144] : 
                                (N177)? btb_q[1209] : 
                                (N179)? btb_q[1274] : 
                                (N181)? btb_q[1339] : 
                                (N183)? btb_q[1404] : 
                                (N185)? btb_q[1469] : 
                                (N187)? btb_q[1534] : 
                                (N189)? btb_q[1599] : 
                                (N191)? btb_q[1664] : 
                                (N193)? btb_q[1729] : 
                                (N195)? btb_q[1794] : 
                                (N197)? btb_q[1859] : 
                                (N199)? btb_q[1924] : 
                                (N201)? btb_q[1989] : 
                                (N203)? btb_q[2054] : 
                                (N142)? btb_q[2119] : 
                                (N144)? btb_q[2184] : 
                                (N146)? btb_q[2249] : 
                                (N148)? btb_q[2314] : 
                                (N150)? btb_q[2379] : 
                                (N152)? btb_q[2444] : 
                                (N154)? btb_q[2509] : 
                                (N156)? btb_q[2574] : 
                                (N158)? btb_q[2639] : 
                                (N160)? btb_q[2704] : 
                                (N162)? btb_q[2769] : 
                                (N164)? btb_q[2834] : 
                                (N166)? btb_q[2899] : 
                                (N168)? btb_q[2964] : 
                                (N170)? btb_q[3029] : 
                                (N172)? btb_q[3094] : 
                                (N174)? btb_q[3159] : 
                                (N176)? btb_q[3224] : 
                                (N178)? btb_q[3289] : 
                                (N180)? btb_q[3354] : 
                                (N182)? btb_q[3419] : 
                                (N184)? btb_q[3484] : 
                                (N186)? btb_q[3549] : 
                                (N188)? btb_q[3614] : 
                                (N190)? btb_q[3679] : 
                                (N192)? btb_q[3744] : 
                                (N194)? btb_q[3809] : 
                                (N196)? btb_q[3874] : 
                                (N198)? btb_q[3939] : 
                                (N200)? btb_q[4004] : 
                                (N202)? btb_q[4069] : 
                                (N204)? btb_q[4134] : 1'b0;
  assign btb_prediction_o[38] = (N141)? btb_q[38] : 
                                (N143)? btb_q[103] : 
                                (N145)? btb_q[168] : 
                                (N147)? btb_q[233] : 
                                (N149)? btb_q[298] : 
                                (N151)? btb_q[363] : 
                                (N153)? btb_q[428] : 
                                (N155)? btb_q[493] : 
                                (N157)? btb_q[558] : 
                                (N159)? btb_q[623] : 
                                (N161)? btb_q[688] : 
                                (N163)? btb_q[753] : 
                                (N165)? btb_q[818] : 
                                (N167)? btb_q[883] : 
                                (N169)? btb_q[948] : 
                                (N171)? btb_q[1013] : 
                                (N173)? btb_q[1078] : 
                                (N175)? btb_q[1143] : 
                                (N177)? btb_q[1208] : 
                                (N179)? btb_q[1273] : 
                                (N181)? btb_q[1338] : 
                                (N183)? btb_q[1403] : 
                                (N185)? btb_q[1468] : 
                                (N187)? btb_q[1533] : 
                                (N189)? btb_q[1598] : 
                                (N191)? btb_q[1663] : 
                                (N193)? btb_q[1728] : 
                                (N195)? btb_q[1793] : 
                                (N197)? btb_q[1858] : 
                                (N199)? btb_q[1923] : 
                                (N201)? btb_q[1988] : 
                                (N203)? btb_q[2053] : 
                                (N142)? btb_q[2118] : 
                                (N144)? btb_q[2183] : 
                                (N146)? btb_q[2248] : 
                                (N148)? btb_q[2313] : 
                                (N150)? btb_q[2378] : 
                                (N152)? btb_q[2443] : 
                                (N154)? btb_q[2508] : 
                                (N156)? btb_q[2573] : 
                                (N158)? btb_q[2638] : 
                                (N160)? btb_q[2703] : 
                                (N162)? btb_q[2768] : 
                                (N164)? btb_q[2833] : 
                                (N166)? btb_q[2898] : 
                                (N168)? btb_q[2963] : 
                                (N170)? btb_q[3028] : 
                                (N172)? btb_q[3093] : 
                                (N174)? btb_q[3158] : 
                                (N176)? btb_q[3223] : 
                                (N178)? btb_q[3288] : 
                                (N180)? btb_q[3353] : 
                                (N182)? btb_q[3418] : 
                                (N184)? btb_q[3483] : 
                                (N186)? btb_q[3548] : 
                                (N188)? btb_q[3613] : 
                                (N190)? btb_q[3678] : 
                                (N192)? btb_q[3743] : 
                                (N194)? btb_q[3808] : 
                                (N196)? btb_q[3873] : 
                                (N198)? btb_q[3938] : 
                                (N200)? btb_q[4003] : 
                                (N202)? btb_q[4068] : 
                                (N204)? btb_q[4133] : 1'b0;
  assign btb_prediction_o[37] = (N141)? btb_q[37] : 
                                (N143)? btb_q[102] : 
                                (N145)? btb_q[167] : 
                                (N147)? btb_q[232] : 
                                (N149)? btb_q[297] : 
                                (N151)? btb_q[362] : 
                                (N153)? btb_q[427] : 
                                (N155)? btb_q[492] : 
                                (N157)? btb_q[557] : 
                                (N159)? btb_q[622] : 
                                (N161)? btb_q[687] : 
                                (N163)? btb_q[752] : 
                                (N165)? btb_q[817] : 
                                (N167)? btb_q[882] : 
                                (N169)? btb_q[947] : 
                                (N171)? btb_q[1012] : 
                                (N173)? btb_q[1077] : 
                                (N175)? btb_q[1142] : 
                                (N177)? btb_q[1207] : 
                                (N179)? btb_q[1272] : 
                                (N181)? btb_q[1337] : 
                                (N183)? btb_q[1402] : 
                                (N185)? btb_q[1467] : 
                                (N187)? btb_q[1532] : 
                                (N189)? btb_q[1597] : 
                                (N191)? btb_q[1662] : 
                                (N193)? btb_q[1727] : 
                                (N195)? btb_q[1792] : 
                                (N197)? btb_q[1857] : 
                                (N199)? btb_q[1922] : 
                                (N201)? btb_q[1987] : 
                                (N203)? btb_q[2052] : 
                                (N142)? btb_q[2117] : 
                                (N144)? btb_q[2182] : 
                                (N146)? btb_q[2247] : 
                                (N148)? btb_q[2312] : 
                                (N150)? btb_q[2377] : 
                                (N152)? btb_q[2442] : 
                                (N154)? btb_q[2507] : 
                                (N156)? btb_q[2572] : 
                                (N158)? btb_q[2637] : 
                                (N160)? btb_q[2702] : 
                                (N162)? btb_q[2767] : 
                                (N164)? btb_q[2832] : 
                                (N166)? btb_q[2897] : 
                                (N168)? btb_q[2962] : 
                                (N170)? btb_q[3027] : 
                                (N172)? btb_q[3092] : 
                                (N174)? btb_q[3157] : 
                                (N176)? btb_q[3222] : 
                                (N178)? btb_q[3287] : 
                                (N180)? btb_q[3352] : 
                                (N182)? btb_q[3417] : 
                                (N184)? btb_q[3482] : 
                                (N186)? btb_q[3547] : 
                                (N188)? btb_q[3612] : 
                                (N190)? btb_q[3677] : 
                                (N192)? btb_q[3742] : 
                                (N194)? btb_q[3807] : 
                                (N196)? btb_q[3872] : 
                                (N198)? btb_q[3937] : 
                                (N200)? btb_q[4002] : 
                                (N202)? btb_q[4067] : 
                                (N204)? btb_q[4132] : 1'b0;
  assign btb_prediction_o[36] = (N141)? btb_q[36] : 
                                (N143)? btb_q[101] : 
                                (N145)? btb_q[166] : 
                                (N147)? btb_q[231] : 
                                (N149)? btb_q[296] : 
                                (N151)? btb_q[361] : 
                                (N153)? btb_q[426] : 
                                (N155)? btb_q[491] : 
                                (N157)? btb_q[556] : 
                                (N159)? btb_q[621] : 
                                (N161)? btb_q[686] : 
                                (N163)? btb_q[751] : 
                                (N165)? btb_q[816] : 
                                (N167)? btb_q[881] : 
                                (N169)? btb_q[946] : 
                                (N171)? btb_q[1011] : 
                                (N173)? btb_q[1076] : 
                                (N175)? btb_q[1141] : 
                                (N177)? btb_q[1206] : 
                                (N179)? btb_q[1271] : 
                                (N181)? btb_q[1336] : 
                                (N183)? btb_q[1401] : 
                                (N185)? btb_q[1466] : 
                                (N187)? btb_q[1531] : 
                                (N189)? btb_q[1596] : 
                                (N191)? btb_q[1661] : 
                                (N193)? btb_q[1726] : 
                                (N195)? btb_q[1791] : 
                                (N197)? btb_q[1856] : 
                                (N199)? btb_q[1921] : 
                                (N201)? btb_q[1986] : 
                                (N203)? btb_q[2051] : 
                                (N142)? btb_q[2116] : 
                                (N144)? btb_q[2181] : 
                                (N146)? btb_q[2246] : 
                                (N148)? btb_q[2311] : 
                                (N150)? btb_q[2376] : 
                                (N152)? btb_q[2441] : 
                                (N154)? btb_q[2506] : 
                                (N156)? btb_q[2571] : 
                                (N158)? btb_q[2636] : 
                                (N160)? btb_q[2701] : 
                                (N162)? btb_q[2766] : 
                                (N164)? btb_q[2831] : 
                                (N166)? btb_q[2896] : 
                                (N168)? btb_q[2961] : 
                                (N170)? btb_q[3026] : 
                                (N172)? btb_q[3091] : 
                                (N174)? btb_q[3156] : 
                                (N176)? btb_q[3221] : 
                                (N178)? btb_q[3286] : 
                                (N180)? btb_q[3351] : 
                                (N182)? btb_q[3416] : 
                                (N184)? btb_q[3481] : 
                                (N186)? btb_q[3546] : 
                                (N188)? btb_q[3611] : 
                                (N190)? btb_q[3676] : 
                                (N192)? btb_q[3741] : 
                                (N194)? btb_q[3806] : 
                                (N196)? btb_q[3871] : 
                                (N198)? btb_q[3936] : 
                                (N200)? btb_q[4001] : 
                                (N202)? btb_q[4066] : 
                                (N204)? btb_q[4131] : 1'b0;
  assign btb_prediction_o[35] = (N141)? btb_q[35] : 
                                (N143)? btb_q[100] : 
                                (N145)? btb_q[165] : 
                                (N147)? btb_q[230] : 
                                (N149)? btb_q[295] : 
                                (N151)? btb_q[360] : 
                                (N153)? btb_q[425] : 
                                (N155)? btb_q[490] : 
                                (N157)? btb_q[555] : 
                                (N159)? btb_q[620] : 
                                (N161)? btb_q[685] : 
                                (N163)? btb_q[750] : 
                                (N165)? btb_q[815] : 
                                (N167)? btb_q[880] : 
                                (N169)? btb_q[945] : 
                                (N171)? btb_q[1010] : 
                                (N173)? btb_q[1075] : 
                                (N175)? btb_q[1140] : 
                                (N177)? btb_q[1205] : 
                                (N179)? btb_q[1270] : 
                                (N181)? btb_q[1335] : 
                                (N183)? btb_q[1400] : 
                                (N185)? btb_q[1465] : 
                                (N187)? btb_q[1530] : 
                                (N189)? btb_q[1595] : 
                                (N191)? btb_q[1660] : 
                                (N193)? btb_q[1725] : 
                                (N195)? btb_q[1790] : 
                                (N197)? btb_q[1855] : 
                                (N199)? btb_q[1920] : 
                                (N201)? btb_q[1985] : 
                                (N203)? btb_q[2050] : 
                                (N142)? btb_q[2115] : 
                                (N144)? btb_q[2180] : 
                                (N146)? btb_q[2245] : 
                                (N148)? btb_q[2310] : 
                                (N150)? btb_q[2375] : 
                                (N152)? btb_q[2440] : 
                                (N154)? btb_q[2505] : 
                                (N156)? btb_q[2570] : 
                                (N158)? btb_q[2635] : 
                                (N160)? btb_q[2700] : 
                                (N162)? btb_q[2765] : 
                                (N164)? btb_q[2830] : 
                                (N166)? btb_q[2895] : 
                                (N168)? btb_q[2960] : 
                                (N170)? btb_q[3025] : 
                                (N172)? btb_q[3090] : 
                                (N174)? btb_q[3155] : 
                                (N176)? btb_q[3220] : 
                                (N178)? btb_q[3285] : 
                                (N180)? btb_q[3350] : 
                                (N182)? btb_q[3415] : 
                                (N184)? btb_q[3480] : 
                                (N186)? btb_q[3545] : 
                                (N188)? btb_q[3610] : 
                                (N190)? btb_q[3675] : 
                                (N192)? btb_q[3740] : 
                                (N194)? btb_q[3805] : 
                                (N196)? btb_q[3870] : 
                                (N198)? btb_q[3935] : 
                                (N200)? btb_q[4000] : 
                                (N202)? btb_q[4065] : 
                                (N204)? btb_q[4130] : 1'b0;
  assign btb_prediction_o[34] = (N141)? btb_q[34] : 
                                (N143)? btb_q[99] : 
                                (N145)? btb_q[164] : 
                                (N147)? btb_q[229] : 
                                (N149)? btb_q[294] : 
                                (N151)? btb_q[359] : 
                                (N153)? btb_q[424] : 
                                (N155)? btb_q[489] : 
                                (N157)? btb_q[554] : 
                                (N159)? btb_q[619] : 
                                (N161)? btb_q[684] : 
                                (N163)? btb_q[749] : 
                                (N165)? btb_q[814] : 
                                (N167)? btb_q[879] : 
                                (N169)? btb_q[944] : 
                                (N171)? btb_q[1009] : 
                                (N173)? btb_q[1074] : 
                                (N175)? btb_q[1139] : 
                                (N177)? btb_q[1204] : 
                                (N179)? btb_q[1269] : 
                                (N181)? btb_q[1334] : 
                                (N183)? btb_q[1399] : 
                                (N185)? btb_q[1464] : 
                                (N187)? btb_q[1529] : 
                                (N189)? btb_q[1594] : 
                                (N191)? btb_q[1659] : 
                                (N193)? btb_q[1724] : 
                                (N195)? btb_q[1789] : 
                                (N197)? btb_q[1854] : 
                                (N199)? btb_q[1919] : 
                                (N201)? btb_q[1984] : 
                                (N203)? btb_q[2049] : 
                                (N142)? btb_q[2114] : 
                                (N144)? btb_q[2179] : 
                                (N146)? btb_q[2244] : 
                                (N148)? btb_q[2309] : 
                                (N150)? btb_q[2374] : 
                                (N152)? btb_q[2439] : 
                                (N154)? btb_q[2504] : 
                                (N156)? btb_q[2569] : 
                                (N158)? btb_q[2634] : 
                                (N160)? btb_q[2699] : 
                                (N162)? btb_q[2764] : 
                                (N164)? btb_q[2829] : 
                                (N166)? btb_q[2894] : 
                                (N168)? btb_q[2959] : 
                                (N170)? btb_q[3024] : 
                                (N172)? btb_q[3089] : 
                                (N174)? btb_q[3154] : 
                                (N176)? btb_q[3219] : 
                                (N178)? btb_q[3284] : 
                                (N180)? btb_q[3349] : 
                                (N182)? btb_q[3414] : 
                                (N184)? btb_q[3479] : 
                                (N186)? btb_q[3544] : 
                                (N188)? btb_q[3609] : 
                                (N190)? btb_q[3674] : 
                                (N192)? btb_q[3739] : 
                                (N194)? btb_q[3804] : 
                                (N196)? btb_q[3869] : 
                                (N198)? btb_q[3934] : 
                                (N200)? btb_q[3999] : 
                                (N202)? btb_q[4064] : 
                                (N204)? btb_q[4129] : 1'b0;
  assign btb_prediction_o[33] = (N141)? btb_q[33] : 
                                (N143)? btb_q[98] : 
                                (N145)? btb_q[163] : 
                                (N147)? btb_q[228] : 
                                (N149)? btb_q[293] : 
                                (N151)? btb_q[358] : 
                                (N153)? btb_q[423] : 
                                (N155)? btb_q[488] : 
                                (N157)? btb_q[553] : 
                                (N159)? btb_q[618] : 
                                (N161)? btb_q[683] : 
                                (N163)? btb_q[748] : 
                                (N165)? btb_q[813] : 
                                (N167)? btb_q[878] : 
                                (N169)? btb_q[943] : 
                                (N171)? btb_q[1008] : 
                                (N173)? btb_q[1073] : 
                                (N175)? btb_q[1138] : 
                                (N177)? btb_q[1203] : 
                                (N179)? btb_q[1268] : 
                                (N181)? btb_q[1333] : 
                                (N183)? btb_q[1398] : 
                                (N185)? btb_q[1463] : 
                                (N187)? btb_q[1528] : 
                                (N189)? btb_q[1593] : 
                                (N191)? btb_q[1658] : 
                                (N193)? btb_q[1723] : 
                                (N195)? btb_q[1788] : 
                                (N197)? btb_q[1853] : 
                                (N199)? btb_q[1918] : 
                                (N201)? btb_q[1983] : 
                                (N203)? btb_q[2048] : 
                                (N142)? btb_q[2113] : 
                                (N144)? btb_q[2178] : 
                                (N146)? btb_q[2243] : 
                                (N148)? btb_q[2308] : 
                                (N150)? btb_q[2373] : 
                                (N152)? btb_q[2438] : 
                                (N154)? btb_q[2503] : 
                                (N156)? btb_q[2568] : 
                                (N158)? btb_q[2633] : 
                                (N160)? btb_q[2698] : 
                                (N162)? btb_q[2763] : 
                                (N164)? btb_q[2828] : 
                                (N166)? btb_q[2893] : 
                                (N168)? btb_q[2958] : 
                                (N170)? btb_q[3023] : 
                                (N172)? btb_q[3088] : 
                                (N174)? btb_q[3153] : 
                                (N176)? btb_q[3218] : 
                                (N178)? btb_q[3283] : 
                                (N180)? btb_q[3348] : 
                                (N182)? btb_q[3413] : 
                                (N184)? btb_q[3478] : 
                                (N186)? btb_q[3543] : 
                                (N188)? btb_q[3608] : 
                                (N190)? btb_q[3673] : 
                                (N192)? btb_q[3738] : 
                                (N194)? btb_q[3803] : 
                                (N196)? btb_q[3868] : 
                                (N198)? btb_q[3933] : 
                                (N200)? btb_q[3998] : 
                                (N202)? btb_q[4063] : 
                                (N204)? btb_q[4128] : 1'b0;
  assign btb_prediction_o[32] = (N141)? btb_q[32] : 
                                (N143)? btb_q[97] : 
                                (N145)? btb_q[162] : 
                                (N147)? btb_q[227] : 
                                (N149)? btb_q[292] : 
                                (N151)? btb_q[357] : 
                                (N153)? btb_q[422] : 
                                (N155)? btb_q[487] : 
                                (N157)? btb_q[552] : 
                                (N159)? btb_q[617] : 
                                (N161)? btb_q[682] : 
                                (N163)? btb_q[747] : 
                                (N165)? btb_q[812] : 
                                (N167)? btb_q[877] : 
                                (N169)? btb_q[942] : 
                                (N171)? btb_q[1007] : 
                                (N173)? btb_q[1072] : 
                                (N175)? btb_q[1137] : 
                                (N177)? btb_q[1202] : 
                                (N179)? btb_q[1267] : 
                                (N181)? btb_q[1332] : 
                                (N183)? btb_q[1397] : 
                                (N185)? btb_q[1462] : 
                                (N187)? btb_q[1527] : 
                                (N189)? btb_q[1592] : 
                                (N191)? btb_q[1657] : 
                                (N193)? btb_q[1722] : 
                                (N195)? btb_q[1787] : 
                                (N197)? btb_q[1852] : 
                                (N199)? btb_q[1917] : 
                                (N201)? btb_q[1982] : 
                                (N203)? btb_q[2047] : 
                                (N142)? btb_q[2112] : 
                                (N144)? btb_q[2177] : 
                                (N146)? btb_q[2242] : 
                                (N148)? btb_q[2307] : 
                                (N150)? btb_q[2372] : 
                                (N152)? btb_q[2437] : 
                                (N154)? btb_q[2502] : 
                                (N156)? btb_q[2567] : 
                                (N158)? btb_q[2632] : 
                                (N160)? btb_q[2697] : 
                                (N162)? btb_q[2762] : 
                                (N164)? btb_q[2827] : 
                                (N166)? btb_q[2892] : 
                                (N168)? btb_q[2957] : 
                                (N170)? btb_q[3022] : 
                                (N172)? btb_q[3087] : 
                                (N174)? btb_q[3152] : 
                                (N176)? btb_q[3217] : 
                                (N178)? btb_q[3282] : 
                                (N180)? btb_q[3347] : 
                                (N182)? btb_q[3412] : 
                                (N184)? btb_q[3477] : 
                                (N186)? btb_q[3542] : 
                                (N188)? btb_q[3607] : 
                                (N190)? btb_q[3672] : 
                                (N192)? btb_q[3737] : 
                                (N194)? btb_q[3802] : 
                                (N196)? btb_q[3867] : 
                                (N198)? btb_q[3932] : 
                                (N200)? btb_q[3997] : 
                                (N202)? btb_q[4062] : 
                                (N204)? btb_q[4127] : 1'b0;
  assign btb_prediction_o[31] = (N141)? btb_q[31] : 
                                (N143)? btb_q[96] : 
                                (N145)? btb_q[161] : 
                                (N147)? btb_q[226] : 
                                (N149)? btb_q[291] : 
                                (N151)? btb_q[356] : 
                                (N153)? btb_q[421] : 
                                (N155)? btb_q[486] : 
                                (N157)? btb_q[551] : 
                                (N159)? btb_q[616] : 
                                (N161)? btb_q[681] : 
                                (N163)? btb_q[746] : 
                                (N165)? btb_q[811] : 
                                (N167)? btb_q[876] : 
                                (N169)? btb_q[941] : 
                                (N171)? btb_q[1006] : 
                                (N173)? btb_q[1071] : 
                                (N175)? btb_q[1136] : 
                                (N177)? btb_q[1201] : 
                                (N179)? btb_q[1266] : 
                                (N181)? btb_q[1331] : 
                                (N183)? btb_q[1396] : 
                                (N185)? btb_q[1461] : 
                                (N187)? btb_q[1526] : 
                                (N189)? btb_q[1591] : 
                                (N191)? btb_q[1656] : 
                                (N193)? btb_q[1721] : 
                                (N195)? btb_q[1786] : 
                                (N197)? btb_q[1851] : 
                                (N199)? btb_q[1916] : 
                                (N201)? btb_q[1981] : 
                                (N203)? btb_q[2046] : 
                                (N142)? btb_q[2111] : 
                                (N144)? btb_q[2176] : 
                                (N146)? btb_q[2241] : 
                                (N148)? btb_q[2306] : 
                                (N150)? btb_q[2371] : 
                                (N152)? btb_q[2436] : 
                                (N154)? btb_q[2501] : 
                                (N156)? btb_q[2566] : 
                                (N158)? btb_q[2631] : 
                                (N160)? btb_q[2696] : 
                                (N162)? btb_q[2761] : 
                                (N164)? btb_q[2826] : 
                                (N166)? btb_q[2891] : 
                                (N168)? btb_q[2956] : 
                                (N170)? btb_q[3021] : 
                                (N172)? btb_q[3086] : 
                                (N174)? btb_q[3151] : 
                                (N176)? btb_q[3216] : 
                                (N178)? btb_q[3281] : 
                                (N180)? btb_q[3346] : 
                                (N182)? btb_q[3411] : 
                                (N184)? btb_q[3476] : 
                                (N186)? btb_q[3541] : 
                                (N188)? btb_q[3606] : 
                                (N190)? btb_q[3671] : 
                                (N192)? btb_q[3736] : 
                                (N194)? btb_q[3801] : 
                                (N196)? btb_q[3866] : 
                                (N198)? btb_q[3931] : 
                                (N200)? btb_q[3996] : 
                                (N202)? btb_q[4061] : 
                                (N204)? btb_q[4126] : 1'b0;
  assign btb_prediction_o[30] = (N141)? btb_q[30] : 
                                (N143)? btb_q[95] : 
                                (N145)? btb_q[160] : 
                                (N147)? btb_q[225] : 
                                (N149)? btb_q[290] : 
                                (N151)? btb_q[355] : 
                                (N153)? btb_q[420] : 
                                (N155)? btb_q[485] : 
                                (N157)? btb_q[550] : 
                                (N159)? btb_q[615] : 
                                (N161)? btb_q[680] : 
                                (N163)? btb_q[745] : 
                                (N165)? btb_q[810] : 
                                (N167)? btb_q[875] : 
                                (N169)? btb_q[940] : 
                                (N171)? btb_q[1005] : 
                                (N173)? btb_q[1070] : 
                                (N175)? btb_q[1135] : 
                                (N177)? btb_q[1200] : 
                                (N179)? btb_q[1265] : 
                                (N181)? btb_q[1330] : 
                                (N183)? btb_q[1395] : 
                                (N185)? btb_q[1460] : 
                                (N187)? btb_q[1525] : 
                                (N189)? btb_q[1590] : 
                                (N191)? btb_q[1655] : 
                                (N193)? btb_q[1720] : 
                                (N195)? btb_q[1785] : 
                                (N197)? btb_q[1850] : 
                                (N199)? btb_q[1915] : 
                                (N201)? btb_q[1980] : 
                                (N203)? btb_q[2045] : 
                                (N142)? btb_q[2110] : 
                                (N144)? btb_q[2175] : 
                                (N146)? btb_q[2240] : 
                                (N148)? btb_q[2305] : 
                                (N150)? btb_q[2370] : 
                                (N152)? btb_q[2435] : 
                                (N154)? btb_q[2500] : 
                                (N156)? btb_q[2565] : 
                                (N158)? btb_q[2630] : 
                                (N160)? btb_q[2695] : 
                                (N162)? btb_q[2760] : 
                                (N164)? btb_q[2825] : 
                                (N166)? btb_q[2890] : 
                                (N168)? btb_q[2955] : 
                                (N170)? btb_q[3020] : 
                                (N172)? btb_q[3085] : 
                                (N174)? btb_q[3150] : 
                                (N176)? btb_q[3215] : 
                                (N178)? btb_q[3280] : 
                                (N180)? btb_q[3345] : 
                                (N182)? btb_q[3410] : 
                                (N184)? btb_q[3475] : 
                                (N186)? btb_q[3540] : 
                                (N188)? btb_q[3605] : 
                                (N190)? btb_q[3670] : 
                                (N192)? btb_q[3735] : 
                                (N194)? btb_q[3800] : 
                                (N196)? btb_q[3865] : 
                                (N198)? btb_q[3930] : 
                                (N200)? btb_q[3995] : 
                                (N202)? btb_q[4060] : 
                                (N204)? btb_q[4125] : 1'b0;
  assign btb_prediction_o[29] = (N141)? btb_q[29] : 
                                (N143)? btb_q[94] : 
                                (N145)? btb_q[159] : 
                                (N147)? btb_q[224] : 
                                (N149)? btb_q[289] : 
                                (N151)? btb_q[354] : 
                                (N153)? btb_q[419] : 
                                (N155)? btb_q[484] : 
                                (N157)? btb_q[549] : 
                                (N159)? btb_q[614] : 
                                (N161)? btb_q[679] : 
                                (N163)? btb_q[744] : 
                                (N165)? btb_q[809] : 
                                (N167)? btb_q[874] : 
                                (N169)? btb_q[939] : 
                                (N171)? btb_q[1004] : 
                                (N173)? btb_q[1069] : 
                                (N175)? btb_q[1134] : 
                                (N177)? btb_q[1199] : 
                                (N179)? btb_q[1264] : 
                                (N181)? btb_q[1329] : 
                                (N183)? btb_q[1394] : 
                                (N185)? btb_q[1459] : 
                                (N187)? btb_q[1524] : 
                                (N189)? btb_q[1589] : 
                                (N191)? btb_q[1654] : 
                                (N193)? btb_q[1719] : 
                                (N195)? btb_q[1784] : 
                                (N197)? btb_q[1849] : 
                                (N199)? btb_q[1914] : 
                                (N201)? btb_q[1979] : 
                                (N203)? btb_q[2044] : 
                                (N142)? btb_q[2109] : 
                                (N144)? btb_q[2174] : 
                                (N146)? btb_q[2239] : 
                                (N148)? btb_q[2304] : 
                                (N150)? btb_q[2369] : 
                                (N152)? btb_q[2434] : 
                                (N154)? btb_q[2499] : 
                                (N156)? btb_q[2564] : 
                                (N158)? btb_q[2629] : 
                                (N160)? btb_q[2694] : 
                                (N162)? btb_q[2759] : 
                                (N164)? btb_q[2824] : 
                                (N166)? btb_q[2889] : 
                                (N168)? btb_q[2954] : 
                                (N170)? btb_q[3019] : 
                                (N172)? btb_q[3084] : 
                                (N174)? btb_q[3149] : 
                                (N176)? btb_q[3214] : 
                                (N178)? btb_q[3279] : 
                                (N180)? btb_q[3344] : 
                                (N182)? btb_q[3409] : 
                                (N184)? btb_q[3474] : 
                                (N186)? btb_q[3539] : 
                                (N188)? btb_q[3604] : 
                                (N190)? btb_q[3669] : 
                                (N192)? btb_q[3734] : 
                                (N194)? btb_q[3799] : 
                                (N196)? btb_q[3864] : 
                                (N198)? btb_q[3929] : 
                                (N200)? btb_q[3994] : 
                                (N202)? btb_q[4059] : 
                                (N204)? btb_q[4124] : 1'b0;
  assign btb_prediction_o[28] = (N141)? btb_q[28] : 
                                (N143)? btb_q[93] : 
                                (N145)? btb_q[158] : 
                                (N147)? btb_q[223] : 
                                (N149)? btb_q[288] : 
                                (N151)? btb_q[353] : 
                                (N153)? btb_q[418] : 
                                (N155)? btb_q[483] : 
                                (N157)? btb_q[548] : 
                                (N159)? btb_q[613] : 
                                (N161)? btb_q[678] : 
                                (N163)? btb_q[743] : 
                                (N165)? btb_q[808] : 
                                (N167)? btb_q[873] : 
                                (N169)? btb_q[938] : 
                                (N171)? btb_q[1003] : 
                                (N173)? btb_q[1068] : 
                                (N175)? btb_q[1133] : 
                                (N177)? btb_q[1198] : 
                                (N179)? btb_q[1263] : 
                                (N181)? btb_q[1328] : 
                                (N183)? btb_q[1393] : 
                                (N185)? btb_q[1458] : 
                                (N187)? btb_q[1523] : 
                                (N189)? btb_q[1588] : 
                                (N191)? btb_q[1653] : 
                                (N193)? btb_q[1718] : 
                                (N195)? btb_q[1783] : 
                                (N197)? btb_q[1848] : 
                                (N199)? btb_q[1913] : 
                                (N201)? btb_q[1978] : 
                                (N203)? btb_q[2043] : 
                                (N142)? btb_q[2108] : 
                                (N144)? btb_q[2173] : 
                                (N146)? btb_q[2238] : 
                                (N148)? btb_q[2303] : 
                                (N150)? btb_q[2368] : 
                                (N152)? btb_q[2433] : 
                                (N154)? btb_q[2498] : 
                                (N156)? btb_q[2563] : 
                                (N158)? btb_q[2628] : 
                                (N160)? btb_q[2693] : 
                                (N162)? btb_q[2758] : 
                                (N164)? btb_q[2823] : 
                                (N166)? btb_q[2888] : 
                                (N168)? btb_q[2953] : 
                                (N170)? btb_q[3018] : 
                                (N172)? btb_q[3083] : 
                                (N174)? btb_q[3148] : 
                                (N176)? btb_q[3213] : 
                                (N178)? btb_q[3278] : 
                                (N180)? btb_q[3343] : 
                                (N182)? btb_q[3408] : 
                                (N184)? btb_q[3473] : 
                                (N186)? btb_q[3538] : 
                                (N188)? btb_q[3603] : 
                                (N190)? btb_q[3668] : 
                                (N192)? btb_q[3733] : 
                                (N194)? btb_q[3798] : 
                                (N196)? btb_q[3863] : 
                                (N198)? btb_q[3928] : 
                                (N200)? btb_q[3993] : 
                                (N202)? btb_q[4058] : 
                                (N204)? btb_q[4123] : 1'b0;
  assign btb_prediction_o[27] = (N141)? btb_q[27] : 
                                (N143)? btb_q[92] : 
                                (N145)? btb_q[157] : 
                                (N147)? btb_q[222] : 
                                (N149)? btb_q[287] : 
                                (N151)? btb_q[352] : 
                                (N153)? btb_q[417] : 
                                (N155)? btb_q[482] : 
                                (N157)? btb_q[547] : 
                                (N159)? btb_q[612] : 
                                (N161)? btb_q[677] : 
                                (N163)? btb_q[742] : 
                                (N165)? btb_q[807] : 
                                (N167)? btb_q[872] : 
                                (N169)? btb_q[937] : 
                                (N171)? btb_q[1002] : 
                                (N173)? btb_q[1067] : 
                                (N175)? btb_q[1132] : 
                                (N177)? btb_q[1197] : 
                                (N179)? btb_q[1262] : 
                                (N181)? btb_q[1327] : 
                                (N183)? btb_q[1392] : 
                                (N185)? btb_q[1457] : 
                                (N187)? btb_q[1522] : 
                                (N189)? btb_q[1587] : 
                                (N191)? btb_q[1652] : 
                                (N193)? btb_q[1717] : 
                                (N195)? btb_q[1782] : 
                                (N197)? btb_q[1847] : 
                                (N199)? btb_q[1912] : 
                                (N201)? btb_q[1977] : 
                                (N203)? btb_q[2042] : 
                                (N142)? btb_q[2107] : 
                                (N144)? btb_q[2172] : 
                                (N146)? btb_q[2237] : 
                                (N148)? btb_q[2302] : 
                                (N150)? btb_q[2367] : 
                                (N152)? btb_q[2432] : 
                                (N154)? btb_q[2497] : 
                                (N156)? btb_q[2562] : 
                                (N158)? btb_q[2627] : 
                                (N160)? btb_q[2692] : 
                                (N162)? btb_q[2757] : 
                                (N164)? btb_q[2822] : 
                                (N166)? btb_q[2887] : 
                                (N168)? btb_q[2952] : 
                                (N170)? btb_q[3017] : 
                                (N172)? btb_q[3082] : 
                                (N174)? btb_q[3147] : 
                                (N176)? btb_q[3212] : 
                                (N178)? btb_q[3277] : 
                                (N180)? btb_q[3342] : 
                                (N182)? btb_q[3407] : 
                                (N184)? btb_q[3472] : 
                                (N186)? btb_q[3537] : 
                                (N188)? btb_q[3602] : 
                                (N190)? btb_q[3667] : 
                                (N192)? btb_q[3732] : 
                                (N194)? btb_q[3797] : 
                                (N196)? btb_q[3862] : 
                                (N198)? btb_q[3927] : 
                                (N200)? btb_q[3992] : 
                                (N202)? btb_q[4057] : 
                                (N204)? btb_q[4122] : 1'b0;
  assign btb_prediction_o[26] = (N141)? btb_q[26] : 
                                (N143)? btb_q[91] : 
                                (N145)? btb_q[156] : 
                                (N147)? btb_q[221] : 
                                (N149)? btb_q[286] : 
                                (N151)? btb_q[351] : 
                                (N153)? btb_q[416] : 
                                (N155)? btb_q[481] : 
                                (N157)? btb_q[546] : 
                                (N159)? btb_q[611] : 
                                (N161)? btb_q[676] : 
                                (N163)? btb_q[741] : 
                                (N165)? btb_q[806] : 
                                (N167)? btb_q[871] : 
                                (N169)? btb_q[936] : 
                                (N171)? btb_q[1001] : 
                                (N173)? btb_q[1066] : 
                                (N175)? btb_q[1131] : 
                                (N177)? btb_q[1196] : 
                                (N179)? btb_q[1261] : 
                                (N181)? btb_q[1326] : 
                                (N183)? btb_q[1391] : 
                                (N185)? btb_q[1456] : 
                                (N187)? btb_q[1521] : 
                                (N189)? btb_q[1586] : 
                                (N191)? btb_q[1651] : 
                                (N193)? btb_q[1716] : 
                                (N195)? btb_q[1781] : 
                                (N197)? btb_q[1846] : 
                                (N199)? btb_q[1911] : 
                                (N201)? btb_q[1976] : 
                                (N203)? btb_q[2041] : 
                                (N142)? btb_q[2106] : 
                                (N144)? btb_q[2171] : 
                                (N146)? btb_q[2236] : 
                                (N148)? btb_q[2301] : 
                                (N150)? btb_q[2366] : 
                                (N152)? btb_q[2431] : 
                                (N154)? btb_q[2496] : 
                                (N156)? btb_q[2561] : 
                                (N158)? btb_q[2626] : 
                                (N160)? btb_q[2691] : 
                                (N162)? btb_q[2756] : 
                                (N164)? btb_q[2821] : 
                                (N166)? btb_q[2886] : 
                                (N168)? btb_q[2951] : 
                                (N170)? btb_q[3016] : 
                                (N172)? btb_q[3081] : 
                                (N174)? btb_q[3146] : 
                                (N176)? btb_q[3211] : 
                                (N178)? btb_q[3276] : 
                                (N180)? btb_q[3341] : 
                                (N182)? btb_q[3406] : 
                                (N184)? btb_q[3471] : 
                                (N186)? btb_q[3536] : 
                                (N188)? btb_q[3601] : 
                                (N190)? btb_q[3666] : 
                                (N192)? btb_q[3731] : 
                                (N194)? btb_q[3796] : 
                                (N196)? btb_q[3861] : 
                                (N198)? btb_q[3926] : 
                                (N200)? btb_q[3991] : 
                                (N202)? btb_q[4056] : 
                                (N204)? btb_q[4121] : 1'b0;
  assign btb_prediction_o[25] = (N141)? btb_q[25] : 
                                (N143)? btb_q[90] : 
                                (N145)? btb_q[155] : 
                                (N147)? btb_q[220] : 
                                (N149)? btb_q[285] : 
                                (N151)? btb_q[350] : 
                                (N153)? btb_q[415] : 
                                (N155)? btb_q[480] : 
                                (N157)? btb_q[545] : 
                                (N159)? btb_q[610] : 
                                (N161)? btb_q[675] : 
                                (N163)? btb_q[740] : 
                                (N165)? btb_q[805] : 
                                (N167)? btb_q[870] : 
                                (N169)? btb_q[935] : 
                                (N171)? btb_q[1000] : 
                                (N173)? btb_q[1065] : 
                                (N175)? btb_q[1130] : 
                                (N177)? btb_q[1195] : 
                                (N179)? btb_q[1260] : 
                                (N181)? btb_q[1325] : 
                                (N183)? btb_q[1390] : 
                                (N185)? btb_q[1455] : 
                                (N187)? btb_q[1520] : 
                                (N189)? btb_q[1585] : 
                                (N191)? btb_q[1650] : 
                                (N193)? btb_q[1715] : 
                                (N195)? btb_q[1780] : 
                                (N197)? btb_q[1845] : 
                                (N199)? btb_q[1910] : 
                                (N201)? btb_q[1975] : 
                                (N203)? btb_q[2040] : 
                                (N142)? btb_q[2105] : 
                                (N144)? btb_q[2170] : 
                                (N146)? btb_q[2235] : 
                                (N148)? btb_q[2300] : 
                                (N150)? btb_q[2365] : 
                                (N152)? btb_q[2430] : 
                                (N154)? btb_q[2495] : 
                                (N156)? btb_q[2560] : 
                                (N158)? btb_q[2625] : 
                                (N160)? btb_q[2690] : 
                                (N162)? btb_q[2755] : 
                                (N164)? btb_q[2820] : 
                                (N166)? btb_q[2885] : 
                                (N168)? btb_q[2950] : 
                                (N170)? btb_q[3015] : 
                                (N172)? btb_q[3080] : 
                                (N174)? btb_q[3145] : 
                                (N176)? btb_q[3210] : 
                                (N178)? btb_q[3275] : 
                                (N180)? btb_q[3340] : 
                                (N182)? btb_q[3405] : 
                                (N184)? btb_q[3470] : 
                                (N186)? btb_q[3535] : 
                                (N188)? btb_q[3600] : 
                                (N190)? btb_q[3665] : 
                                (N192)? btb_q[3730] : 
                                (N194)? btb_q[3795] : 
                                (N196)? btb_q[3860] : 
                                (N198)? btb_q[3925] : 
                                (N200)? btb_q[3990] : 
                                (N202)? btb_q[4055] : 
                                (N204)? btb_q[4120] : 1'b0;
  assign btb_prediction_o[24] = (N141)? btb_q[24] : 
                                (N143)? btb_q[89] : 
                                (N145)? btb_q[154] : 
                                (N147)? btb_q[219] : 
                                (N149)? btb_q[284] : 
                                (N151)? btb_q[349] : 
                                (N153)? btb_q[414] : 
                                (N155)? btb_q[479] : 
                                (N157)? btb_q[544] : 
                                (N159)? btb_q[609] : 
                                (N161)? btb_q[674] : 
                                (N163)? btb_q[739] : 
                                (N165)? btb_q[804] : 
                                (N167)? btb_q[869] : 
                                (N169)? btb_q[934] : 
                                (N171)? btb_q[999] : 
                                (N173)? btb_q[1064] : 
                                (N175)? btb_q[1129] : 
                                (N177)? btb_q[1194] : 
                                (N179)? btb_q[1259] : 
                                (N181)? btb_q[1324] : 
                                (N183)? btb_q[1389] : 
                                (N185)? btb_q[1454] : 
                                (N187)? btb_q[1519] : 
                                (N189)? btb_q[1584] : 
                                (N191)? btb_q[1649] : 
                                (N193)? btb_q[1714] : 
                                (N195)? btb_q[1779] : 
                                (N197)? btb_q[1844] : 
                                (N199)? btb_q[1909] : 
                                (N201)? btb_q[1974] : 
                                (N203)? btb_q[2039] : 
                                (N142)? btb_q[2104] : 
                                (N144)? btb_q[2169] : 
                                (N146)? btb_q[2234] : 
                                (N148)? btb_q[2299] : 
                                (N150)? btb_q[2364] : 
                                (N152)? btb_q[2429] : 
                                (N154)? btb_q[2494] : 
                                (N156)? btb_q[2559] : 
                                (N158)? btb_q[2624] : 
                                (N160)? btb_q[2689] : 
                                (N162)? btb_q[2754] : 
                                (N164)? btb_q[2819] : 
                                (N166)? btb_q[2884] : 
                                (N168)? btb_q[2949] : 
                                (N170)? btb_q[3014] : 
                                (N172)? btb_q[3079] : 
                                (N174)? btb_q[3144] : 
                                (N176)? btb_q[3209] : 
                                (N178)? btb_q[3274] : 
                                (N180)? btb_q[3339] : 
                                (N182)? btb_q[3404] : 
                                (N184)? btb_q[3469] : 
                                (N186)? btb_q[3534] : 
                                (N188)? btb_q[3599] : 
                                (N190)? btb_q[3664] : 
                                (N192)? btb_q[3729] : 
                                (N194)? btb_q[3794] : 
                                (N196)? btb_q[3859] : 
                                (N198)? btb_q[3924] : 
                                (N200)? btb_q[3989] : 
                                (N202)? btb_q[4054] : 
                                (N204)? btb_q[4119] : 1'b0;
  assign btb_prediction_o[23] = (N141)? btb_q[23] : 
                                (N143)? btb_q[88] : 
                                (N145)? btb_q[153] : 
                                (N147)? btb_q[218] : 
                                (N149)? btb_q[283] : 
                                (N151)? btb_q[348] : 
                                (N153)? btb_q[413] : 
                                (N155)? btb_q[478] : 
                                (N157)? btb_q[543] : 
                                (N159)? btb_q[608] : 
                                (N161)? btb_q[673] : 
                                (N163)? btb_q[738] : 
                                (N165)? btb_q[803] : 
                                (N167)? btb_q[868] : 
                                (N169)? btb_q[933] : 
                                (N171)? btb_q[998] : 
                                (N173)? btb_q[1063] : 
                                (N175)? btb_q[1128] : 
                                (N177)? btb_q[1193] : 
                                (N179)? btb_q[1258] : 
                                (N181)? btb_q[1323] : 
                                (N183)? btb_q[1388] : 
                                (N185)? btb_q[1453] : 
                                (N187)? btb_q[1518] : 
                                (N189)? btb_q[1583] : 
                                (N191)? btb_q[1648] : 
                                (N193)? btb_q[1713] : 
                                (N195)? btb_q[1778] : 
                                (N197)? btb_q[1843] : 
                                (N199)? btb_q[1908] : 
                                (N201)? btb_q[1973] : 
                                (N203)? btb_q[2038] : 
                                (N142)? btb_q[2103] : 
                                (N144)? btb_q[2168] : 
                                (N146)? btb_q[2233] : 
                                (N148)? btb_q[2298] : 
                                (N150)? btb_q[2363] : 
                                (N152)? btb_q[2428] : 
                                (N154)? btb_q[2493] : 
                                (N156)? btb_q[2558] : 
                                (N158)? btb_q[2623] : 
                                (N160)? btb_q[2688] : 
                                (N162)? btb_q[2753] : 
                                (N164)? btb_q[2818] : 
                                (N166)? btb_q[2883] : 
                                (N168)? btb_q[2948] : 
                                (N170)? btb_q[3013] : 
                                (N172)? btb_q[3078] : 
                                (N174)? btb_q[3143] : 
                                (N176)? btb_q[3208] : 
                                (N178)? btb_q[3273] : 
                                (N180)? btb_q[3338] : 
                                (N182)? btb_q[3403] : 
                                (N184)? btb_q[3468] : 
                                (N186)? btb_q[3533] : 
                                (N188)? btb_q[3598] : 
                                (N190)? btb_q[3663] : 
                                (N192)? btb_q[3728] : 
                                (N194)? btb_q[3793] : 
                                (N196)? btb_q[3858] : 
                                (N198)? btb_q[3923] : 
                                (N200)? btb_q[3988] : 
                                (N202)? btb_q[4053] : 
                                (N204)? btb_q[4118] : 1'b0;
  assign btb_prediction_o[22] = (N141)? btb_q[22] : 
                                (N143)? btb_q[87] : 
                                (N145)? btb_q[152] : 
                                (N147)? btb_q[217] : 
                                (N149)? btb_q[282] : 
                                (N151)? btb_q[347] : 
                                (N153)? btb_q[412] : 
                                (N155)? btb_q[477] : 
                                (N157)? btb_q[542] : 
                                (N159)? btb_q[607] : 
                                (N161)? btb_q[672] : 
                                (N163)? btb_q[737] : 
                                (N165)? btb_q[802] : 
                                (N167)? btb_q[867] : 
                                (N169)? btb_q[932] : 
                                (N171)? btb_q[997] : 
                                (N173)? btb_q[1062] : 
                                (N175)? btb_q[1127] : 
                                (N177)? btb_q[1192] : 
                                (N179)? btb_q[1257] : 
                                (N181)? btb_q[1322] : 
                                (N183)? btb_q[1387] : 
                                (N185)? btb_q[1452] : 
                                (N187)? btb_q[1517] : 
                                (N189)? btb_q[1582] : 
                                (N191)? btb_q[1647] : 
                                (N193)? btb_q[1712] : 
                                (N195)? btb_q[1777] : 
                                (N197)? btb_q[1842] : 
                                (N199)? btb_q[1907] : 
                                (N201)? btb_q[1972] : 
                                (N203)? btb_q[2037] : 
                                (N142)? btb_q[2102] : 
                                (N144)? btb_q[2167] : 
                                (N146)? btb_q[2232] : 
                                (N148)? btb_q[2297] : 
                                (N150)? btb_q[2362] : 
                                (N152)? btb_q[2427] : 
                                (N154)? btb_q[2492] : 
                                (N156)? btb_q[2557] : 
                                (N158)? btb_q[2622] : 
                                (N160)? btb_q[2687] : 
                                (N162)? btb_q[2752] : 
                                (N164)? btb_q[2817] : 
                                (N166)? btb_q[2882] : 
                                (N168)? btb_q[2947] : 
                                (N170)? btb_q[3012] : 
                                (N172)? btb_q[3077] : 
                                (N174)? btb_q[3142] : 
                                (N176)? btb_q[3207] : 
                                (N178)? btb_q[3272] : 
                                (N180)? btb_q[3337] : 
                                (N182)? btb_q[3402] : 
                                (N184)? btb_q[3467] : 
                                (N186)? btb_q[3532] : 
                                (N188)? btb_q[3597] : 
                                (N190)? btb_q[3662] : 
                                (N192)? btb_q[3727] : 
                                (N194)? btb_q[3792] : 
                                (N196)? btb_q[3857] : 
                                (N198)? btb_q[3922] : 
                                (N200)? btb_q[3987] : 
                                (N202)? btb_q[4052] : 
                                (N204)? btb_q[4117] : 1'b0;
  assign btb_prediction_o[21] = (N141)? btb_q[21] : 
                                (N143)? btb_q[86] : 
                                (N145)? btb_q[151] : 
                                (N147)? btb_q[216] : 
                                (N149)? btb_q[281] : 
                                (N151)? btb_q[346] : 
                                (N153)? btb_q[411] : 
                                (N155)? btb_q[476] : 
                                (N157)? btb_q[541] : 
                                (N159)? btb_q[606] : 
                                (N161)? btb_q[671] : 
                                (N163)? btb_q[736] : 
                                (N165)? btb_q[801] : 
                                (N167)? btb_q[866] : 
                                (N169)? btb_q[931] : 
                                (N171)? btb_q[996] : 
                                (N173)? btb_q[1061] : 
                                (N175)? btb_q[1126] : 
                                (N177)? btb_q[1191] : 
                                (N179)? btb_q[1256] : 
                                (N181)? btb_q[1321] : 
                                (N183)? btb_q[1386] : 
                                (N185)? btb_q[1451] : 
                                (N187)? btb_q[1516] : 
                                (N189)? btb_q[1581] : 
                                (N191)? btb_q[1646] : 
                                (N193)? btb_q[1711] : 
                                (N195)? btb_q[1776] : 
                                (N197)? btb_q[1841] : 
                                (N199)? btb_q[1906] : 
                                (N201)? btb_q[1971] : 
                                (N203)? btb_q[2036] : 
                                (N142)? btb_q[2101] : 
                                (N144)? btb_q[2166] : 
                                (N146)? btb_q[2231] : 
                                (N148)? btb_q[2296] : 
                                (N150)? btb_q[2361] : 
                                (N152)? btb_q[2426] : 
                                (N154)? btb_q[2491] : 
                                (N156)? btb_q[2556] : 
                                (N158)? btb_q[2621] : 
                                (N160)? btb_q[2686] : 
                                (N162)? btb_q[2751] : 
                                (N164)? btb_q[2816] : 
                                (N166)? btb_q[2881] : 
                                (N168)? btb_q[2946] : 
                                (N170)? btb_q[3011] : 
                                (N172)? btb_q[3076] : 
                                (N174)? btb_q[3141] : 
                                (N176)? btb_q[3206] : 
                                (N178)? btb_q[3271] : 
                                (N180)? btb_q[3336] : 
                                (N182)? btb_q[3401] : 
                                (N184)? btb_q[3466] : 
                                (N186)? btb_q[3531] : 
                                (N188)? btb_q[3596] : 
                                (N190)? btb_q[3661] : 
                                (N192)? btb_q[3726] : 
                                (N194)? btb_q[3791] : 
                                (N196)? btb_q[3856] : 
                                (N198)? btb_q[3921] : 
                                (N200)? btb_q[3986] : 
                                (N202)? btb_q[4051] : 
                                (N204)? btb_q[4116] : 1'b0;
  assign btb_prediction_o[20] = (N141)? btb_q[20] : 
                                (N143)? btb_q[85] : 
                                (N145)? btb_q[150] : 
                                (N147)? btb_q[215] : 
                                (N149)? btb_q[280] : 
                                (N151)? btb_q[345] : 
                                (N153)? btb_q[410] : 
                                (N155)? btb_q[475] : 
                                (N157)? btb_q[540] : 
                                (N159)? btb_q[605] : 
                                (N161)? btb_q[670] : 
                                (N163)? btb_q[735] : 
                                (N165)? btb_q[800] : 
                                (N167)? btb_q[865] : 
                                (N169)? btb_q[930] : 
                                (N171)? btb_q[995] : 
                                (N173)? btb_q[1060] : 
                                (N175)? btb_q[1125] : 
                                (N177)? btb_q[1190] : 
                                (N179)? btb_q[1255] : 
                                (N181)? btb_q[1320] : 
                                (N183)? btb_q[1385] : 
                                (N185)? btb_q[1450] : 
                                (N187)? btb_q[1515] : 
                                (N189)? btb_q[1580] : 
                                (N191)? btb_q[1645] : 
                                (N193)? btb_q[1710] : 
                                (N195)? btb_q[1775] : 
                                (N197)? btb_q[1840] : 
                                (N199)? btb_q[1905] : 
                                (N201)? btb_q[1970] : 
                                (N203)? btb_q[2035] : 
                                (N142)? btb_q[2100] : 
                                (N144)? btb_q[2165] : 
                                (N146)? btb_q[2230] : 
                                (N148)? btb_q[2295] : 
                                (N150)? btb_q[2360] : 
                                (N152)? btb_q[2425] : 
                                (N154)? btb_q[2490] : 
                                (N156)? btb_q[2555] : 
                                (N158)? btb_q[2620] : 
                                (N160)? btb_q[2685] : 
                                (N162)? btb_q[2750] : 
                                (N164)? btb_q[2815] : 
                                (N166)? btb_q[2880] : 
                                (N168)? btb_q[2945] : 
                                (N170)? btb_q[3010] : 
                                (N172)? btb_q[3075] : 
                                (N174)? btb_q[3140] : 
                                (N176)? btb_q[3205] : 
                                (N178)? btb_q[3270] : 
                                (N180)? btb_q[3335] : 
                                (N182)? btb_q[3400] : 
                                (N184)? btb_q[3465] : 
                                (N186)? btb_q[3530] : 
                                (N188)? btb_q[3595] : 
                                (N190)? btb_q[3660] : 
                                (N192)? btb_q[3725] : 
                                (N194)? btb_q[3790] : 
                                (N196)? btb_q[3855] : 
                                (N198)? btb_q[3920] : 
                                (N200)? btb_q[3985] : 
                                (N202)? btb_q[4050] : 
                                (N204)? btb_q[4115] : 1'b0;
  assign btb_prediction_o[19] = (N141)? btb_q[19] : 
                                (N143)? btb_q[84] : 
                                (N145)? btb_q[149] : 
                                (N147)? btb_q[214] : 
                                (N149)? btb_q[279] : 
                                (N151)? btb_q[344] : 
                                (N153)? btb_q[409] : 
                                (N155)? btb_q[474] : 
                                (N157)? btb_q[539] : 
                                (N159)? btb_q[604] : 
                                (N161)? btb_q[669] : 
                                (N163)? btb_q[734] : 
                                (N165)? btb_q[799] : 
                                (N167)? btb_q[864] : 
                                (N169)? btb_q[929] : 
                                (N171)? btb_q[994] : 
                                (N173)? btb_q[1059] : 
                                (N175)? btb_q[1124] : 
                                (N177)? btb_q[1189] : 
                                (N179)? btb_q[1254] : 
                                (N181)? btb_q[1319] : 
                                (N183)? btb_q[1384] : 
                                (N185)? btb_q[1449] : 
                                (N187)? btb_q[1514] : 
                                (N189)? btb_q[1579] : 
                                (N191)? btb_q[1644] : 
                                (N193)? btb_q[1709] : 
                                (N195)? btb_q[1774] : 
                                (N197)? btb_q[1839] : 
                                (N199)? btb_q[1904] : 
                                (N201)? btb_q[1969] : 
                                (N203)? btb_q[2034] : 
                                (N142)? btb_q[2099] : 
                                (N144)? btb_q[2164] : 
                                (N146)? btb_q[2229] : 
                                (N148)? btb_q[2294] : 
                                (N150)? btb_q[2359] : 
                                (N152)? btb_q[2424] : 
                                (N154)? btb_q[2489] : 
                                (N156)? btb_q[2554] : 
                                (N158)? btb_q[2619] : 
                                (N160)? btb_q[2684] : 
                                (N162)? btb_q[2749] : 
                                (N164)? btb_q[2814] : 
                                (N166)? btb_q[2879] : 
                                (N168)? btb_q[2944] : 
                                (N170)? btb_q[3009] : 
                                (N172)? btb_q[3074] : 
                                (N174)? btb_q[3139] : 
                                (N176)? btb_q[3204] : 
                                (N178)? btb_q[3269] : 
                                (N180)? btb_q[3334] : 
                                (N182)? btb_q[3399] : 
                                (N184)? btb_q[3464] : 
                                (N186)? btb_q[3529] : 
                                (N188)? btb_q[3594] : 
                                (N190)? btb_q[3659] : 
                                (N192)? btb_q[3724] : 
                                (N194)? btb_q[3789] : 
                                (N196)? btb_q[3854] : 
                                (N198)? btb_q[3919] : 
                                (N200)? btb_q[3984] : 
                                (N202)? btb_q[4049] : 
                                (N204)? btb_q[4114] : 1'b0;
  assign btb_prediction_o[18] = (N141)? btb_q[18] : 
                                (N143)? btb_q[83] : 
                                (N145)? btb_q[148] : 
                                (N147)? btb_q[213] : 
                                (N149)? btb_q[278] : 
                                (N151)? btb_q[343] : 
                                (N153)? btb_q[408] : 
                                (N155)? btb_q[473] : 
                                (N157)? btb_q[538] : 
                                (N159)? btb_q[603] : 
                                (N161)? btb_q[668] : 
                                (N163)? btb_q[733] : 
                                (N165)? btb_q[798] : 
                                (N167)? btb_q[863] : 
                                (N169)? btb_q[928] : 
                                (N171)? btb_q[993] : 
                                (N173)? btb_q[1058] : 
                                (N175)? btb_q[1123] : 
                                (N177)? btb_q[1188] : 
                                (N179)? btb_q[1253] : 
                                (N181)? btb_q[1318] : 
                                (N183)? btb_q[1383] : 
                                (N185)? btb_q[1448] : 
                                (N187)? btb_q[1513] : 
                                (N189)? btb_q[1578] : 
                                (N191)? btb_q[1643] : 
                                (N193)? btb_q[1708] : 
                                (N195)? btb_q[1773] : 
                                (N197)? btb_q[1838] : 
                                (N199)? btb_q[1903] : 
                                (N201)? btb_q[1968] : 
                                (N203)? btb_q[2033] : 
                                (N142)? btb_q[2098] : 
                                (N144)? btb_q[2163] : 
                                (N146)? btb_q[2228] : 
                                (N148)? btb_q[2293] : 
                                (N150)? btb_q[2358] : 
                                (N152)? btb_q[2423] : 
                                (N154)? btb_q[2488] : 
                                (N156)? btb_q[2553] : 
                                (N158)? btb_q[2618] : 
                                (N160)? btb_q[2683] : 
                                (N162)? btb_q[2748] : 
                                (N164)? btb_q[2813] : 
                                (N166)? btb_q[2878] : 
                                (N168)? btb_q[2943] : 
                                (N170)? btb_q[3008] : 
                                (N172)? btb_q[3073] : 
                                (N174)? btb_q[3138] : 
                                (N176)? btb_q[3203] : 
                                (N178)? btb_q[3268] : 
                                (N180)? btb_q[3333] : 
                                (N182)? btb_q[3398] : 
                                (N184)? btb_q[3463] : 
                                (N186)? btb_q[3528] : 
                                (N188)? btb_q[3593] : 
                                (N190)? btb_q[3658] : 
                                (N192)? btb_q[3723] : 
                                (N194)? btb_q[3788] : 
                                (N196)? btb_q[3853] : 
                                (N198)? btb_q[3918] : 
                                (N200)? btb_q[3983] : 
                                (N202)? btb_q[4048] : 
                                (N204)? btb_q[4113] : 1'b0;
  assign btb_prediction_o[17] = (N141)? btb_q[17] : 
                                (N143)? btb_q[82] : 
                                (N145)? btb_q[147] : 
                                (N147)? btb_q[212] : 
                                (N149)? btb_q[277] : 
                                (N151)? btb_q[342] : 
                                (N153)? btb_q[407] : 
                                (N155)? btb_q[472] : 
                                (N157)? btb_q[537] : 
                                (N159)? btb_q[602] : 
                                (N161)? btb_q[667] : 
                                (N163)? btb_q[732] : 
                                (N165)? btb_q[797] : 
                                (N167)? btb_q[862] : 
                                (N169)? btb_q[927] : 
                                (N171)? btb_q[992] : 
                                (N173)? btb_q[1057] : 
                                (N175)? btb_q[1122] : 
                                (N177)? btb_q[1187] : 
                                (N179)? btb_q[1252] : 
                                (N181)? btb_q[1317] : 
                                (N183)? btb_q[1382] : 
                                (N185)? btb_q[1447] : 
                                (N187)? btb_q[1512] : 
                                (N189)? btb_q[1577] : 
                                (N191)? btb_q[1642] : 
                                (N193)? btb_q[1707] : 
                                (N195)? btb_q[1772] : 
                                (N197)? btb_q[1837] : 
                                (N199)? btb_q[1902] : 
                                (N201)? btb_q[1967] : 
                                (N203)? btb_q[2032] : 
                                (N142)? btb_q[2097] : 
                                (N144)? btb_q[2162] : 
                                (N146)? btb_q[2227] : 
                                (N148)? btb_q[2292] : 
                                (N150)? btb_q[2357] : 
                                (N152)? btb_q[2422] : 
                                (N154)? btb_q[2487] : 
                                (N156)? btb_q[2552] : 
                                (N158)? btb_q[2617] : 
                                (N160)? btb_q[2682] : 
                                (N162)? btb_q[2747] : 
                                (N164)? btb_q[2812] : 
                                (N166)? btb_q[2877] : 
                                (N168)? btb_q[2942] : 
                                (N170)? btb_q[3007] : 
                                (N172)? btb_q[3072] : 
                                (N174)? btb_q[3137] : 
                                (N176)? btb_q[3202] : 
                                (N178)? btb_q[3267] : 
                                (N180)? btb_q[3332] : 
                                (N182)? btb_q[3397] : 
                                (N184)? btb_q[3462] : 
                                (N186)? btb_q[3527] : 
                                (N188)? btb_q[3592] : 
                                (N190)? btb_q[3657] : 
                                (N192)? btb_q[3722] : 
                                (N194)? btb_q[3787] : 
                                (N196)? btb_q[3852] : 
                                (N198)? btb_q[3917] : 
                                (N200)? btb_q[3982] : 
                                (N202)? btb_q[4047] : 
                                (N204)? btb_q[4112] : 1'b0;
  assign btb_prediction_o[16] = (N141)? btb_q[16] : 
                                (N143)? btb_q[81] : 
                                (N145)? btb_q[146] : 
                                (N147)? btb_q[211] : 
                                (N149)? btb_q[276] : 
                                (N151)? btb_q[341] : 
                                (N153)? btb_q[406] : 
                                (N155)? btb_q[471] : 
                                (N157)? btb_q[536] : 
                                (N159)? btb_q[601] : 
                                (N161)? btb_q[666] : 
                                (N163)? btb_q[731] : 
                                (N165)? btb_q[796] : 
                                (N167)? btb_q[861] : 
                                (N169)? btb_q[926] : 
                                (N171)? btb_q[991] : 
                                (N173)? btb_q[1056] : 
                                (N175)? btb_q[1121] : 
                                (N177)? btb_q[1186] : 
                                (N179)? btb_q[1251] : 
                                (N181)? btb_q[1316] : 
                                (N183)? btb_q[1381] : 
                                (N185)? btb_q[1446] : 
                                (N187)? btb_q[1511] : 
                                (N189)? btb_q[1576] : 
                                (N191)? btb_q[1641] : 
                                (N193)? btb_q[1706] : 
                                (N195)? btb_q[1771] : 
                                (N197)? btb_q[1836] : 
                                (N199)? btb_q[1901] : 
                                (N201)? btb_q[1966] : 
                                (N203)? btb_q[2031] : 
                                (N142)? btb_q[2096] : 
                                (N144)? btb_q[2161] : 
                                (N146)? btb_q[2226] : 
                                (N148)? btb_q[2291] : 
                                (N150)? btb_q[2356] : 
                                (N152)? btb_q[2421] : 
                                (N154)? btb_q[2486] : 
                                (N156)? btb_q[2551] : 
                                (N158)? btb_q[2616] : 
                                (N160)? btb_q[2681] : 
                                (N162)? btb_q[2746] : 
                                (N164)? btb_q[2811] : 
                                (N166)? btb_q[2876] : 
                                (N168)? btb_q[2941] : 
                                (N170)? btb_q[3006] : 
                                (N172)? btb_q[3071] : 
                                (N174)? btb_q[3136] : 
                                (N176)? btb_q[3201] : 
                                (N178)? btb_q[3266] : 
                                (N180)? btb_q[3331] : 
                                (N182)? btb_q[3396] : 
                                (N184)? btb_q[3461] : 
                                (N186)? btb_q[3526] : 
                                (N188)? btb_q[3591] : 
                                (N190)? btb_q[3656] : 
                                (N192)? btb_q[3721] : 
                                (N194)? btb_q[3786] : 
                                (N196)? btb_q[3851] : 
                                (N198)? btb_q[3916] : 
                                (N200)? btb_q[3981] : 
                                (N202)? btb_q[4046] : 
                                (N204)? btb_q[4111] : 1'b0;
  assign btb_prediction_o[15] = (N141)? btb_q[15] : 
                                (N143)? btb_q[80] : 
                                (N145)? btb_q[145] : 
                                (N147)? btb_q[210] : 
                                (N149)? btb_q[275] : 
                                (N151)? btb_q[340] : 
                                (N153)? btb_q[405] : 
                                (N155)? btb_q[470] : 
                                (N157)? btb_q[535] : 
                                (N159)? btb_q[600] : 
                                (N161)? btb_q[665] : 
                                (N163)? btb_q[730] : 
                                (N165)? btb_q[795] : 
                                (N167)? btb_q[860] : 
                                (N169)? btb_q[925] : 
                                (N171)? btb_q[990] : 
                                (N173)? btb_q[1055] : 
                                (N175)? btb_q[1120] : 
                                (N177)? btb_q[1185] : 
                                (N179)? btb_q[1250] : 
                                (N181)? btb_q[1315] : 
                                (N183)? btb_q[1380] : 
                                (N185)? btb_q[1445] : 
                                (N187)? btb_q[1510] : 
                                (N189)? btb_q[1575] : 
                                (N191)? btb_q[1640] : 
                                (N193)? btb_q[1705] : 
                                (N195)? btb_q[1770] : 
                                (N197)? btb_q[1835] : 
                                (N199)? btb_q[1900] : 
                                (N201)? btb_q[1965] : 
                                (N203)? btb_q[2030] : 
                                (N142)? btb_q[2095] : 
                                (N144)? btb_q[2160] : 
                                (N146)? btb_q[2225] : 
                                (N148)? btb_q[2290] : 
                                (N150)? btb_q[2355] : 
                                (N152)? btb_q[2420] : 
                                (N154)? btb_q[2485] : 
                                (N156)? btb_q[2550] : 
                                (N158)? btb_q[2615] : 
                                (N160)? btb_q[2680] : 
                                (N162)? btb_q[2745] : 
                                (N164)? btb_q[2810] : 
                                (N166)? btb_q[2875] : 
                                (N168)? btb_q[2940] : 
                                (N170)? btb_q[3005] : 
                                (N172)? btb_q[3070] : 
                                (N174)? btb_q[3135] : 
                                (N176)? btb_q[3200] : 
                                (N178)? btb_q[3265] : 
                                (N180)? btb_q[3330] : 
                                (N182)? btb_q[3395] : 
                                (N184)? btb_q[3460] : 
                                (N186)? btb_q[3525] : 
                                (N188)? btb_q[3590] : 
                                (N190)? btb_q[3655] : 
                                (N192)? btb_q[3720] : 
                                (N194)? btb_q[3785] : 
                                (N196)? btb_q[3850] : 
                                (N198)? btb_q[3915] : 
                                (N200)? btb_q[3980] : 
                                (N202)? btb_q[4045] : 
                                (N204)? btb_q[4110] : 1'b0;
  assign btb_prediction_o[14] = (N141)? btb_q[14] : 
                                (N143)? btb_q[79] : 
                                (N145)? btb_q[144] : 
                                (N147)? btb_q[209] : 
                                (N149)? btb_q[274] : 
                                (N151)? btb_q[339] : 
                                (N153)? btb_q[404] : 
                                (N155)? btb_q[469] : 
                                (N157)? btb_q[534] : 
                                (N159)? btb_q[599] : 
                                (N161)? btb_q[664] : 
                                (N163)? btb_q[729] : 
                                (N165)? btb_q[794] : 
                                (N167)? btb_q[859] : 
                                (N169)? btb_q[924] : 
                                (N171)? btb_q[989] : 
                                (N173)? btb_q[1054] : 
                                (N175)? btb_q[1119] : 
                                (N177)? btb_q[1184] : 
                                (N179)? btb_q[1249] : 
                                (N181)? btb_q[1314] : 
                                (N183)? btb_q[1379] : 
                                (N185)? btb_q[1444] : 
                                (N187)? btb_q[1509] : 
                                (N189)? btb_q[1574] : 
                                (N191)? btb_q[1639] : 
                                (N193)? btb_q[1704] : 
                                (N195)? btb_q[1769] : 
                                (N197)? btb_q[1834] : 
                                (N199)? btb_q[1899] : 
                                (N201)? btb_q[1964] : 
                                (N203)? btb_q[2029] : 
                                (N142)? btb_q[2094] : 
                                (N144)? btb_q[2159] : 
                                (N146)? btb_q[2224] : 
                                (N148)? btb_q[2289] : 
                                (N150)? btb_q[2354] : 
                                (N152)? btb_q[2419] : 
                                (N154)? btb_q[2484] : 
                                (N156)? btb_q[2549] : 
                                (N158)? btb_q[2614] : 
                                (N160)? btb_q[2679] : 
                                (N162)? btb_q[2744] : 
                                (N164)? btb_q[2809] : 
                                (N166)? btb_q[2874] : 
                                (N168)? btb_q[2939] : 
                                (N170)? btb_q[3004] : 
                                (N172)? btb_q[3069] : 
                                (N174)? btb_q[3134] : 
                                (N176)? btb_q[3199] : 
                                (N178)? btb_q[3264] : 
                                (N180)? btb_q[3329] : 
                                (N182)? btb_q[3394] : 
                                (N184)? btb_q[3459] : 
                                (N186)? btb_q[3524] : 
                                (N188)? btb_q[3589] : 
                                (N190)? btb_q[3654] : 
                                (N192)? btb_q[3719] : 
                                (N194)? btb_q[3784] : 
                                (N196)? btb_q[3849] : 
                                (N198)? btb_q[3914] : 
                                (N200)? btb_q[3979] : 
                                (N202)? btb_q[4044] : 
                                (N204)? btb_q[4109] : 1'b0;
  assign btb_prediction_o[13] = (N141)? btb_q[13] : 
                                (N143)? btb_q[78] : 
                                (N145)? btb_q[143] : 
                                (N147)? btb_q[208] : 
                                (N149)? btb_q[273] : 
                                (N151)? btb_q[338] : 
                                (N153)? btb_q[403] : 
                                (N155)? btb_q[468] : 
                                (N157)? btb_q[533] : 
                                (N159)? btb_q[598] : 
                                (N161)? btb_q[663] : 
                                (N163)? btb_q[728] : 
                                (N165)? btb_q[793] : 
                                (N167)? btb_q[858] : 
                                (N169)? btb_q[923] : 
                                (N171)? btb_q[988] : 
                                (N173)? btb_q[1053] : 
                                (N175)? btb_q[1118] : 
                                (N177)? btb_q[1183] : 
                                (N179)? btb_q[1248] : 
                                (N181)? btb_q[1313] : 
                                (N183)? btb_q[1378] : 
                                (N185)? btb_q[1443] : 
                                (N187)? btb_q[1508] : 
                                (N189)? btb_q[1573] : 
                                (N191)? btb_q[1638] : 
                                (N193)? btb_q[1703] : 
                                (N195)? btb_q[1768] : 
                                (N197)? btb_q[1833] : 
                                (N199)? btb_q[1898] : 
                                (N201)? btb_q[1963] : 
                                (N203)? btb_q[2028] : 
                                (N142)? btb_q[2093] : 
                                (N144)? btb_q[2158] : 
                                (N146)? btb_q[2223] : 
                                (N148)? btb_q[2288] : 
                                (N150)? btb_q[2353] : 
                                (N152)? btb_q[2418] : 
                                (N154)? btb_q[2483] : 
                                (N156)? btb_q[2548] : 
                                (N158)? btb_q[2613] : 
                                (N160)? btb_q[2678] : 
                                (N162)? btb_q[2743] : 
                                (N164)? btb_q[2808] : 
                                (N166)? btb_q[2873] : 
                                (N168)? btb_q[2938] : 
                                (N170)? btb_q[3003] : 
                                (N172)? btb_q[3068] : 
                                (N174)? btb_q[3133] : 
                                (N176)? btb_q[3198] : 
                                (N178)? btb_q[3263] : 
                                (N180)? btb_q[3328] : 
                                (N182)? btb_q[3393] : 
                                (N184)? btb_q[3458] : 
                                (N186)? btb_q[3523] : 
                                (N188)? btb_q[3588] : 
                                (N190)? btb_q[3653] : 
                                (N192)? btb_q[3718] : 
                                (N194)? btb_q[3783] : 
                                (N196)? btb_q[3848] : 
                                (N198)? btb_q[3913] : 
                                (N200)? btb_q[3978] : 
                                (N202)? btb_q[4043] : 
                                (N204)? btb_q[4108] : 1'b0;
  assign btb_prediction_o[12] = (N141)? btb_q[12] : 
                                (N143)? btb_q[77] : 
                                (N145)? btb_q[142] : 
                                (N147)? btb_q[207] : 
                                (N149)? btb_q[272] : 
                                (N151)? btb_q[337] : 
                                (N153)? btb_q[402] : 
                                (N155)? btb_q[467] : 
                                (N157)? btb_q[532] : 
                                (N159)? btb_q[597] : 
                                (N161)? btb_q[662] : 
                                (N163)? btb_q[727] : 
                                (N165)? btb_q[792] : 
                                (N167)? btb_q[857] : 
                                (N169)? btb_q[922] : 
                                (N171)? btb_q[987] : 
                                (N173)? btb_q[1052] : 
                                (N175)? btb_q[1117] : 
                                (N177)? btb_q[1182] : 
                                (N179)? btb_q[1247] : 
                                (N181)? btb_q[1312] : 
                                (N183)? btb_q[1377] : 
                                (N185)? btb_q[1442] : 
                                (N187)? btb_q[1507] : 
                                (N189)? btb_q[1572] : 
                                (N191)? btb_q[1637] : 
                                (N193)? btb_q[1702] : 
                                (N195)? btb_q[1767] : 
                                (N197)? btb_q[1832] : 
                                (N199)? btb_q[1897] : 
                                (N201)? btb_q[1962] : 
                                (N203)? btb_q[2027] : 
                                (N142)? btb_q[2092] : 
                                (N144)? btb_q[2157] : 
                                (N146)? btb_q[2222] : 
                                (N148)? btb_q[2287] : 
                                (N150)? btb_q[2352] : 
                                (N152)? btb_q[2417] : 
                                (N154)? btb_q[2482] : 
                                (N156)? btb_q[2547] : 
                                (N158)? btb_q[2612] : 
                                (N160)? btb_q[2677] : 
                                (N162)? btb_q[2742] : 
                                (N164)? btb_q[2807] : 
                                (N166)? btb_q[2872] : 
                                (N168)? btb_q[2937] : 
                                (N170)? btb_q[3002] : 
                                (N172)? btb_q[3067] : 
                                (N174)? btb_q[3132] : 
                                (N176)? btb_q[3197] : 
                                (N178)? btb_q[3262] : 
                                (N180)? btb_q[3327] : 
                                (N182)? btb_q[3392] : 
                                (N184)? btb_q[3457] : 
                                (N186)? btb_q[3522] : 
                                (N188)? btb_q[3587] : 
                                (N190)? btb_q[3652] : 
                                (N192)? btb_q[3717] : 
                                (N194)? btb_q[3782] : 
                                (N196)? btb_q[3847] : 
                                (N198)? btb_q[3912] : 
                                (N200)? btb_q[3977] : 
                                (N202)? btb_q[4042] : 
                                (N204)? btb_q[4107] : 1'b0;
  assign btb_prediction_o[11] = (N141)? btb_q[11] : 
                                (N143)? btb_q[76] : 
                                (N145)? btb_q[141] : 
                                (N147)? btb_q[206] : 
                                (N149)? btb_q[271] : 
                                (N151)? btb_q[336] : 
                                (N153)? btb_q[401] : 
                                (N155)? btb_q[466] : 
                                (N157)? btb_q[531] : 
                                (N159)? btb_q[596] : 
                                (N161)? btb_q[661] : 
                                (N163)? btb_q[726] : 
                                (N165)? btb_q[791] : 
                                (N167)? btb_q[856] : 
                                (N169)? btb_q[921] : 
                                (N171)? btb_q[986] : 
                                (N173)? btb_q[1051] : 
                                (N175)? btb_q[1116] : 
                                (N177)? btb_q[1181] : 
                                (N179)? btb_q[1246] : 
                                (N181)? btb_q[1311] : 
                                (N183)? btb_q[1376] : 
                                (N185)? btb_q[1441] : 
                                (N187)? btb_q[1506] : 
                                (N189)? btb_q[1571] : 
                                (N191)? btb_q[1636] : 
                                (N193)? btb_q[1701] : 
                                (N195)? btb_q[1766] : 
                                (N197)? btb_q[1831] : 
                                (N199)? btb_q[1896] : 
                                (N201)? btb_q[1961] : 
                                (N203)? btb_q[2026] : 
                                (N142)? btb_q[2091] : 
                                (N144)? btb_q[2156] : 
                                (N146)? btb_q[2221] : 
                                (N148)? btb_q[2286] : 
                                (N150)? btb_q[2351] : 
                                (N152)? btb_q[2416] : 
                                (N154)? btb_q[2481] : 
                                (N156)? btb_q[2546] : 
                                (N158)? btb_q[2611] : 
                                (N160)? btb_q[2676] : 
                                (N162)? btb_q[2741] : 
                                (N164)? btb_q[2806] : 
                                (N166)? btb_q[2871] : 
                                (N168)? btb_q[2936] : 
                                (N170)? btb_q[3001] : 
                                (N172)? btb_q[3066] : 
                                (N174)? btb_q[3131] : 
                                (N176)? btb_q[3196] : 
                                (N178)? btb_q[3261] : 
                                (N180)? btb_q[3326] : 
                                (N182)? btb_q[3391] : 
                                (N184)? btb_q[3456] : 
                                (N186)? btb_q[3521] : 
                                (N188)? btb_q[3586] : 
                                (N190)? btb_q[3651] : 
                                (N192)? btb_q[3716] : 
                                (N194)? btb_q[3781] : 
                                (N196)? btb_q[3846] : 
                                (N198)? btb_q[3911] : 
                                (N200)? btb_q[3976] : 
                                (N202)? btb_q[4041] : 
                                (N204)? btb_q[4106] : 1'b0;
  assign btb_prediction_o[10] = (N141)? btb_q[10] : 
                                (N143)? btb_q[75] : 
                                (N145)? btb_q[140] : 
                                (N147)? btb_q[205] : 
                                (N149)? btb_q[270] : 
                                (N151)? btb_q[335] : 
                                (N153)? btb_q[400] : 
                                (N155)? btb_q[465] : 
                                (N157)? btb_q[530] : 
                                (N159)? btb_q[595] : 
                                (N161)? btb_q[660] : 
                                (N163)? btb_q[725] : 
                                (N165)? btb_q[790] : 
                                (N167)? btb_q[855] : 
                                (N169)? btb_q[920] : 
                                (N171)? btb_q[985] : 
                                (N173)? btb_q[1050] : 
                                (N175)? btb_q[1115] : 
                                (N177)? btb_q[1180] : 
                                (N179)? btb_q[1245] : 
                                (N181)? btb_q[1310] : 
                                (N183)? btb_q[1375] : 
                                (N185)? btb_q[1440] : 
                                (N187)? btb_q[1505] : 
                                (N189)? btb_q[1570] : 
                                (N191)? btb_q[1635] : 
                                (N193)? btb_q[1700] : 
                                (N195)? btb_q[1765] : 
                                (N197)? btb_q[1830] : 
                                (N199)? btb_q[1895] : 
                                (N201)? btb_q[1960] : 
                                (N203)? btb_q[2025] : 
                                (N142)? btb_q[2090] : 
                                (N144)? btb_q[2155] : 
                                (N146)? btb_q[2220] : 
                                (N148)? btb_q[2285] : 
                                (N150)? btb_q[2350] : 
                                (N152)? btb_q[2415] : 
                                (N154)? btb_q[2480] : 
                                (N156)? btb_q[2545] : 
                                (N158)? btb_q[2610] : 
                                (N160)? btb_q[2675] : 
                                (N162)? btb_q[2740] : 
                                (N164)? btb_q[2805] : 
                                (N166)? btb_q[2870] : 
                                (N168)? btb_q[2935] : 
                                (N170)? btb_q[3000] : 
                                (N172)? btb_q[3065] : 
                                (N174)? btb_q[3130] : 
                                (N176)? btb_q[3195] : 
                                (N178)? btb_q[3260] : 
                                (N180)? btb_q[3325] : 
                                (N182)? btb_q[3390] : 
                                (N184)? btb_q[3455] : 
                                (N186)? btb_q[3520] : 
                                (N188)? btb_q[3585] : 
                                (N190)? btb_q[3650] : 
                                (N192)? btb_q[3715] : 
                                (N194)? btb_q[3780] : 
                                (N196)? btb_q[3845] : 
                                (N198)? btb_q[3910] : 
                                (N200)? btb_q[3975] : 
                                (N202)? btb_q[4040] : 
                                (N204)? btb_q[4105] : 1'b0;
  assign btb_prediction_o[9] = (N141)? btb_q[9] : 
                               (N143)? btb_q[74] : 
                               (N145)? btb_q[139] : 
                               (N147)? btb_q[204] : 
                               (N149)? btb_q[269] : 
                               (N151)? btb_q[334] : 
                               (N153)? btb_q[399] : 
                               (N155)? btb_q[464] : 
                               (N157)? btb_q[529] : 
                               (N159)? btb_q[594] : 
                               (N161)? btb_q[659] : 
                               (N163)? btb_q[724] : 
                               (N165)? btb_q[789] : 
                               (N167)? btb_q[854] : 
                               (N169)? btb_q[919] : 
                               (N171)? btb_q[984] : 
                               (N173)? btb_q[1049] : 
                               (N175)? btb_q[1114] : 
                               (N177)? btb_q[1179] : 
                               (N179)? btb_q[1244] : 
                               (N181)? btb_q[1309] : 
                               (N183)? btb_q[1374] : 
                               (N185)? btb_q[1439] : 
                               (N187)? btb_q[1504] : 
                               (N189)? btb_q[1569] : 
                               (N191)? btb_q[1634] : 
                               (N193)? btb_q[1699] : 
                               (N195)? btb_q[1764] : 
                               (N197)? btb_q[1829] : 
                               (N199)? btb_q[1894] : 
                               (N201)? btb_q[1959] : 
                               (N203)? btb_q[2024] : 
                               (N142)? btb_q[2089] : 
                               (N144)? btb_q[2154] : 
                               (N146)? btb_q[2219] : 
                               (N148)? btb_q[2284] : 
                               (N150)? btb_q[2349] : 
                               (N152)? btb_q[2414] : 
                               (N154)? btb_q[2479] : 
                               (N156)? btb_q[2544] : 
                               (N158)? btb_q[2609] : 
                               (N160)? btb_q[2674] : 
                               (N162)? btb_q[2739] : 
                               (N164)? btb_q[2804] : 
                               (N166)? btb_q[2869] : 
                               (N168)? btb_q[2934] : 
                               (N170)? btb_q[2999] : 
                               (N172)? btb_q[3064] : 
                               (N174)? btb_q[3129] : 
                               (N176)? btb_q[3194] : 
                               (N178)? btb_q[3259] : 
                               (N180)? btb_q[3324] : 
                               (N182)? btb_q[3389] : 
                               (N184)? btb_q[3454] : 
                               (N186)? btb_q[3519] : 
                               (N188)? btb_q[3584] : 
                               (N190)? btb_q[3649] : 
                               (N192)? btb_q[3714] : 
                               (N194)? btb_q[3779] : 
                               (N196)? btb_q[3844] : 
                               (N198)? btb_q[3909] : 
                               (N200)? btb_q[3974] : 
                               (N202)? btb_q[4039] : 
                               (N204)? btb_q[4104] : 1'b0;
  assign btb_prediction_o[8] = (N141)? btb_q[8] : 
                               (N143)? btb_q[73] : 
                               (N145)? btb_q[138] : 
                               (N147)? btb_q[203] : 
                               (N149)? btb_q[268] : 
                               (N151)? btb_q[333] : 
                               (N153)? btb_q[398] : 
                               (N155)? btb_q[463] : 
                               (N157)? btb_q[528] : 
                               (N159)? btb_q[593] : 
                               (N161)? btb_q[658] : 
                               (N163)? btb_q[723] : 
                               (N165)? btb_q[788] : 
                               (N167)? btb_q[853] : 
                               (N169)? btb_q[918] : 
                               (N171)? btb_q[983] : 
                               (N173)? btb_q[1048] : 
                               (N175)? btb_q[1113] : 
                               (N177)? btb_q[1178] : 
                               (N179)? btb_q[1243] : 
                               (N181)? btb_q[1308] : 
                               (N183)? btb_q[1373] : 
                               (N185)? btb_q[1438] : 
                               (N187)? btb_q[1503] : 
                               (N189)? btb_q[1568] : 
                               (N191)? btb_q[1633] : 
                               (N193)? btb_q[1698] : 
                               (N195)? btb_q[1763] : 
                               (N197)? btb_q[1828] : 
                               (N199)? btb_q[1893] : 
                               (N201)? btb_q[1958] : 
                               (N203)? btb_q[2023] : 
                               (N142)? btb_q[2088] : 
                               (N144)? btb_q[2153] : 
                               (N146)? btb_q[2218] : 
                               (N148)? btb_q[2283] : 
                               (N150)? btb_q[2348] : 
                               (N152)? btb_q[2413] : 
                               (N154)? btb_q[2478] : 
                               (N156)? btb_q[2543] : 
                               (N158)? btb_q[2608] : 
                               (N160)? btb_q[2673] : 
                               (N162)? btb_q[2738] : 
                               (N164)? btb_q[2803] : 
                               (N166)? btb_q[2868] : 
                               (N168)? btb_q[2933] : 
                               (N170)? btb_q[2998] : 
                               (N172)? btb_q[3063] : 
                               (N174)? btb_q[3128] : 
                               (N176)? btb_q[3193] : 
                               (N178)? btb_q[3258] : 
                               (N180)? btb_q[3323] : 
                               (N182)? btb_q[3388] : 
                               (N184)? btb_q[3453] : 
                               (N186)? btb_q[3518] : 
                               (N188)? btb_q[3583] : 
                               (N190)? btb_q[3648] : 
                               (N192)? btb_q[3713] : 
                               (N194)? btb_q[3778] : 
                               (N196)? btb_q[3843] : 
                               (N198)? btb_q[3908] : 
                               (N200)? btb_q[3973] : 
                               (N202)? btb_q[4038] : 
                               (N204)? btb_q[4103] : 1'b0;
  assign btb_prediction_o[7] = (N141)? btb_q[7] : 
                               (N143)? btb_q[72] : 
                               (N145)? btb_q[137] : 
                               (N147)? btb_q[202] : 
                               (N149)? btb_q[267] : 
                               (N151)? btb_q[332] : 
                               (N153)? btb_q[397] : 
                               (N155)? btb_q[462] : 
                               (N157)? btb_q[527] : 
                               (N159)? btb_q[592] : 
                               (N161)? btb_q[657] : 
                               (N163)? btb_q[722] : 
                               (N165)? btb_q[787] : 
                               (N167)? btb_q[852] : 
                               (N169)? btb_q[917] : 
                               (N171)? btb_q[982] : 
                               (N173)? btb_q[1047] : 
                               (N175)? btb_q[1112] : 
                               (N177)? btb_q[1177] : 
                               (N179)? btb_q[1242] : 
                               (N181)? btb_q[1307] : 
                               (N183)? btb_q[1372] : 
                               (N185)? btb_q[1437] : 
                               (N187)? btb_q[1502] : 
                               (N189)? btb_q[1567] : 
                               (N191)? btb_q[1632] : 
                               (N193)? btb_q[1697] : 
                               (N195)? btb_q[1762] : 
                               (N197)? btb_q[1827] : 
                               (N199)? btb_q[1892] : 
                               (N201)? btb_q[1957] : 
                               (N203)? btb_q[2022] : 
                               (N142)? btb_q[2087] : 
                               (N144)? btb_q[2152] : 
                               (N146)? btb_q[2217] : 
                               (N148)? btb_q[2282] : 
                               (N150)? btb_q[2347] : 
                               (N152)? btb_q[2412] : 
                               (N154)? btb_q[2477] : 
                               (N156)? btb_q[2542] : 
                               (N158)? btb_q[2607] : 
                               (N160)? btb_q[2672] : 
                               (N162)? btb_q[2737] : 
                               (N164)? btb_q[2802] : 
                               (N166)? btb_q[2867] : 
                               (N168)? btb_q[2932] : 
                               (N170)? btb_q[2997] : 
                               (N172)? btb_q[3062] : 
                               (N174)? btb_q[3127] : 
                               (N176)? btb_q[3192] : 
                               (N178)? btb_q[3257] : 
                               (N180)? btb_q[3322] : 
                               (N182)? btb_q[3387] : 
                               (N184)? btb_q[3452] : 
                               (N186)? btb_q[3517] : 
                               (N188)? btb_q[3582] : 
                               (N190)? btb_q[3647] : 
                               (N192)? btb_q[3712] : 
                               (N194)? btb_q[3777] : 
                               (N196)? btb_q[3842] : 
                               (N198)? btb_q[3907] : 
                               (N200)? btb_q[3972] : 
                               (N202)? btb_q[4037] : 
                               (N204)? btb_q[4102] : 1'b0;
  assign btb_prediction_o[6] = (N141)? btb_q[6] : 
                               (N143)? btb_q[71] : 
                               (N145)? btb_q[136] : 
                               (N147)? btb_q[201] : 
                               (N149)? btb_q[266] : 
                               (N151)? btb_q[331] : 
                               (N153)? btb_q[396] : 
                               (N155)? btb_q[461] : 
                               (N157)? btb_q[526] : 
                               (N159)? btb_q[591] : 
                               (N161)? btb_q[656] : 
                               (N163)? btb_q[721] : 
                               (N165)? btb_q[786] : 
                               (N167)? btb_q[851] : 
                               (N169)? btb_q[916] : 
                               (N171)? btb_q[981] : 
                               (N173)? btb_q[1046] : 
                               (N175)? btb_q[1111] : 
                               (N177)? btb_q[1176] : 
                               (N179)? btb_q[1241] : 
                               (N181)? btb_q[1306] : 
                               (N183)? btb_q[1371] : 
                               (N185)? btb_q[1436] : 
                               (N187)? btb_q[1501] : 
                               (N189)? btb_q[1566] : 
                               (N191)? btb_q[1631] : 
                               (N193)? btb_q[1696] : 
                               (N195)? btb_q[1761] : 
                               (N197)? btb_q[1826] : 
                               (N199)? btb_q[1891] : 
                               (N201)? btb_q[1956] : 
                               (N203)? btb_q[2021] : 
                               (N142)? btb_q[2086] : 
                               (N144)? btb_q[2151] : 
                               (N146)? btb_q[2216] : 
                               (N148)? btb_q[2281] : 
                               (N150)? btb_q[2346] : 
                               (N152)? btb_q[2411] : 
                               (N154)? btb_q[2476] : 
                               (N156)? btb_q[2541] : 
                               (N158)? btb_q[2606] : 
                               (N160)? btb_q[2671] : 
                               (N162)? btb_q[2736] : 
                               (N164)? btb_q[2801] : 
                               (N166)? btb_q[2866] : 
                               (N168)? btb_q[2931] : 
                               (N170)? btb_q[2996] : 
                               (N172)? btb_q[3061] : 
                               (N174)? btb_q[3126] : 
                               (N176)? btb_q[3191] : 
                               (N178)? btb_q[3256] : 
                               (N180)? btb_q[3321] : 
                               (N182)? btb_q[3386] : 
                               (N184)? btb_q[3451] : 
                               (N186)? btb_q[3516] : 
                               (N188)? btb_q[3581] : 
                               (N190)? btb_q[3646] : 
                               (N192)? btb_q[3711] : 
                               (N194)? btb_q[3776] : 
                               (N196)? btb_q[3841] : 
                               (N198)? btb_q[3906] : 
                               (N200)? btb_q[3971] : 
                               (N202)? btb_q[4036] : 
                               (N204)? btb_q[4101] : 1'b0;
  assign btb_prediction_o[5] = (N141)? btb_q[5] : 
                               (N143)? btb_q[70] : 
                               (N145)? btb_q[135] : 
                               (N147)? btb_q[200] : 
                               (N149)? btb_q[265] : 
                               (N151)? btb_q[330] : 
                               (N153)? btb_q[395] : 
                               (N155)? btb_q[460] : 
                               (N157)? btb_q[525] : 
                               (N159)? btb_q[590] : 
                               (N161)? btb_q[655] : 
                               (N163)? btb_q[720] : 
                               (N165)? btb_q[785] : 
                               (N167)? btb_q[850] : 
                               (N169)? btb_q[915] : 
                               (N171)? btb_q[980] : 
                               (N173)? btb_q[1045] : 
                               (N175)? btb_q[1110] : 
                               (N177)? btb_q[1175] : 
                               (N179)? btb_q[1240] : 
                               (N181)? btb_q[1305] : 
                               (N183)? btb_q[1370] : 
                               (N185)? btb_q[1435] : 
                               (N187)? btb_q[1500] : 
                               (N189)? btb_q[1565] : 
                               (N191)? btb_q[1630] : 
                               (N193)? btb_q[1695] : 
                               (N195)? btb_q[1760] : 
                               (N197)? btb_q[1825] : 
                               (N199)? btb_q[1890] : 
                               (N201)? btb_q[1955] : 
                               (N203)? btb_q[2020] : 
                               (N142)? btb_q[2085] : 
                               (N144)? btb_q[2150] : 
                               (N146)? btb_q[2215] : 
                               (N148)? btb_q[2280] : 
                               (N150)? btb_q[2345] : 
                               (N152)? btb_q[2410] : 
                               (N154)? btb_q[2475] : 
                               (N156)? btb_q[2540] : 
                               (N158)? btb_q[2605] : 
                               (N160)? btb_q[2670] : 
                               (N162)? btb_q[2735] : 
                               (N164)? btb_q[2800] : 
                               (N166)? btb_q[2865] : 
                               (N168)? btb_q[2930] : 
                               (N170)? btb_q[2995] : 
                               (N172)? btb_q[3060] : 
                               (N174)? btb_q[3125] : 
                               (N176)? btb_q[3190] : 
                               (N178)? btb_q[3255] : 
                               (N180)? btb_q[3320] : 
                               (N182)? btb_q[3385] : 
                               (N184)? btb_q[3450] : 
                               (N186)? btb_q[3515] : 
                               (N188)? btb_q[3580] : 
                               (N190)? btb_q[3645] : 
                               (N192)? btb_q[3710] : 
                               (N194)? btb_q[3775] : 
                               (N196)? btb_q[3840] : 
                               (N198)? btb_q[3905] : 
                               (N200)? btb_q[3970] : 
                               (N202)? btb_q[4035] : 
                               (N204)? btb_q[4100] : 1'b0;
  assign btb_prediction_o[4] = (N141)? btb_q[4] : 
                               (N143)? btb_q[69] : 
                               (N145)? btb_q[134] : 
                               (N147)? btb_q[199] : 
                               (N149)? btb_q[264] : 
                               (N151)? btb_q[329] : 
                               (N153)? btb_q[394] : 
                               (N155)? btb_q[459] : 
                               (N157)? btb_q[524] : 
                               (N159)? btb_q[589] : 
                               (N161)? btb_q[654] : 
                               (N163)? btb_q[719] : 
                               (N165)? btb_q[784] : 
                               (N167)? btb_q[849] : 
                               (N169)? btb_q[914] : 
                               (N171)? btb_q[979] : 
                               (N173)? btb_q[1044] : 
                               (N175)? btb_q[1109] : 
                               (N177)? btb_q[1174] : 
                               (N179)? btb_q[1239] : 
                               (N181)? btb_q[1304] : 
                               (N183)? btb_q[1369] : 
                               (N185)? btb_q[1434] : 
                               (N187)? btb_q[1499] : 
                               (N189)? btb_q[1564] : 
                               (N191)? btb_q[1629] : 
                               (N193)? btb_q[1694] : 
                               (N195)? btb_q[1759] : 
                               (N197)? btb_q[1824] : 
                               (N199)? btb_q[1889] : 
                               (N201)? btb_q[1954] : 
                               (N203)? btb_q[2019] : 
                               (N142)? btb_q[2084] : 
                               (N144)? btb_q[2149] : 
                               (N146)? btb_q[2214] : 
                               (N148)? btb_q[2279] : 
                               (N150)? btb_q[2344] : 
                               (N152)? btb_q[2409] : 
                               (N154)? btb_q[2474] : 
                               (N156)? btb_q[2539] : 
                               (N158)? btb_q[2604] : 
                               (N160)? btb_q[2669] : 
                               (N162)? btb_q[2734] : 
                               (N164)? btb_q[2799] : 
                               (N166)? btb_q[2864] : 
                               (N168)? btb_q[2929] : 
                               (N170)? btb_q[2994] : 
                               (N172)? btb_q[3059] : 
                               (N174)? btb_q[3124] : 
                               (N176)? btb_q[3189] : 
                               (N178)? btb_q[3254] : 
                               (N180)? btb_q[3319] : 
                               (N182)? btb_q[3384] : 
                               (N184)? btb_q[3449] : 
                               (N186)? btb_q[3514] : 
                               (N188)? btb_q[3579] : 
                               (N190)? btb_q[3644] : 
                               (N192)? btb_q[3709] : 
                               (N194)? btb_q[3774] : 
                               (N196)? btb_q[3839] : 
                               (N198)? btb_q[3904] : 
                               (N200)? btb_q[3969] : 
                               (N202)? btb_q[4034] : 
                               (N204)? btb_q[4099] : 1'b0;
  assign btb_prediction_o[3] = (N141)? btb_q[3] : 
                               (N143)? btb_q[68] : 
                               (N145)? btb_q[133] : 
                               (N147)? btb_q[198] : 
                               (N149)? btb_q[263] : 
                               (N151)? btb_q[328] : 
                               (N153)? btb_q[393] : 
                               (N155)? btb_q[458] : 
                               (N157)? btb_q[523] : 
                               (N159)? btb_q[588] : 
                               (N161)? btb_q[653] : 
                               (N163)? btb_q[718] : 
                               (N165)? btb_q[783] : 
                               (N167)? btb_q[848] : 
                               (N169)? btb_q[913] : 
                               (N171)? btb_q[978] : 
                               (N173)? btb_q[1043] : 
                               (N175)? btb_q[1108] : 
                               (N177)? btb_q[1173] : 
                               (N179)? btb_q[1238] : 
                               (N181)? btb_q[1303] : 
                               (N183)? btb_q[1368] : 
                               (N185)? btb_q[1433] : 
                               (N187)? btb_q[1498] : 
                               (N189)? btb_q[1563] : 
                               (N191)? btb_q[1628] : 
                               (N193)? btb_q[1693] : 
                               (N195)? btb_q[1758] : 
                               (N197)? btb_q[1823] : 
                               (N199)? btb_q[1888] : 
                               (N201)? btb_q[1953] : 
                               (N203)? btb_q[2018] : 
                               (N142)? btb_q[2083] : 
                               (N144)? btb_q[2148] : 
                               (N146)? btb_q[2213] : 
                               (N148)? btb_q[2278] : 
                               (N150)? btb_q[2343] : 
                               (N152)? btb_q[2408] : 
                               (N154)? btb_q[2473] : 
                               (N156)? btb_q[2538] : 
                               (N158)? btb_q[2603] : 
                               (N160)? btb_q[2668] : 
                               (N162)? btb_q[2733] : 
                               (N164)? btb_q[2798] : 
                               (N166)? btb_q[2863] : 
                               (N168)? btb_q[2928] : 
                               (N170)? btb_q[2993] : 
                               (N172)? btb_q[3058] : 
                               (N174)? btb_q[3123] : 
                               (N176)? btb_q[3188] : 
                               (N178)? btb_q[3253] : 
                               (N180)? btb_q[3318] : 
                               (N182)? btb_q[3383] : 
                               (N184)? btb_q[3448] : 
                               (N186)? btb_q[3513] : 
                               (N188)? btb_q[3578] : 
                               (N190)? btb_q[3643] : 
                               (N192)? btb_q[3708] : 
                               (N194)? btb_q[3773] : 
                               (N196)? btb_q[3838] : 
                               (N198)? btb_q[3903] : 
                               (N200)? btb_q[3968] : 
                               (N202)? btb_q[4033] : 
                               (N204)? btb_q[4098] : 1'b0;
  assign btb_prediction_o[2] = (N141)? btb_q[2] : 
                               (N143)? btb_q[67] : 
                               (N145)? btb_q[132] : 
                               (N147)? btb_q[197] : 
                               (N149)? btb_q[262] : 
                               (N151)? btb_q[327] : 
                               (N153)? btb_q[392] : 
                               (N155)? btb_q[457] : 
                               (N157)? btb_q[522] : 
                               (N159)? btb_q[587] : 
                               (N161)? btb_q[652] : 
                               (N163)? btb_q[717] : 
                               (N165)? btb_q[782] : 
                               (N167)? btb_q[847] : 
                               (N169)? btb_q[912] : 
                               (N171)? btb_q[977] : 
                               (N173)? btb_q[1042] : 
                               (N175)? btb_q[1107] : 
                               (N177)? btb_q[1172] : 
                               (N179)? btb_q[1237] : 
                               (N181)? btb_q[1302] : 
                               (N183)? btb_q[1367] : 
                               (N185)? btb_q[1432] : 
                               (N187)? btb_q[1497] : 
                               (N189)? btb_q[1562] : 
                               (N191)? btb_q[1627] : 
                               (N193)? btb_q[1692] : 
                               (N195)? btb_q[1757] : 
                               (N197)? btb_q[1822] : 
                               (N199)? btb_q[1887] : 
                               (N201)? btb_q[1952] : 
                               (N203)? btb_q[2017] : 
                               (N142)? btb_q[2082] : 
                               (N144)? btb_q[2147] : 
                               (N146)? btb_q[2212] : 
                               (N148)? btb_q[2277] : 
                               (N150)? btb_q[2342] : 
                               (N152)? btb_q[2407] : 
                               (N154)? btb_q[2472] : 
                               (N156)? btb_q[2537] : 
                               (N158)? btb_q[2602] : 
                               (N160)? btb_q[2667] : 
                               (N162)? btb_q[2732] : 
                               (N164)? btb_q[2797] : 
                               (N166)? btb_q[2862] : 
                               (N168)? btb_q[2927] : 
                               (N170)? btb_q[2992] : 
                               (N172)? btb_q[3057] : 
                               (N174)? btb_q[3122] : 
                               (N176)? btb_q[3187] : 
                               (N178)? btb_q[3252] : 
                               (N180)? btb_q[3317] : 
                               (N182)? btb_q[3382] : 
                               (N184)? btb_q[3447] : 
                               (N186)? btb_q[3512] : 
                               (N188)? btb_q[3577] : 
                               (N190)? btb_q[3642] : 
                               (N192)? btb_q[3707] : 
                               (N194)? btb_q[3772] : 
                               (N196)? btb_q[3837] : 
                               (N198)? btb_q[3902] : 
                               (N200)? btb_q[3967] : 
                               (N202)? btb_q[4032] : 
                               (N204)? btb_q[4097] : 1'b0;
  assign btb_prediction_o[1] = (N141)? btb_q[1] : 
                               (N143)? btb_q[66] : 
                               (N145)? btb_q[131] : 
                               (N147)? btb_q[196] : 
                               (N149)? btb_q[261] : 
                               (N151)? btb_q[326] : 
                               (N153)? btb_q[391] : 
                               (N155)? btb_q[456] : 
                               (N157)? btb_q[521] : 
                               (N159)? btb_q[586] : 
                               (N161)? btb_q[651] : 
                               (N163)? btb_q[716] : 
                               (N165)? btb_q[781] : 
                               (N167)? btb_q[846] : 
                               (N169)? btb_q[911] : 
                               (N171)? btb_q[976] : 
                               (N173)? btb_q[1041] : 
                               (N175)? btb_q[1106] : 
                               (N177)? btb_q[1171] : 
                               (N179)? btb_q[1236] : 
                               (N181)? btb_q[1301] : 
                               (N183)? btb_q[1366] : 
                               (N185)? btb_q[1431] : 
                               (N187)? btb_q[1496] : 
                               (N189)? btb_q[1561] : 
                               (N191)? btb_q[1626] : 
                               (N193)? btb_q[1691] : 
                               (N195)? btb_q[1756] : 
                               (N197)? btb_q[1821] : 
                               (N199)? btb_q[1886] : 
                               (N201)? btb_q[1951] : 
                               (N203)? btb_q[2016] : 
                               (N142)? btb_q[2081] : 
                               (N144)? btb_q[2146] : 
                               (N146)? btb_q[2211] : 
                               (N148)? btb_q[2276] : 
                               (N150)? btb_q[2341] : 
                               (N152)? btb_q[2406] : 
                               (N154)? btb_q[2471] : 
                               (N156)? btb_q[2536] : 
                               (N158)? btb_q[2601] : 
                               (N160)? btb_q[2666] : 
                               (N162)? btb_q[2731] : 
                               (N164)? btb_q[2796] : 
                               (N166)? btb_q[2861] : 
                               (N168)? btb_q[2926] : 
                               (N170)? btb_q[2991] : 
                               (N172)? btb_q[3056] : 
                               (N174)? btb_q[3121] : 
                               (N176)? btb_q[3186] : 
                               (N178)? btb_q[3251] : 
                               (N180)? btb_q[3316] : 
                               (N182)? btb_q[3381] : 
                               (N184)? btb_q[3446] : 
                               (N186)? btb_q[3511] : 
                               (N188)? btb_q[3576] : 
                               (N190)? btb_q[3641] : 
                               (N192)? btb_q[3706] : 
                               (N194)? btb_q[3771] : 
                               (N196)? btb_q[3836] : 
                               (N198)? btb_q[3901] : 
                               (N200)? btb_q[3966] : 
                               (N202)? btb_q[4031] : 
                               (N204)? btb_q[4096] : 1'b0;
  assign btb_prediction_o[0] = (N141)? btb_q[0] : 
                               (N143)? btb_q[65] : 
                               (N145)? btb_q[130] : 
                               (N147)? btb_q[195] : 
                               (N149)? btb_q[260] : 
                               (N151)? btb_q[325] : 
                               (N153)? btb_q[390] : 
                               (N155)? btb_q[455] : 
                               (N157)? btb_q[520] : 
                               (N159)? btb_q[585] : 
                               (N161)? btb_q[650] : 
                               (N163)? btb_q[715] : 
                               (N165)? btb_q[780] : 
                               (N167)? btb_q[845] : 
                               (N169)? btb_q[910] : 
                               (N171)? btb_q[975] : 
                               (N173)? btb_q[1040] : 
                               (N175)? btb_q[1105] : 
                               (N177)? btb_q[1170] : 
                               (N179)? btb_q[1235] : 
                               (N181)? btb_q[1300] : 
                               (N183)? btb_q[1365] : 
                               (N185)? btb_q[1430] : 
                               (N187)? btb_q[1495] : 
                               (N189)? btb_q[1560] : 
                               (N191)? btb_q[1625] : 
                               (N193)? btb_q[1690] : 
                               (N195)? btb_q[1755] : 
                               (N197)? btb_q[1820] : 
                               (N199)? btb_q[1885] : 
                               (N201)? btb_q[1950] : 
                               (N203)? btb_q[2015] : 
                               (N142)? btb_q[2080] : 
                               (N144)? btb_q[2145] : 
                               (N146)? btb_q[2210] : 
                               (N148)? btb_q[2275] : 
                               (N150)? btb_q[2340] : 
                               (N152)? btb_q[2405] : 
                               (N154)? btb_q[2470] : 
                               (N156)? btb_q[2535] : 
                               (N158)? btb_q[2600] : 
                               (N160)? btb_q[2665] : 
                               (N162)? btb_q[2730] : 
                               (N164)? btb_q[2795] : 
                               (N166)? btb_q[2860] : 
                               (N168)? btb_q[2925] : 
                               (N170)? btb_q[2990] : 
                               (N172)? btb_q[3055] : 
                               (N174)? btb_q[3120] : 
                               (N176)? btb_q[3185] : 
                               (N178)? btb_q[3250] : 
                               (N180)? btb_q[3315] : 
                               (N182)? btb_q[3380] : 
                               (N184)? btb_q[3445] : 
                               (N186)? btb_q[3510] : 
                               (N188)? btb_q[3575] : 
                               (N190)? btb_q[3640] : 
                               (N192)? btb_q[3705] : 
                               (N194)? btb_q[3770] : 
                               (N196)? btb_q[3835] : 
                               (N198)? btb_q[3900] : 
                               (N200)? btb_q[3965] : 
                               (N202)? btb_q[4030] : 
                               (N204)? btb_q[4095] : 1'b0;

  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4159] <= 1'b0;
    end else if(N595) begin
      btb_q[4159] <= N593;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4158] <= 1'b0;
    end else if(N601) begin
      btb_q[4158] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4157] <= 1'b0;
    end else if(N607) begin
      btb_q[4157] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4156] <= 1'b0;
    end else if(N613) begin
      btb_q[4156] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4155] <= 1'b0;
    end else if(N619) begin
      btb_q[4155] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4154] <= 1'b0;
    end else if(N625) begin
      btb_q[4154] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4153] <= 1'b0;
    end else if(N631) begin
      btb_q[4153] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4152] <= 1'b0;
    end else if(N637) begin
      btb_q[4152] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4151] <= 1'b0;
    end else if(N643) begin
      btb_q[4151] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4150] <= 1'b0;
    end else if(N649) begin
      btb_q[4150] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4149] <= 1'b0;
    end else if(N655) begin
      btb_q[4149] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4148] <= 1'b0;
    end else if(N661) begin
      btb_q[4148] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4147] <= 1'b0;
    end else if(N667) begin
      btb_q[4147] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4146] <= 1'b0;
    end else if(N673) begin
      btb_q[4146] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4145] <= 1'b0;
    end else if(N679) begin
      btb_q[4145] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4144] <= 1'b0;
    end else if(N685) begin
      btb_q[4144] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4143] <= 1'b0;
    end else if(N691) begin
      btb_q[4143] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4142] <= 1'b0;
    end else if(N697) begin
      btb_q[4142] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4141] <= 1'b0;
    end else if(N703) begin
      btb_q[4141] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4140] <= 1'b0;
    end else if(N709) begin
      btb_q[4140] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4139] <= 1'b0;
    end else if(N715) begin
      btb_q[4139] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4138] <= 1'b0;
    end else if(N721) begin
      btb_q[4138] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4137] <= 1'b0;
    end else if(N727) begin
      btb_q[4137] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4136] <= 1'b0;
    end else if(N733) begin
      btb_q[4136] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4135] <= 1'b0;
    end else if(N739) begin
      btb_q[4135] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4134] <= 1'b0;
    end else if(N745) begin
      btb_q[4134] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4133] <= 1'b0;
    end else if(N751) begin
      btb_q[4133] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4132] <= 1'b0;
    end else if(N757) begin
      btb_q[4132] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4131] <= 1'b0;
    end else if(N763) begin
      btb_q[4131] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4130] <= 1'b0;
    end else if(N769) begin
      btb_q[4130] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4129] <= 1'b0;
    end else if(N775) begin
      btb_q[4129] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4128] <= 1'b0;
    end else if(N781) begin
      btb_q[4128] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4127] <= 1'b0;
    end else if(N787) begin
      btb_q[4127] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4126] <= 1'b0;
    end else if(N793) begin
      btb_q[4126] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4125] <= 1'b0;
    end else if(N799) begin
      btb_q[4125] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4124] <= 1'b0;
    end else if(N805) begin
      btb_q[4124] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4123] <= 1'b0;
    end else if(N811) begin
      btb_q[4123] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4122] <= 1'b0;
    end else if(N817) begin
      btb_q[4122] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4121] <= 1'b0;
    end else if(N823) begin
      btb_q[4121] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4120] <= 1'b0;
    end else if(N829) begin
      btb_q[4120] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4119] <= 1'b0;
    end else if(N835) begin
      btb_q[4119] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4118] <= 1'b0;
    end else if(N841) begin
      btb_q[4118] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4117] <= 1'b0;
    end else if(N841) begin
      btb_q[4117] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4116] <= 1'b0;
    end else if(N841) begin
      btb_q[4116] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4115] <= 1'b0;
    end else if(N841) begin
      btb_q[4115] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4114] <= 1'b0;
    end else if(N841) begin
      btb_q[4114] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4113] <= 1'b0;
    end else if(N841) begin
      btb_q[4113] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4112] <= 1'b0;
    end else if(N841) begin
      btb_q[4112] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4111] <= 1'b0;
    end else if(N841) begin
      btb_q[4111] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4110] <= 1'b0;
    end else if(N841) begin
      btb_q[4110] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4109] <= 1'b0;
    end else if(N841) begin
      btb_q[4109] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4108] <= 1'b0;
    end else if(N841) begin
      btb_q[4108] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4107] <= 1'b0;
    end else if(N841) begin
      btb_q[4107] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4106] <= 1'b0;
    end else if(N841) begin
      btb_q[4106] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4105] <= 1'b0;
    end else if(N841) begin
      btb_q[4105] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4104] <= 1'b0;
    end else if(N841) begin
      btb_q[4104] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4103] <= 1'b0;
    end else if(N841) begin
      btb_q[4103] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4102] <= 1'b0;
    end else if(N841) begin
      btb_q[4102] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4101] <= 1'b0;
    end else if(N841) begin
      btb_q[4101] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4100] <= 1'b0;
    end else if(N841) begin
      btb_q[4100] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4099] <= 1'b0;
    end else if(N841) begin
      btb_q[4099] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4098] <= 1'b0;
    end else if(N841) begin
      btb_q[4098] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4097] <= 1'b0;
    end else if(N841) begin
      btb_q[4097] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4096] <= 1'b0;
    end else if(N841) begin
      btb_q[4096] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4095] <= 1'b0;
    end else if(N841) begin
      btb_q[4095] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4094] <= 1'b0;
    end else if(N842) begin
      btb_q[4094] <= N592;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4093] <= 1'b0;
    end else if(N846) begin
      btb_q[4093] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4092] <= 1'b0;
    end else if(N846) begin
      btb_q[4092] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4091] <= 1'b0;
    end else if(N846) begin
      btb_q[4091] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4090] <= 1'b0;
    end else if(N846) begin
      btb_q[4090] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4089] <= 1'b0;
    end else if(N846) begin
      btb_q[4089] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4088] <= 1'b0;
    end else if(N846) begin
      btb_q[4088] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4087] <= 1'b0;
    end else if(N846) begin
      btb_q[4087] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4086] <= 1'b0;
    end else if(N846) begin
      btb_q[4086] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4085] <= 1'b0;
    end else if(N846) begin
      btb_q[4085] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4084] <= 1'b0;
    end else if(N846) begin
      btb_q[4084] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4083] <= 1'b0;
    end else if(N846) begin
      btb_q[4083] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4082] <= 1'b0;
    end else if(N846) begin
      btb_q[4082] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4081] <= 1'b0;
    end else if(N846) begin
      btb_q[4081] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4080] <= 1'b0;
    end else if(N846) begin
      btb_q[4080] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4079] <= 1'b0;
    end else if(N846) begin
      btb_q[4079] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4078] <= 1'b0;
    end else if(N846) begin
      btb_q[4078] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4077] <= 1'b0;
    end else if(N846) begin
      btb_q[4077] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4076] <= 1'b0;
    end else if(N846) begin
      btb_q[4076] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4075] <= 1'b0;
    end else if(N846) begin
      btb_q[4075] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4074] <= 1'b0;
    end else if(N846) begin
      btb_q[4074] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4073] <= 1'b0;
    end else if(N846) begin
      btb_q[4073] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4072] <= 1'b0;
    end else if(N846) begin
      btb_q[4072] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4071] <= 1'b0;
    end else if(N846) begin
      btb_q[4071] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4070] <= 1'b0;
    end else if(N846) begin
      btb_q[4070] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4069] <= 1'b0;
    end else if(N846) begin
      btb_q[4069] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4068] <= 1'b0;
    end else if(N846) begin
      btb_q[4068] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4067] <= 1'b0;
    end else if(N846) begin
      btb_q[4067] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4066] <= 1'b0;
    end else if(N846) begin
      btb_q[4066] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4065] <= 1'b0;
    end else if(N846) begin
      btb_q[4065] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4064] <= 1'b0;
    end else if(N846) begin
      btb_q[4064] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4063] <= 1'b0;
    end else if(N846) begin
      btb_q[4063] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4062] <= 1'b0;
    end else if(N846) begin
      btb_q[4062] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4061] <= 1'b0;
    end else if(N846) begin
      btb_q[4061] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4060] <= 1'b0;
    end else if(N846) begin
      btb_q[4060] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4059] <= 1'b0;
    end else if(N846) begin
      btb_q[4059] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4058] <= 1'b0;
    end else if(N849) begin
      btb_q[4058] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4057] <= 1'b0;
    end else if(N849) begin
      btb_q[4057] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4056] <= 1'b0;
    end else if(N849) begin
      btb_q[4056] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4055] <= 1'b0;
    end else if(N849) begin
      btb_q[4055] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4054] <= 1'b0;
    end else if(N849) begin
      btb_q[4054] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4053] <= 1'b0;
    end else if(N849) begin
      btb_q[4053] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4052] <= 1'b0;
    end else if(N849) begin
      btb_q[4052] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4051] <= 1'b0;
    end else if(N849) begin
      btb_q[4051] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4050] <= 1'b0;
    end else if(N849) begin
      btb_q[4050] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4049] <= 1'b0;
    end else if(N849) begin
      btb_q[4049] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4048] <= 1'b0;
    end else if(N849) begin
      btb_q[4048] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4047] <= 1'b0;
    end else if(N849) begin
      btb_q[4047] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4046] <= 1'b0;
    end else if(N849) begin
      btb_q[4046] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4045] <= 1'b0;
    end else if(N849) begin
      btb_q[4045] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4044] <= 1'b0;
    end else if(N849) begin
      btb_q[4044] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4043] <= 1'b0;
    end else if(N849) begin
      btb_q[4043] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4042] <= 1'b0;
    end else if(N849) begin
      btb_q[4042] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4041] <= 1'b0;
    end else if(N849) begin
      btb_q[4041] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4040] <= 1'b0;
    end else if(N849) begin
      btb_q[4040] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4039] <= 1'b0;
    end else if(N849) begin
      btb_q[4039] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4038] <= 1'b0;
    end else if(N849) begin
      btb_q[4038] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4037] <= 1'b0;
    end else if(N849) begin
      btb_q[4037] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4036] <= 1'b0;
    end else if(N849) begin
      btb_q[4036] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4035] <= 1'b0;
    end else if(N849) begin
      btb_q[4035] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4034] <= 1'b0;
    end else if(N849) begin
      btb_q[4034] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4033] <= 1'b0;
    end else if(N849) begin
      btb_q[4033] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4032] <= 1'b0;
    end else if(N849) begin
      btb_q[4032] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4031] <= 1'b0;
    end else if(N849) begin
      btb_q[4031] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4030] <= 1'b0;
    end else if(N849) begin
      btb_q[4030] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4029] <= 1'b0;
    end else if(N850) begin
      btb_q[4029] <= N591;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4028] <= 1'b0;
    end else if(N854) begin
      btb_q[4028] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4027] <= 1'b0;
    end else if(N854) begin
      btb_q[4027] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4026] <= 1'b0;
    end else if(N854) begin
      btb_q[4026] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4025] <= 1'b0;
    end else if(N854) begin
      btb_q[4025] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4024] <= 1'b0;
    end else if(N854) begin
      btb_q[4024] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4023] <= 1'b0;
    end else if(N854) begin
      btb_q[4023] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4022] <= 1'b0;
    end else if(N854) begin
      btb_q[4022] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4021] <= 1'b0;
    end else if(N854) begin
      btb_q[4021] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4020] <= 1'b0;
    end else if(N858) begin
      btb_q[4020] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4019] <= 1'b0;
    end else if(N858) begin
      btb_q[4019] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4018] <= 1'b0;
    end else if(N858) begin
      btb_q[4018] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4017] <= 1'b0;
    end else if(N858) begin
      btb_q[4017] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4016] <= 1'b0;
    end else if(N858) begin
      btb_q[4016] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4015] <= 1'b0;
    end else if(N858) begin
      btb_q[4015] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4014] <= 1'b0;
    end else if(N858) begin
      btb_q[4014] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4013] <= 1'b0;
    end else if(N858) begin
      btb_q[4013] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4012] <= 1'b0;
    end else if(N858) begin
      btb_q[4012] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4011] <= 1'b0;
    end else if(N858) begin
      btb_q[4011] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4010] <= 1'b0;
    end else if(N858) begin
      btb_q[4010] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4009] <= 1'b0;
    end else if(N858) begin
      btb_q[4009] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4008] <= 1'b0;
    end else if(N858) begin
      btb_q[4008] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4007] <= 1'b0;
    end else if(N858) begin
      btb_q[4007] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4006] <= 1'b0;
    end else if(N858) begin
      btb_q[4006] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4005] <= 1'b0;
    end else if(N858) begin
      btb_q[4005] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4004] <= 1'b0;
    end else if(N858) begin
      btb_q[4004] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4003] <= 1'b0;
    end else if(N858) begin
      btb_q[4003] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4002] <= 1'b0;
    end else if(N858) begin
      btb_q[4002] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4001] <= 1'b0;
    end else if(N858) begin
      btb_q[4001] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4000] <= 1'b0;
    end else if(N858) begin
      btb_q[4000] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3999] <= 1'b0;
    end else if(N858) begin
      btb_q[3999] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3998] <= 1'b0;
    end else if(N858) begin
      btb_q[3998] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3997] <= 1'b0;
    end else if(N858) begin
      btb_q[3997] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3996] <= 1'b0;
    end else if(N858) begin
      btb_q[3996] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3995] <= 1'b0;
    end else if(N858) begin
      btb_q[3995] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3994] <= 1'b0;
    end else if(N858) begin
      btb_q[3994] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3993] <= 1'b0;
    end else if(N858) begin
      btb_q[3993] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3992] <= 1'b0;
    end else if(N858) begin
      btb_q[3992] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3991] <= 1'b0;
    end else if(N858) begin
      btb_q[3991] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3990] <= 1'b0;
    end else if(N858) begin
      btb_q[3990] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3989] <= 1'b0;
    end else if(N858) begin
      btb_q[3989] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3988] <= 1'b0;
    end else if(N858) begin
      btb_q[3988] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3987] <= 1'b0;
    end else if(N858) begin
      btb_q[3987] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3986] <= 1'b0;
    end else if(N858) begin
      btb_q[3986] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3985] <= 1'b0;
    end else if(N858) begin
      btb_q[3985] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3984] <= 1'b0;
    end else if(N858) begin
      btb_q[3984] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3983] <= 1'b0;
    end else if(N858) begin
      btb_q[3983] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3982] <= 1'b0;
    end else if(N858) begin
      btb_q[3982] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3981] <= 1'b0;
    end else if(N858) begin
      btb_q[3981] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3980] <= 1'b0;
    end else if(N858) begin
      btb_q[3980] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3979] <= 1'b0;
    end else if(N858) begin
      btb_q[3979] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3978] <= 1'b0;
    end else if(N858) begin
      btb_q[3978] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3977] <= 1'b0;
    end else if(N858) begin
      btb_q[3977] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3976] <= 1'b0;
    end else if(N858) begin
      btb_q[3976] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3975] <= 1'b0;
    end else if(N858) begin
      btb_q[3975] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3974] <= 1'b0;
    end else if(N858) begin
      btb_q[3974] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3973] <= 1'b0;
    end else if(N858) begin
      btb_q[3973] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3972] <= 1'b0;
    end else if(N858) begin
      btb_q[3972] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3971] <= 1'b0;
    end else if(N858) begin
      btb_q[3971] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3970] <= 1'b0;
    end else if(N858) begin
      btb_q[3970] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3969] <= 1'b0;
    end else if(N858) begin
      btb_q[3969] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3968] <= 1'b0;
    end else if(N858) begin
      btb_q[3968] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3967] <= 1'b0;
    end else if(N858) begin
      btb_q[3967] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3966] <= 1'b0;
    end else if(N858) begin
      btb_q[3966] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3965] <= 1'b0;
    end else if(N858) begin
      btb_q[3965] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3964] <= 1'b0;
    end else if(N850) begin
      btb_q[3964] <= N590;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3963] <= 1'b0;
    end else if(N862) begin
      btb_q[3963] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3962] <= 1'b0;
    end else if(N862) begin
      btb_q[3962] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3961] <= 1'b0;
    end else if(N862) begin
      btb_q[3961] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3960] <= 1'b0;
    end else if(N862) begin
      btb_q[3960] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3959] <= 1'b0;
    end else if(N865) begin
      btb_q[3959] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3958] <= 1'b0;
    end else if(N865) begin
      btb_q[3958] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3957] <= 1'b0;
    end else if(N866) begin
      btb_q[3957] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3956] <= 1'b0;
    end else if(N866) begin
      btb_q[3956] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3955] <= 1'b0;
    end else if(N866) begin
      btb_q[3955] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3954] <= 1'b0;
    end else if(N866) begin
      btb_q[3954] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3953] <= 1'b0;
    end else if(N866) begin
      btb_q[3953] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3952] <= 1'b0;
    end else if(N866) begin
      btb_q[3952] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3951] <= 1'b0;
    end else if(N866) begin
      btb_q[3951] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3950] <= 1'b0;
    end else if(N866) begin
      btb_q[3950] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3949] <= 1'b0;
    end else if(N866) begin
      btb_q[3949] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3948] <= 1'b0;
    end else if(N866) begin
      btb_q[3948] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3947] <= 1'b0;
    end else if(N866) begin
      btb_q[3947] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3946] <= 1'b0;
    end else if(N866) begin
      btb_q[3946] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3945] <= 1'b0;
    end else if(N866) begin
      btb_q[3945] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3944] <= 1'b0;
    end else if(N866) begin
      btb_q[3944] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3943] <= 1'b0;
    end else if(N866) begin
      btb_q[3943] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3942] <= 1'b0;
    end else if(N866) begin
      btb_q[3942] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3941] <= 1'b0;
    end else if(N866) begin
      btb_q[3941] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3940] <= 1'b0;
    end else if(N866) begin
      btb_q[3940] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3939] <= 1'b0;
    end else if(N866) begin
      btb_q[3939] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3938] <= 1'b0;
    end else if(N866) begin
      btb_q[3938] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3937] <= 1'b0;
    end else if(N866) begin
      btb_q[3937] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3936] <= 1'b0;
    end else if(N866) begin
      btb_q[3936] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3935] <= 1'b0;
    end else if(N866) begin
      btb_q[3935] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3934] <= 1'b0;
    end else if(N866) begin
      btb_q[3934] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3933] <= 1'b0;
    end else if(N866) begin
      btb_q[3933] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3932] <= 1'b0;
    end else if(N866) begin
      btb_q[3932] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3931] <= 1'b0;
    end else if(N866) begin
      btb_q[3931] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3930] <= 1'b0;
    end else if(N866) begin
      btb_q[3930] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3929] <= 1'b0;
    end else if(N866) begin
      btb_q[3929] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3928] <= 1'b0;
    end else if(N866) begin
      btb_q[3928] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3927] <= 1'b0;
    end else if(N866) begin
      btb_q[3927] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3926] <= 1'b0;
    end else if(N866) begin
      btb_q[3926] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3925] <= 1'b0;
    end else if(N866) begin
      btb_q[3925] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3924] <= 1'b0;
    end else if(N866) begin
      btb_q[3924] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3923] <= 1'b0;
    end else if(N866) begin
      btb_q[3923] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3922] <= 1'b0;
    end else if(N866) begin
      btb_q[3922] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3921] <= 1'b0;
    end else if(N866) begin
      btb_q[3921] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3920] <= 1'b0;
    end else if(N870) begin
      btb_q[3920] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3919] <= 1'b0;
    end else if(N870) begin
      btb_q[3919] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3918] <= 1'b0;
    end else if(N870) begin
      btb_q[3918] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3917] <= 1'b0;
    end else if(N870) begin
      btb_q[3917] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3916] <= 1'b0;
    end else if(N870) begin
      btb_q[3916] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3915] <= 1'b0;
    end else if(N870) begin
      btb_q[3915] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3914] <= 1'b0;
    end else if(N870) begin
      btb_q[3914] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3913] <= 1'b0;
    end else if(N870) begin
      btb_q[3913] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3912] <= 1'b0;
    end else if(N870) begin
      btb_q[3912] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3911] <= 1'b0;
    end else if(N870) begin
      btb_q[3911] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3910] <= 1'b0;
    end else if(N870) begin
      btb_q[3910] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3909] <= 1'b0;
    end else if(N870) begin
      btb_q[3909] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3908] <= 1'b0;
    end else if(N870) begin
      btb_q[3908] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3907] <= 1'b0;
    end else if(N870) begin
      btb_q[3907] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3906] <= 1'b0;
    end else if(N870) begin
      btb_q[3906] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3905] <= 1'b0;
    end else if(N870) begin
      btb_q[3905] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3904] <= 1'b0;
    end else if(N870) begin
      btb_q[3904] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3903] <= 1'b0;
    end else if(N870) begin
      btb_q[3903] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3902] <= 1'b0;
    end else if(N870) begin
      btb_q[3902] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3901] <= 1'b0;
    end else if(N870) begin
      btb_q[3901] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3900] <= 1'b0;
    end else if(N870) begin
      btb_q[3900] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3899] <= 1'b0;
    end else if(N871) begin
      btb_q[3899] <= N589;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3898] <= 1'b0;
    end else if(N875) begin
      btb_q[3898] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3897] <= 1'b0;
    end else if(N875) begin
      btb_q[3897] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3896] <= 1'b0;
    end else if(N875) begin
      btb_q[3896] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3895] <= 1'b0;
    end else if(N875) begin
      btb_q[3895] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3894] <= 1'b0;
    end else if(N875) begin
      btb_q[3894] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3893] <= 1'b0;
    end else if(N875) begin
      btb_q[3893] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3892] <= 1'b0;
    end else if(N875) begin
      btb_q[3892] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3891] <= 1'b0;
    end else if(N875) begin
      btb_q[3891] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3890] <= 1'b0;
    end else if(N875) begin
      btb_q[3890] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3889] <= 1'b0;
    end else if(N875) begin
      btb_q[3889] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3888] <= 1'b0;
    end else if(N875) begin
      btb_q[3888] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3887] <= 1'b0;
    end else if(N875) begin
      btb_q[3887] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3886] <= 1'b0;
    end else if(N875) begin
      btb_q[3886] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3885] <= 1'b0;
    end else if(N875) begin
      btb_q[3885] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3884] <= 1'b0;
    end else if(N875) begin
      btb_q[3884] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3883] <= 1'b0;
    end else if(N875) begin
      btb_q[3883] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3882] <= 1'b0;
    end else if(N875) begin
      btb_q[3882] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3881] <= 1'b0;
    end else if(N875) begin
      btb_q[3881] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3880] <= 1'b0;
    end else if(N875) begin
      btb_q[3880] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3879] <= 1'b0;
    end else if(N875) begin
      btb_q[3879] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3878] <= 1'b0;
    end else if(N875) begin
      btb_q[3878] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3877] <= 1'b0;
    end else if(N875) begin
      btb_q[3877] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3876] <= 1'b0;
    end else if(N875) begin
      btb_q[3876] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3875] <= 1'b0;
    end else if(N875) begin
      btb_q[3875] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3874] <= 1'b0;
    end else if(N875) begin
      btb_q[3874] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3873] <= 1'b0;
    end else if(N875) begin
      btb_q[3873] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3872] <= 1'b0;
    end else if(N875) begin
      btb_q[3872] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3871] <= 1'b0;
    end else if(N875) begin
      btb_q[3871] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3870] <= 1'b0;
    end else if(N875) begin
      btb_q[3870] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3869] <= 1'b0;
    end else if(N875) begin
      btb_q[3869] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3868] <= 1'b0;
    end else if(N875) begin
      btb_q[3868] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3867] <= 1'b0;
    end else if(N875) begin
      btb_q[3867] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3866] <= 1'b0;
    end else if(N875) begin
      btb_q[3866] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3865] <= 1'b0;
    end else if(N875) begin
      btb_q[3865] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3864] <= 1'b0;
    end else if(N875) begin
      btb_q[3864] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3863] <= 1'b0;
    end else if(N875) begin
      btb_q[3863] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3862] <= 1'b0;
    end else if(N875) begin
      btb_q[3862] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3861] <= 1'b0;
    end else if(N875) begin
      btb_q[3861] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3860] <= 1'b0;
    end else if(N878) begin
      btb_q[3860] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3859] <= 1'b0;
    end else if(N878) begin
      btb_q[3859] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3858] <= 1'b0;
    end else if(N878) begin
      btb_q[3858] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3857] <= 1'b0;
    end else if(N879) begin
      btb_q[3857] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3856] <= 1'b0;
    end else if(N879) begin
      btb_q[3856] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3855] <= 1'b0;
    end else if(N879) begin
      btb_q[3855] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3854] <= 1'b0;
    end else if(N879) begin
      btb_q[3854] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3853] <= 1'b0;
    end else if(N879) begin
      btb_q[3853] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3852] <= 1'b0;
    end else if(N879) begin
      btb_q[3852] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3851] <= 1'b0;
    end else if(N879) begin
      btb_q[3851] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3850] <= 1'b0;
    end else if(N879) begin
      btb_q[3850] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3849] <= 1'b0;
    end else if(N879) begin
      btb_q[3849] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3848] <= 1'b0;
    end else if(N879) begin
      btb_q[3848] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3847] <= 1'b0;
    end else if(N879) begin
      btb_q[3847] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3846] <= 1'b0;
    end else if(N879) begin
      btb_q[3846] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3845] <= 1'b0;
    end else if(N879) begin
      btb_q[3845] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3844] <= 1'b0;
    end else if(N879) begin
      btb_q[3844] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3843] <= 1'b0;
    end else if(N879) begin
      btb_q[3843] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3842] <= 1'b0;
    end else if(N879) begin
      btb_q[3842] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3841] <= 1'b0;
    end else if(N879) begin
      btb_q[3841] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3840] <= 1'b0;
    end else if(N879) begin
      btb_q[3840] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3839] <= 1'b0;
    end else if(N879) begin
      btb_q[3839] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3838] <= 1'b0;
    end else if(N879) begin
      btb_q[3838] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3837] <= 1'b0;
    end else if(N879) begin
      btb_q[3837] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3836] <= 1'b0;
    end else if(N879) begin
      btb_q[3836] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3835] <= 1'b0;
    end else if(N879) begin
      btb_q[3835] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3834] <= 1'b0;
    end else if(N880) begin
      btb_q[3834] <= N588;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3833] <= 1'b0;
    end else if(N884) begin
      btb_q[3833] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3832] <= 1'b0;
    end else if(N884) begin
      btb_q[3832] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3831] <= 1'b0;
    end else if(N884) begin
      btb_q[3831] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3830] <= 1'b0;
    end else if(N884) begin
      btb_q[3830] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3829] <= 1'b0;
    end else if(N884) begin
      btb_q[3829] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3828] <= 1'b0;
    end else if(N884) begin
      btb_q[3828] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3827] <= 1'b0;
    end else if(N884) begin
      btb_q[3827] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3826] <= 1'b0;
    end else if(N884) begin
      btb_q[3826] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3825] <= 1'b0;
    end else if(N884) begin
      btb_q[3825] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3824] <= 1'b0;
    end else if(N884) begin
      btb_q[3824] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3823] <= 1'b0;
    end else if(N884) begin
      btb_q[3823] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3822] <= 1'b0;
    end else if(N884) begin
      btb_q[3822] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3821] <= 1'b0;
    end else if(N884) begin
      btb_q[3821] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3820] <= 1'b0;
    end else if(N884) begin
      btb_q[3820] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3819] <= 1'b0;
    end else if(N888) begin
      btb_q[3819] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3818] <= 1'b0;
    end else if(N888) begin
      btb_q[3818] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3817] <= 1'b0;
    end else if(N888) begin
      btb_q[3817] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3816] <= 1'b0;
    end else if(N888) begin
      btb_q[3816] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3815] <= 1'b0;
    end else if(N888) begin
      btb_q[3815] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3814] <= 1'b0;
    end else if(N888) begin
      btb_q[3814] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3813] <= 1'b0;
    end else if(N888) begin
      btb_q[3813] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3812] <= 1'b0;
    end else if(N888) begin
      btb_q[3812] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3811] <= 1'b0;
    end else if(N888) begin
      btb_q[3811] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3810] <= 1'b0;
    end else if(N888) begin
      btb_q[3810] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3809] <= 1'b0;
    end else if(N888) begin
      btb_q[3809] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3808] <= 1'b0;
    end else if(N888) begin
      btb_q[3808] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3807] <= 1'b0;
    end else if(N888) begin
      btb_q[3807] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3806] <= 1'b0;
    end else if(N888) begin
      btb_q[3806] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3805] <= 1'b0;
    end else if(N888) begin
      btb_q[3805] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3804] <= 1'b0;
    end else if(N888) begin
      btb_q[3804] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3803] <= 1'b0;
    end else if(N888) begin
      btb_q[3803] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3802] <= 1'b0;
    end else if(N888) begin
      btb_q[3802] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3801] <= 1'b0;
    end else if(N888) begin
      btb_q[3801] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3800] <= 1'b0;
    end else if(N888) begin
      btb_q[3800] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3799] <= 1'b0;
    end else if(N888) begin
      btb_q[3799] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3798] <= 1'b0;
    end else if(N888) begin
      btb_q[3798] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3797] <= 1'b0;
    end else if(N888) begin
      btb_q[3797] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3796] <= 1'b0;
    end else if(N888) begin
      btb_q[3796] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3795] <= 1'b0;
    end else if(N888) begin
      btb_q[3795] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3794] <= 1'b0;
    end else if(N888) begin
      btb_q[3794] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3793] <= 1'b0;
    end else if(N888) begin
      btb_q[3793] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3792] <= 1'b0;
    end else if(N888) begin
      btb_q[3792] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3791] <= 1'b0;
    end else if(N888) begin
      btb_q[3791] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3790] <= 1'b0;
    end else if(N888) begin
      btb_q[3790] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3789] <= 1'b0;
    end else if(N888) begin
      btb_q[3789] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3788] <= 1'b0;
    end else if(N888) begin
      btb_q[3788] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3787] <= 1'b0;
    end else if(N888) begin
      btb_q[3787] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3786] <= 1'b0;
    end else if(N888) begin
      btb_q[3786] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3785] <= 1'b0;
    end else if(N888) begin
      btb_q[3785] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3784] <= 1'b0;
    end else if(N888) begin
      btb_q[3784] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3783] <= 1'b0;
    end else if(N888) begin
      btb_q[3783] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3782] <= 1'b0;
    end else if(N888) begin
      btb_q[3782] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3781] <= 1'b0;
    end else if(N888) begin
      btb_q[3781] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3780] <= 1'b0;
    end else if(N888) begin
      btb_q[3780] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3779] <= 1'b0;
    end else if(N888) begin
      btb_q[3779] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3778] <= 1'b0;
    end else if(N888) begin
      btb_q[3778] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3777] <= 1'b0;
    end else if(N888) begin
      btb_q[3777] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3776] <= 1'b0;
    end else if(N888) begin
      btb_q[3776] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3775] <= 1'b0;
    end else if(N888) begin
      btb_q[3775] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3774] <= 1'b0;
    end else if(N888) begin
      btb_q[3774] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3773] <= 1'b0;
    end else if(N888) begin
      btb_q[3773] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3772] <= 1'b0;
    end else if(N888) begin
      btb_q[3772] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3771] <= 1'b0;
    end else if(N888) begin
      btb_q[3771] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3770] <= 1'b0;
    end else if(N888) begin
      btb_q[3770] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3769] <= 1'b0;
    end else if(N880) begin
      btb_q[3769] <= N587;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3768] <= 1'b0;
    end else if(N892) begin
      btb_q[3768] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3767] <= 1'b0;
    end else if(N892) begin
      btb_q[3767] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3766] <= 1'b0;
    end else if(N892) begin
      btb_q[3766] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3765] <= 1'b0;
    end else if(N892) begin
      btb_q[3765] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3764] <= 1'b0;
    end else if(N892) begin
      btb_q[3764] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3763] <= 1'b0;
    end else if(N892) begin
      btb_q[3763] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3762] <= 1'b0;
    end else if(N892) begin
      btb_q[3762] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3761] <= 1'b0;
    end else if(N895) begin
      btb_q[3761] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3760] <= 1'b0;
    end else if(N895) begin
      btb_q[3760] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3759] <= 1'b0;
    end else if(N895) begin
      btb_q[3759] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3758] <= 1'b0;
    end else if(N895) begin
      btb_q[3758] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3757] <= 1'b0;
    end else if(N895) begin
      btb_q[3757] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3756] <= 1'b0;
    end else if(N896) begin
      btb_q[3756] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3755] <= 1'b0;
    end else if(N896) begin
      btb_q[3755] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3754] <= 1'b0;
    end else if(N896) begin
      btb_q[3754] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3753] <= 1'b0;
    end else if(N896) begin
      btb_q[3753] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3752] <= 1'b0;
    end else if(N896) begin
      btb_q[3752] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3751] <= 1'b0;
    end else if(N896) begin
      btb_q[3751] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3750] <= 1'b0;
    end else if(N896) begin
      btb_q[3750] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3749] <= 1'b0;
    end else if(N896) begin
      btb_q[3749] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3748] <= 1'b0;
    end else if(N896) begin
      btb_q[3748] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3747] <= 1'b0;
    end else if(N896) begin
      btb_q[3747] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3746] <= 1'b0;
    end else if(N896) begin
      btb_q[3746] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3745] <= 1'b0;
    end else if(N896) begin
      btb_q[3745] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3744] <= 1'b0;
    end else if(N896) begin
      btb_q[3744] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3743] <= 1'b0;
    end else if(N896) begin
      btb_q[3743] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3742] <= 1'b0;
    end else if(N896) begin
      btb_q[3742] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3741] <= 1'b0;
    end else if(N896) begin
      btb_q[3741] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3740] <= 1'b0;
    end else if(N896) begin
      btb_q[3740] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3739] <= 1'b0;
    end else if(N896) begin
      btb_q[3739] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3738] <= 1'b0;
    end else if(N896) begin
      btb_q[3738] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3737] <= 1'b0;
    end else if(N896) begin
      btb_q[3737] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3736] <= 1'b0;
    end else if(N896) begin
      btb_q[3736] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3735] <= 1'b0;
    end else if(N896) begin
      btb_q[3735] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3734] <= 1'b0;
    end else if(N896) begin
      btb_q[3734] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3733] <= 1'b0;
    end else if(N896) begin
      btb_q[3733] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3732] <= 1'b0;
    end else if(N896) begin
      btb_q[3732] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3731] <= 1'b0;
    end else if(N896) begin
      btb_q[3731] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3730] <= 1'b0;
    end else if(N896) begin
      btb_q[3730] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3729] <= 1'b0;
    end else if(N896) begin
      btb_q[3729] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3728] <= 1'b0;
    end else if(N896) begin
      btb_q[3728] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3727] <= 1'b0;
    end else if(N896) begin
      btb_q[3727] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3726] <= 1'b0;
    end else if(N896) begin
      btb_q[3726] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3725] <= 1'b0;
    end else if(N896) begin
      btb_q[3725] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3724] <= 1'b0;
    end else if(N896) begin
      btb_q[3724] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3723] <= 1'b0;
    end else if(N896) begin
      btb_q[3723] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3722] <= 1'b0;
    end else if(N896) begin
      btb_q[3722] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3721] <= 1'b0;
    end else if(N896) begin
      btb_q[3721] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3720] <= 1'b0;
    end else if(N896) begin
      btb_q[3720] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3719] <= 1'b0;
    end else if(N900) begin
      btb_q[3719] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3718] <= 1'b0;
    end else if(N900) begin
      btb_q[3718] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3717] <= 1'b0;
    end else if(N900) begin
      btb_q[3717] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3716] <= 1'b0;
    end else if(N900) begin
      btb_q[3716] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3715] <= 1'b0;
    end else if(N900) begin
      btb_q[3715] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3714] <= 1'b0;
    end else if(N900) begin
      btb_q[3714] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3713] <= 1'b0;
    end else if(N900) begin
      btb_q[3713] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3712] <= 1'b0;
    end else if(N900) begin
      btb_q[3712] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3711] <= 1'b0;
    end else if(N900) begin
      btb_q[3711] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3710] <= 1'b0;
    end else if(N900) begin
      btb_q[3710] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3709] <= 1'b0;
    end else if(N900) begin
      btb_q[3709] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3708] <= 1'b0;
    end else if(N900) begin
      btb_q[3708] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3707] <= 1'b0;
    end else if(N900) begin
      btb_q[3707] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3706] <= 1'b0;
    end else if(N900) begin
      btb_q[3706] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3705] <= 1'b0;
    end else if(N900) begin
      btb_q[3705] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3704] <= 1'b0;
    end else if(N901) begin
      btb_q[3704] <= N586;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3703] <= 1'b0;
    end else if(N905) begin
      btb_q[3703] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3702] <= 1'b0;
    end else if(N905) begin
      btb_q[3702] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3701] <= 1'b0;
    end else if(N905) begin
      btb_q[3701] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3700] <= 1'b0;
    end else if(N905) begin
      btb_q[3700] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3699] <= 1'b0;
    end else if(N905) begin
      btb_q[3699] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3698] <= 1'b0;
    end else if(N905) begin
      btb_q[3698] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3697] <= 1'b0;
    end else if(N905) begin
      btb_q[3697] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3696] <= 1'b0;
    end else if(N905) begin
      btb_q[3696] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3695] <= 1'b0;
    end else if(N905) begin
      btb_q[3695] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3694] <= 1'b0;
    end else if(N905) begin
      btb_q[3694] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3693] <= 1'b0;
    end else if(N905) begin
      btb_q[3693] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3692] <= 1'b0;
    end else if(N905) begin
      btb_q[3692] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3691] <= 1'b0;
    end else if(N905) begin
      btb_q[3691] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3690] <= 1'b0;
    end else if(N905) begin
      btb_q[3690] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3689] <= 1'b0;
    end else if(N905) begin
      btb_q[3689] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3688] <= 1'b0;
    end else if(N905) begin
      btb_q[3688] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3687] <= 1'b0;
    end else if(N905) begin
      btb_q[3687] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3686] <= 1'b0;
    end else if(N905) begin
      btb_q[3686] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3685] <= 1'b0;
    end else if(N905) begin
      btb_q[3685] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3684] <= 1'b0;
    end else if(N905) begin
      btb_q[3684] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3683] <= 1'b0;
    end else if(N905) begin
      btb_q[3683] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3682] <= 1'b0;
    end else if(N905) begin
      btb_q[3682] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3681] <= 1'b0;
    end else if(N905) begin
      btb_q[3681] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3680] <= 1'b0;
    end else if(N905) begin
      btb_q[3680] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3679] <= 1'b0;
    end else if(N905) begin
      btb_q[3679] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3678] <= 1'b0;
    end else if(N905) begin
      btb_q[3678] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3677] <= 1'b0;
    end else if(N905) begin
      btb_q[3677] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3676] <= 1'b0;
    end else if(N905) begin
      btb_q[3676] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3675] <= 1'b0;
    end else if(N905) begin
      btb_q[3675] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3674] <= 1'b0;
    end else if(N905) begin
      btb_q[3674] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3673] <= 1'b0;
    end else if(N905) begin
      btb_q[3673] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3672] <= 1'b0;
    end else if(N905) begin
      btb_q[3672] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3671] <= 1'b0;
    end else if(N905) begin
      btb_q[3671] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3670] <= 1'b0;
    end else if(N905) begin
      btb_q[3670] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3669] <= 1'b0;
    end else if(N905) begin
      btb_q[3669] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3668] <= 1'b0;
    end else if(N905) begin
      btb_q[3668] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3667] <= 1'b0;
    end else if(N905) begin
      btb_q[3667] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3666] <= 1'b0;
    end else if(N905) begin
      btb_q[3666] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3665] <= 1'b0;
    end else if(N905) begin
      btb_q[3665] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3664] <= 1'b0;
    end else if(N905) begin
      btb_q[3664] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3663] <= 1'b0;
    end else if(N905) begin
      btb_q[3663] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3662] <= 1'b0;
    end else if(N908) begin
      btb_q[3662] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3661] <= 1'b0;
    end else if(N908) begin
      btb_q[3661] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3660] <= 1'b0;
    end else if(N908) begin
      btb_q[3660] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3659] <= 1'b0;
    end else if(N908) begin
      btb_q[3659] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3658] <= 1'b0;
    end else if(N908) begin
      btb_q[3658] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3657] <= 1'b0;
    end else if(N908) begin
      btb_q[3657] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3656] <= 1'b0;
    end else if(N909) begin
      btb_q[3656] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3655] <= 1'b0;
    end else if(N909) begin
      btb_q[3655] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3654] <= 1'b0;
    end else if(N909) begin
      btb_q[3654] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3653] <= 1'b0;
    end else if(N909) begin
      btb_q[3653] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3652] <= 1'b0;
    end else if(N909) begin
      btb_q[3652] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3651] <= 1'b0;
    end else if(N909) begin
      btb_q[3651] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3650] <= 1'b0;
    end else if(N909) begin
      btb_q[3650] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3649] <= 1'b0;
    end else if(N909) begin
      btb_q[3649] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3648] <= 1'b0;
    end else if(N909) begin
      btb_q[3648] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3647] <= 1'b0;
    end else if(N909) begin
      btb_q[3647] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3646] <= 1'b0;
    end else if(N909) begin
      btb_q[3646] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3645] <= 1'b0;
    end else if(N909) begin
      btb_q[3645] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3644] <= 1'b0;
    end else if(N909) begin
      btb_q[3644] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3643] <= 1'b0;
    end else if(N909) begin
      btb_q[3643] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3642] <= 1'b0;
    end else if(N909) begin
      btb_q[3642] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3641] <= 1'b0;
    end else if(N909) begin
      btb_q[3641] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3640] <= 1'b0;
    end else if(N909) begin
      btb_q[3640] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3639] <= 1'b0;
    end else if(N910) begin
      btb_q[3639] <= N585;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3638] <= 1'b0;
    end else if(N914) begin
      btb_q[3638] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3637] <= 1'b0;
    end else if(N914) begin
      btb_q[3637] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3636] <= 1'b0;
    end else if(N914) begin
      btb_q[3636] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3635] <= 1'b0;
    end else if(N914) begin
      btb_q[3635] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3634] <= 1'b0;
    end else if(N914) begin
      btb_q[3634] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3633] <= 1'b0;
    end else if(N914) begin
      btb_q[3633] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3632] <= 1'b0;
    end else if(N914) begin
      btb_q[3632] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3631] <= 1'b0;
    end else if(N914) begin
      btb_q[3631] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3630] <= 1'b0;
    end else if(N914) begin
      btb_q[3630] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3629] <= 1'b0;
    end else if(N914) begin
      btb_q[3629] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3628] <= 1'b0;
    end else if(N914) begin
      btb_q[3628] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3627] <= 1'b0;
    end else if(N914) begin
      btb_q[3627] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3626] <= 1'b0;
    end else if(N914) begin
      btb_q[3626] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3625] <= 1'b0;
    end else if(N914) begin
      btb_q[3625] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3624] <= 1'b0;
    end else if(N914) begin
      btb_q[3624] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3623] <= 1'b0;
    end else if(N914) begin
      btb_q[3623] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3622] <= 1'b0;
    end else if(N914) begin
      btb_q[3622] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3621] <= 1'b0;
    end else if(N914) begin
      btb_q[3621] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3620] <= 1'b0;
    end else if(N914) begin
      btb_q[3620] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3619] <= 1'b0;
    end else if(N914) begin
      btb_q[3619] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3618] <= 1'b0;
    end else if(N918) begin
      btb_q[3618] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3617] <= 1'b0;
    end else if(N918) begin
      btb_q[3617] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3616] <= 1'b0;
    end else if(N918) begin
      btb_q[3616] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3615] <= 1'b0;
    end else if(N918) begin
      btb_q[3615] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3614] <= 1'b0;
    end else if(N918) begin
      btb_q[3614] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3613] <= 1'b0;
    end else if(N918) begin
      btb_q[3613] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3612] <= 1'b0;
    end else if(N918) begin
      btb_q[3612] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3611] <= 1'b0;
    end else if(N918) begin
      btb_q[3611] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3610] <= 1'b0;
    end else if(N918) begin
      btb_q[3610] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3609] <= 1'b0;
    end else if(N918) begin
      btb_q[3609] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3608] <= 1'b0;
    end else if(N918) begin
      btb_q[3608] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3607] <= 1'b0;
    end else if(N918) begin
      btb_q[3607] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3606] <= 1'b0;
    end else if(N918) begin
      btb_q[3606] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3605] <= 1'b0;
    end else if(N918) begin
      btb_q[3605] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3604] <= 1'b0;
    end else if(N918) begin
      btb_q[3604] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3603] <= 1'b0;
    end else if(N918) begin
      btb_q[3603] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3602] <= 1'b0;
    end else if(N918) begin
      btb_q[3602] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3601] <= 1'b0;
    end else if(N918) begin
      btb_q[3601] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3600] <= 1'b0;
    end else if(N918) begin
      btb_q[3600] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3599] <= 1'b0;
    end else if(N918) begin
      btb_q[3599] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3598] <= 1'b0;
    end else if(N918) begin
      btb_q[3598] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3597] <= 1'b0;
    end else if(N918) begin
      btb_q[3597] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3596] <= 1'b0;
    end else if(N918) begin
      btb_q[3596] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3595] <= 1'b0;
    end else if(N918) begin
      btb_q[3595] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3594] <= 1'b0;
    end else if(N918) begin
      btb_q[3594] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3593] <= 1'b0;
    end else if(N918) begin
      btb_q[3593] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3592] <= 1'b0;
    end else if(N918) begin
      btb_q[3592] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3591] <= 1'b0;
    end else if(N918) begin
      btb_q[3591] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3590] <= 1'b0;
    end else if(N918) begin
      btb_q[3590] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3589] <= 1'b0;
    end else if(N918) begin
      btb_q[3589] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3588] <= 1'b0;
    end else if(N918) begin
      btb_q[3588] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3587] <= 1'b0;
    end else if(N918) begin
      btb_q[3587] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3586] <= 1'b0;
    end else if(N918) begin
      btb_q[3586] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3585] <= 1'b0;
    end else if(N918) begin
      btb_q[3585] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3584] <= 1'b0;
    end else if(N918) begin
      btb_q[3584] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3583] <= 1'b0;
    end else if(N918) begin
      btb_q[3583] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3582] <= 1'b0;
    end else if(N918) begin
      btb_q[3582] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3581] <= 1'b0;
    end else if(N918) begin
      btb_q[3581] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3580] <= 1'b0;
    end else if(N918) begin
      btb_q[3580] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3579] <= 1'b0;
    end else if(N918) begin
      btb_q[3579] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3578] <= 1'b0;
    end else if(N918) begin
      btb_q[3578] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3577] <= 1'b0;
    end else if(N918) begin
      btb_q[3577] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3576] <= 1'b0;
    end else if(N918) begin
      btb_q[3576] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3575] <= 1'b0;
    end else if(N918) begin
      btb_q[3575] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3574] <= 1'b0;
    end else if(N910) begin
      btb_q[3574] <= N584;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3573] <= 1'b0;
    end else if(N922) begin
      btb_q[3573] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3572] <= 1'b0;
    end else if(N922) begin
      btb_q[3572] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3571] <= 1'b0;
    end else if(N922) begin
      btb_q[3571] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3570] <= 1'b0;
    end else if(N922) begin
      btb_q[3570] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3569] <= 1'b0;
    end else if(N922) begin
      btb_q[3569] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3568] <= 1'b0;
    end else if(N922) begin
      btb_q[3568] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3567] <= 1'b0;
    end else if(N922) begin
      btb_q[3567] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3566] <= 1'b0;
    end else if(N922) begin
      btb_q[3566] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3565] <= 1'b0;
    end else if(N922) begin
      btb_q[3565] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3564] <= 1'b0;
    end else if(N922) begin
      btb_q[3564] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3563] <= 1'b0;
    end else if(N925) begin
      btb_q[3563] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3562] <= 1'b0;
    end else if(N925) begin
      btb_q[3562] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3561] <= 1'b0;
    end else if(N925) begin
      btb_q[3561] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3560] <= 1'b0;
    end else if(N925) begin
      btb_q[3560] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3559] <= 1'b0;
    end else if(N925) begin
      btb_q[3559] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3558] <= 1'b0;
    end else if(N925) begin
      btb_q[3558] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3557] <= 1'b0;
    end else if(N925) begin
      btb_q[3557] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3556] <= 1'b0;
    end else if(N925) begin
      btb_q[3556] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3555] <= 1'b0;
    end else if(N926) begin
      btb_q[3555] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3554] <= 1'b0;
    end else if(N926) begin
      btb_q[3554] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3553] <= 1'b0;
    end else if(N926) begin
      btb_q[3553] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3552] <= 1'b0;
    end else if(N926) begin
      btb_q[3552] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3551] <= 1'b0;
    end else if(N926) begin
      btb_q[3551] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3550] <= 1'b0;
    end else if(N926) begin
      btb_q[3550] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3549] <= 1'b0;
    end else if(N926) begin
      btb_q[3549] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3548] <= 1'b0;
    end else if(N926) begin
      btb_q[3548] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3547] <= 1'b0;
    end else if(N926) begin
      btb_q[3547] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3546] <= 1'b0;
    end else if(N926) begin
      btb_q[3546] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3545] <= 1'b0;
    end else if(N926) begin
      btb_q[3545] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3544] <= 1'b0;
    end else if(N926) begin
      btb_q[3544] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3543] <= 1'b0;
    end else if(N926) begin
      btb_q[3543] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3542] <= 1'b0;
    end else if(N926) begin
      btb_q[3542] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3541] <= 1'b0;
    end else if(N926) begin
      btb_q[3541] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3540] <= 1'b0;
    end else if(N926) begin
      btb_q[3540] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3539] <= 1'b0;
    end else if(N926) begin
      btb_q[3539] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3538] <= 1'b0;
    end else if(N926) begin
      btb_q[3538] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3537] <= 1'b0;
    end else if(N926) begin
      btb_q[3537] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3536] <= 1'b0;
    end else if(N926) begin
      btb_q[3536] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3535] <= 1'b0;
    end else if(N926) begin
      btb_q[3535] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3534] <= 1'b0;
    end else if(N926) begin
      btb_q[3534] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3533] <= 1'b0;
    end else if(N926) begin
      btb_q[3533] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3532] <= 1'b0;
    end else if(N926) begin
      btb_q[3532] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3531] <= 1'b0;
    end else if(N926) begin
      btb_q[3531] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3530] <= 1'b0;
    end else if(N926) begin
      btb_q[3530] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3529] <= 1'b0;
    end else if(N926) begin
      btb_q[3529] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3528] <= 1'b0;
    end else if(N926) begin
      btb_q[3528] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3527] <= 1'b0;
    end else if(N926) begin
      btb_q[3527] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3526] <= 1'b0;
    end else if(N926) begin
      btb_q[3526] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3525] <= 1'b0;
    end else if(N926) begin
      btb_q[3525] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3524] <= 1'b0;
    end else if(N926) begin
      btb_q[3524] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3523] <= 1'b0;
    end else if(N926) begin
      btb_q[3523] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3522] <= 1'b0;
    end else if(N926) begin
      btb_q[3522] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3521] <= 1'b0;
    end else if(N926) begin
      btb_q[3521] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3520] <= 1'b0;
    end else if(N926) begin
      btb_q[3520] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3519] <= 1'b0;
    end else if(N926) begin
      btb_q[3519] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3518] <= 1'b0;
    end else if(N930) begin
      btb_q[3518] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3517] <= 1'b0;
    end else if(N930) begin
      btb_q[3517] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3516] <= 1'b0;
    end else if(N930) begin
      btb_q[3516] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3515] <= 1'b0;
    end else if(N930) begin
      btb_q[3515] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3514] <= 1'b0;
    end else if(N930) begin
      btb_q[3514] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3513] <= 1'b0;
    end else if(N930) begin
      btb_q[3513] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3512] <= 1'b0;
    end else if(N930) begin
      btb_q[3512] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3511] <= 1'b0;
    end else if(N930) begin
      btb_q[3511] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3510] <= 1'b0;
    end else if(N930) begin
      btb_q[3510] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3509] <= 1'b0;
    end else if(N931) begin
      btb_q[3509] <= N583;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3508] <= 1'b0;
    end else if(N935) begin
      btb_q[3508] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3507] <= 1'b0;
    end else if(N935) begin
      btb_q[3507] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3506] <= 1'b0;
    end else if(N935) begin
      btb_q[3506] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3505] <= 1'b0;
    end else if(N935) begin
      btb_q[3505] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3504] <= 1'b0;
    end else if(N935) begin
      btb_q[3504] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3503] <= 1'b0;
    end else if(N935) begin
      btb_q[3503] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3502] <= 1'b0;
    end else if(N935) begin
      btb_q[3502] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3501] <= 1'b0;
    end else if(N935) begin
      btb_q[3501] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3500] <= 1'b0;
    end else if(N935) begin
      btb_q[3500] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3499] <= 1'b0;
    end else if(N935) begin
      btb_q[3499] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3498] <= 1'b0;
    end else if(N935) begin
      btb_q[3498] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3497] <= 1'b0;
    end else if(N935) begin
      btb_q[3497] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3496] <= 1'b0;
    end else if(N935) begin
      btb_q[3496] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3495] <= 1'b0;
    end else if(N935) begin
      btb_q[3495] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3494] <= 1'b0;
    end else if(N935) begin
      btb_q[3494] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3493] <= 1'b0;
    end else if(N935) begin
      btb_q[3493] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3492] <= 1'b0;
    end else if(N935) begin
      btb_q[3492] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3491] <= 1'b0;
    end else if(N935) begin
      btb_q[3491] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3490] <= 1'b0;
    end else if(N935) begin
      btb_q[3490] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3489] <= 1'b0;
    end else if(N935) begin
      btb_q[3489] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3488] <= 1'b0;
    end else if(N935) begin
      btb_q[3488] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3487] <= 1'b0;
    end else if(N935) begin
      btb_q[3487] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3486] <= 1'b0;
    end else if(N935) begin
      btb_q[3486] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3485] <= 1'b0;
    end else if(N935) begin
      btb_q[3485] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3484] <= 1'b0;
    end else if(N935) begin
      btb_q[3484] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3483] <= 1'b0;
    end else if(N935) begin
      btb_q[3483] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3482] <= 1'b0;
    end else if(N935) begin
      btb_q[3482] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3481] <= 1'b0;
    end else if(N935) begin
      btb_q[3481] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3480] <= 1'b0;
    end else if(N935) begin
      btb_q[3480] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3479] <= 1'b0;
    end else if(N935) begin
      btb_q[3479] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3478] <= 1'b0;
    end else if(N935) begin
      btb_q[3478] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3477] <= 1'b0;
    end else if(N935) begin
      btb_q[3477] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3476] <= 1'b0;
    end else if(N935) begin
      btb_q[3476] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3475] <= 1'b0;
    end else if(N935) begin
      btb_q[3475] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3474] <= 1'b0;
    end else if(N935) begin
      btb_q[3474] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3473] <= 1'b0;
    end else if(N935) begin
      btb_q[3473] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3472] <= 1'b0;
    end else if(N935) begin
      btb_q[3472] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3471] <= 1'b0;
    end else if(N935) begin
      btb_q[3471] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3470] <= 1'b0;
    end else if(N935) begin
      btb_q[3470] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3469] <= 1'b0;
    end else if(N935) begin
      btb_q[3469] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3468] <= 1'b0;
    end else if(N935) begin
      btb_q[3468] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3467] <= 1'b0;
    end else if(N935) begin
      btb_q[3467] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3466] <= 1'b0;
    end else if(N935) begin
      btb_q[3466] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3465] <= 1'b0;
    end else if(N935) begin
      btb_q[3465] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3464] <= 1'b0;
    end else if(N938) begin
      btb_q[3464] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3463] <= 1'b0;
    end else if(N938) begin
      btb_q[3463] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3462] <= 1'b0;
    end else if(N938) begin
      btb_q[3462] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3461] <= 1'b0;
    end else if(N938) begin
      btb_q[3461] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3460] <= 1'b0;
    end else if(N938) begin
      btb_q[3460] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3459] <= 1'b0;
    end else if(N938) begin
      btb_q[3459] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3458] <= 1'b0;
    end else if(N938) begin
      btb_q[3458] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3457] <= 1'b0;
    end else if(N938) begin
      btb_q[3457] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3456] <= 1'b0;
    end else if(N938) begin
      btb_q[3456] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3455] <= 1'b0;
    end else if(N939) begin
      btb_q[3455] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3454] <= 1'b0;
    end else if(N939) begin
      btb_q[3454] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3453] <= 1'b0;
    end else if(N939) begin
      btb_q[3453] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3452] <= 1'b0;
    end else if(N939) begin
      btb_q[3452] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3451] <= 1'b0;
    end else if(N939) begin
      btb_q[3451] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3450] <= 1'b0;
    end else if(N939) begin
      btb_q[3450] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3449] <= 1'b0;
    end else if(N939) begin
      btb_q[3449] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3448] <= 1'b0;
    end else if(N939) begin
      btb_q[3448] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3447] <= 1'b0;
    end else if(N939) begin
      btb_q[3447] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3446] <= 1'b0;
    end else if(N939) begin
      btb_q[3446] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3445] <= 1'b0;
    end else if(N939) begin
      btb_q[3445] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3444] <= 1'b0;
    end else if(N940) begin
      btb_q[3444] <= N582;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3443] <= 1'b0;
    end else if(N944) begin
      btb_q[3443] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3442] <= 1'b0;
    end else if(N944) begin
      btb_q[3442] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3441] <= 1'b0;
    end else if(N944) begin
      btb_q[3441] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3440] <= 1'b0;
    end else if(N944) begin
      btb_q[3440] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3439] <= 1'b0;
    end else if(N944) begin
      btb_q[3439] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3438] <= 1'b0;
    end else if(N944) begin
      btb_q[3438] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3437] <= 1'b0;
    end else if(N944) begin
      btb_q[3437] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3436] <= 1'b0;
    end else if(N944) begin
      btb_q[3436] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3435] <= 1'b0;
    end else if(N944) begin
      btb_q[3435] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3434] <= 1'b0;
    end else if(N944) begin
      btb_q[3434] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3433] <= 1'b0;
    end else if(N944) begin
      btb_q[3433] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3432] <= 1'b0;
    end else if(N944) begin
      btb_q[3432] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3431] <= 1'b0;
    end else if(N944) begin
      btb_q[3431] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3430] <= 1'b0;
    end else if(N944) begin
      btb_q[3430] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3429] <= 1'b0;
    end else if(N944) begin
      btb_q[3429] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3428] <= 1'b0;
    end else if(N944) begin
      btb_q[3428] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3427] <= 1'b0;
    end else if(N944) begin
      btb_q[3427] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3426] <= 1'b0;
    end else if(N944) begin
      btb_q[3426] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3425] <= 1'b0;
    end else if(N944) begin
      btb_q[3425] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3424] <= 1'b0;
    end else if(N944) begin
      btb_q[3424] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3423] <= 1'b0;
    end else if(N944) begin
      btb_q[3423] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3422] <= 1'b0;
    end else if(N944) begin
      btb_q[3422] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3421] <= 1'b0;
    end else if(N944) begin
      btb_q[3421] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3420] <= 1'b0;
    end else if(N944) begin
      btb_q[3420] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3419] <= 1'b0;
    end else if(N944) begin
      btb_q[3419] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3418] <= 1'b0;
    end else if(N944) begin
      btb_q[3418] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3417] <= 1'b0;
    end else if(N948) begin
      btb_q[3417] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3416] <= 1'b0;
    end else if(N948) begin
      btb_q[3416] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3415] <= 1'b0;
    end else if(N948) begin
      btb_q[3415] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3414] <= 1'b0;
    end else if(N948) begin
      btb_q[3414] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3413] <= 1'b0;
    end else if(N948) begin
      btb_q[3413] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3412] <= 1'b0;
    end else if(N948) begin
      btb_q[3412] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3411] <= 1'b0;
    end else if(N948) begin
      btb_q[3411] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3410] <= 1'b0;
    end else if(N948) begin
      btb_q[3410] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3409] <= 1'b0;
    end else if(N948) begin
      btb_q[3409] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3408] <= 1'b0;
    end else if(N948) begin
      btb_q[3408] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3407] <= 1'b0;
    end else if(N948) begin
      btb_q[3407] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3406] <= 1'b0;
    end else if(N948) begin
      btb_q[3406] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3405] <= 1'b0;
    end else if(N948) begin
      btb_q[3405] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3404] <= 1'b0;
    end else if(N948) begin
      btb_q[3404] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3403] <= 1'b0;
    end else if(N948) begin
      btb_q[3403] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3402] <= 1'b0;
    end else if(N948) begin
      btb_q[3402] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3401] <= 1'b0;
    end else if(N948) begin
      btb_q[3401] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3400] <= 1'b0;
    end else if(N948) begin
      btb_q[3400] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3399] <= 1'b0;
    end else if(N948) begin
      btb_q[3399] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3398] <= 1'b0;
    end else if(N948) begin
      btb_q[3398] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3397] <= 1'b0;
    end else if(N948) begin
      btb_q[3397] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3396] <= 1'b0;
    end else if(N948) begin
      btb_q[3396] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3395] <= 1'b0;
    end else if(N948) begin
      btb_q[3395] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3394] <= 1'b0;
    end else if(N948) begin
      btb_q[3394] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3393] <= 1'b0;
    end else if(N948) begin
      btb_q[3393] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3392] <= 1'b0;
    end else if(N948) begin
      btb_q[3392] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3391] <= 1'b0;
    end else if(N948) begin
      btb_q[3391] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3390] <= 1'b0;
    end else if(N948) begin
      btb_q[3390] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3389] <= 1'b0;
    end else if(N948) begin
      btb_q[3389] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3388] <= 1'b0;
    end else if(N948) begin
      btb_q[3388] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3387] <= 1'b0;
    end else if(N948) begin
      btb_q[3387] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3386] <= 1'b0;
    end else if(N948) begin
      btb_q[3386] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3385] <= 1'b0;
    end else if(N948) begin
      btb_q[3385] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3384] <= 1'b0;
    end else if(N948) begin
      btb_q[3384] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3383] <= 1'b0;
    end else if(N948) begin
      btb_q[3383] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3382] <= 1'b0;
    end else if(N948) begin
      btb_q[3382] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3381] <= 1'b0;
    end else if(N948) begin
      btb_q[3381] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3380] <= 1'b0;
    end else if(N948) begin
      btb_q[3380] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3379] <= 1'b0;
    end else if(N940) begin
      btb_q[3379] <= N581;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3378] <= 1'b0;
    end else if(N952) begin
      btb_q[3378] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3377] <= 1'b0;
    end else if(N952) begin
      btb_q[3377] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3376] <= 1'b0;
    end else if(N952) begin
      btb_q[3376] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3375] <= 1'b0;
    end else if(N952) begin
      btb_q[3375] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3374] <= 1'b0;
    end else if(N952) begin
      btb_q[3374] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3373] <= 1'b0;
    end else if(N952) begin
      btb_q[3373] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3372] <= 1'b0;
    end else if(N952) begin
      btb_q[3372] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3371] <= 1'b0;
    end else if(N952) begin
      btb_q[3371] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3370] <= 1'b0;
    end else if(N952) begin
      btb_q[3370] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3369] <= 1'b0;
    end else if(N952) begin
      btb_q[3369] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3368] <= 1'b0;
    end else if(N952) begin
      btb_q[3368] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3367] <= 1'b0;
    end else if(N952) begin
      btb_q[3367] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3366] <= 1'b0;
    end else if(N952) begin
      btb_q[3366] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3365] <= 1'b0;
    end else if(N955) begin
      btb_q[3365] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3364] <= 1'b0;
    end else if(N955) begin
      btb_q[3364] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3363] <= 1'b0;
    end else if(N955) begin
      btb_q[3363] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3362] <= 1'b0;
    end else if(N955) begin
      btb_q[3362] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3361] <= 1'b0;
    end else if(N955) begin
      btb_q[3361] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3360] <= 1'b0;
    end else if(N955) begin
      btb_q[3360] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3359] <= 1'b0;
    end else if(N955) begin
      btb_q[3359] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3358] <= 1'b0;
    end else if(N955) begin
      btb_q[3358] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3357] <= 1'b0;
    end else if(N955) begin
      btb_q[3357] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3356] <= 1'b0;
    end else if(N955) begin
      btb_q[3356] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3355] <= 1'b0;
    end else if(N955) begin
      btb_q[3355] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3354] <= 1'b0;
    end else if(N956) begin
      btb_q[3354] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3353] <= 1'b0;
    end else if(N956) begin
      btb_q[3353] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3352] <= 1'b0;
    end else if(N956) begin
      btb_q[3352] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3351] <= 1'b0;
    end else if(N956) begin
      btb_q[3351] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3350] <= 1'b0;
    end else if(N956) begin
      btb_q[3350] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3349] <= 1'b0;
    end else if(N956) begin
      btb_q[3349] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3348] <= 1'b0;
    end else if(N956) begin
      btb_q[3348] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3347] <= 1'b0;
    end else if(N956) begin
      btb_q[3347] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3346] <= 1'b0;
    end else if(N956) begin
      btb_q[3346] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3345] <= 1'b0;
    end else if(N956) begin
      btb_q[3345] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3344] <= 1'b0;
    end else if(N956) begin
      btb_q[3344] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3343] <= 1'b0;
    end else if(N956) begin
      btb_q[3343] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3342] <= 1'b0;
    end else if(N956) begin
      btb_q[3342] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3341] <= 1'b0;
    end else if(N956) begin
      btb_q[3341] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3340] <= 1'b0;
    end else if(N956) begin
      btb_q[3340] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3339] <= 1'b0;
    end else if(N956) begin
      btb_q[3339] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3338] <= 1'b0;
    end else if(N956) begin
      btb_q[3338] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3337] <= 1'b0;
    end else if(N956) begin
      btb_q[3337] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3336] <= 1'b0;
    end else if(N956) begin
      btb_q[3336] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3335] <= 1'b0;
    end else if(N956) begin
      btb_q[3335] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3334] <= 1'b0;
    end else if(N956) begin
      btb_q[3334] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3333] <= 1'b0;
    end else if(N956) begin
      btb_q[3333] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3332] <= 1'b0;
    end else if(N956) begin
      btb_q[3332] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3331] <= 1'b0;
    end else if(N956) begin
      btb_q[3331] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3330] <= 1'b0;
    end else if(N956) begin
      btb_q[3330] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3329] <= 1'b0;
    end else if(N956) begin
      btb_q[3329] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3328] <= 1'b0;
    end else if(N956) begin
      btb_q[3328] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3327] <= 1'b0;
    end else if(N956) begin
      btb_q[3327] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3326] <= 1'b0;
    end else if(N956) begin
      btb_q[3326] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3325] <= 1'b0;
    end else if(N956) begin
      btb_q[3325] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3324] <= 1'b0;
    end else if(N956) begin
      btb_q[3324] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3323] <= 1'b0;
    end else if(N956) begin
      btb_q[3323] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3322] <= 1'b0;
    end else if(N956) begin
      btb_q[3322] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3321] <= 1'b0;
    end else if(N956) begin
      btb_q[3321] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3320] <= 1'b0;
    end else if(N956) begin
      btb_q[3320] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3319] <= 1'b0;
    end else if(N956) begin
      btb_q[3319] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3318] <= 1'b0;
    end else if(N956) begin
      btb_q[3318] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3317] <= 1'b0;
    end else if(N960) begin
      btb_q[3317] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3316] <= 1'b0;
    end else if(N960) begin
      btb_q[3316] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3315] <= 1'b0;
    end else if(N960) begin
      btb_q[3315] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3314] <= 1'b0;
    end else if(N961) begin
      btb_q[3314] <= N580;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3313] <= 1'b0;
    end else if(N965) begin
      btb_q[3313] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3312] <= 1'b0;
    end else if(N965) begin
      btb_q[3312] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3311] <= 1'b0;
    end else if(N965) begin
      btb_q[3311] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3310] <= 1'b0;
    end else if(N965) begin
      btb_q[3310] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3309] <= 1'b0;
    end else if(N965) begin
      btb_q[3309] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3308] <= 1'b0;
    end else if(N965) begin
      btb_q[3308] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3307] <= 1'b0;
    end else if(N965) begin
      btb_q[3307] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3306] <= 1'b0;
    end else if(N965) begin
      btb_q[3306] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3305] <= 1'b0;
    end else if(N965) begin
      btb_q[3305] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3304] <= 1'b0;
    end else if(N965) begin
      btb_q[3304] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3303] <= 1'b0;
    end else if(N965) begin
      btb_q[3303] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3302] <= 1'b0;
    end else if(N965) begin
      btb_q[3302] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3301] <= 1'b0;
    end else if(N965) begin
      btb_q[3301] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3300] <= 1'b0;
    end else if(N965) begin
      btb_q[3300] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3299] <= 1'b0;
    end else if(N965) begin
      btb_q[3299] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3298] <= 1'b0;
    end else if(N965) begin
      btb_q[3298] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3297] <= 1'b0;
    end else if(N965) begin
      btb_q[3297] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3296] <= 1'b0;
    end else if(N965) begin
      btb_q[3296] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3295] <= 1'b0;
    end else if(N965) begin
      btb_q[3295] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3294] <= 1'b0;
    end else if(N965) begin
      btb_q[3294] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3293] <= 1'b0;
    end else if(N965) begin
      btb_q[3293] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3292] <= 1'b0;
    end else if(N965) begin
      btb_q[3292] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3291] <= 1'b0;
    end else if(N965) begin
      btb_q[3291] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3290] <= 1'b0;
    end else if(N965) begin
      btb_q[3290] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3289] <= 1'b0;
    end else if(N965) begin
      btb_q[3289] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3288] <= 1'b0;
    end else if(N965) begin
      btb_q[3288] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3287] <= 1'b0;
    end else if(N965) begin
      btb_q[3287] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3286] <= 1'b0;
    end else if(N965) begin
      btb_q[3286] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3285] <= 1'b0;
    end else if(N965) begin
      btb_q[3285] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3284] <= 1'b0;
    end else if(N965) begin
      btb_q[3284] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3283] <= 1'b0;
    end else if(N965) begin
      btb_q[3283] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3282] <= 1'b0;
    end else if(N965) begin
      btb_q[3282] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3281] <= 1'b0;
    end else if(N965) begin
      btb_q[3281] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3280] <= 1'b0;
    end else if(N965) begin
      btb_q[3280] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3279] <= 1'b0;
    end else if(N965) begin
      btb_q[3279] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3278] <= 1'b0;
    end else if(N965) begin
      btb_q[3278] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3277] <= 1'b0;
    end else if(N965) begin
      btb_q[3277] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3276] <= 1'b0;
    end else if(N965) begin
      btb_q[3276] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3275] <= 1'b0;
    end else if(N965) begin
      btb_q[3275] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3274] <= 1'b0;
    end else if(N965) begin
      btb_q[3274] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3273] <= 1'b0;
    end else if(N965) begin
      btb_q[3273] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3272] <= 1'b0;
    end else if(N965) begin
      btb_q[3272] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3271] <= 1'b0;
    end else if(N965) begin
      btb_q[3271] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3270] <= 1'b0;
    end else if(N965) begin
      btb_q[3270] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3269] <= 1'b0;
    end else if(N965) begin
      btb_q[3269] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3268] <= 1'b0;
    end else if(N965) begin
      btb_q[3268] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3267] <= 1'b0;
    end else if(N965) begin
      btb_q[3267] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3266] <= 1'b0;
    end else if(N968) begin
      btb_q[3266] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3265] <= 1'b0;
    end else if(N968) begin
      btb_q[3265] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3264] <= 1'b0;
    end else if(N968) begin
      btb_q[3264] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3263] <= 1'b0;
    end else if(N968) begin
      btb_q[3263] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3262] <= 1'b0;
    end else if(N968) begin
      btb_q[3262] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3261] <= 1'b0;
    end else if(N968) begin
      btb_q[3261] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3260] <= 1'b0;
    end else if(N968) begin
      btb_q[3260] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3259] <= 1'b0;
    end else if(N968) begin
      btb_q[3259] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3258] <= 1'b0;
    end else if(N968) begin
      btb_q[3258] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3257] <= 1'b0;
    end else if(N968) begin
      btb_q[3257] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3256] <= 1'b0;
    end else if(N968) begin
      btb_q[3256] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3255] <= 1'b0;
    end else if(N968) begin
      btb_q[3255] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3254] <= 1'b0;
    end else if(N969) begin
      btb_q[3254] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3253] <= 1'b0;
    end else if(N969) begin
      btb_q[3253] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3252] <= 1'b0;
    end else if(N969) begin
      btb_q[3252] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3251] <= 1'b0;
    end else if(N969) begin
      btb_q[3251] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3250] <= 1'b0;
    end else if(N969) begin
      btb_q[3250] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3249] <= 1'b0;
    end else if(N970) begin
      btb_q[3249] <= N579;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3248] <= 1'b0;
    end else if(N974) begin
      btb_q[3248] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3247] <= 1'b0;
    end else if(N974) begin
      btb_q[3247] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3246] <= 1'b0;
    end else if(N974) begin
      btb_q[3246] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3245] <= 1'b0;
    end else if(N974) begin
      btb_q[3245] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3244] <= 1'b0;
    end else if(N974) begin
      btb_q[3244] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3243] <= 1'b0;
    end else if(N974) begin
      btb_q[3243] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3242] <= 1'b0;
    end else if(N974) begin
      btb_q[3242] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3241] <= 1'b0;
    end else if(N974) begin
      btb_q[3241] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3240] <= 1'b0;
    end else if(N974) begin
      btb_q[3240] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3239] <= 1'b0;
    end else if(N974) begin
      btb_q[3239] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3238] <= 1'b0;
    end else if(N974) begin
      btb_q[3238] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3237] <= 1'b0;
    end else if(N974) begin
      btb_q[3237] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3236] <= 1'b0;
    end else if(N974) begin
      btb_q[3236] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3235] <= 1'b0;
    end else if(N974) begin
      btb_q[3235] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3234] <= 1'b0;
    end else if(N974) begin
      btb_q[3234] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3233] <= 1'b0;
    end else if(N974) begin
      btb_q[3233] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3232] <= 1'b0;
    end else if(N974) begin
      btb_q[3232] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3231] <= 1'b0;
    end else if(N974) begin
      btb_q[3231] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3230] <= 1'b0;
    end else if(N974) begin
      btb_q[3230] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3229] <= 1'b0;
    end else if(N974) begin
      btb_q[3229] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3228] <= 1'b0;
    end else if(N974) begin
      btb_q[3228] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3227] <= 1'b0;
    end else if(N974) begin
      btb_q[3227] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3226] <= 1'b0;
    end else if(N974) begin
      btb_q[3226] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3225] <= 1'b0;
    end else if(N974) begin
      btb_q[3225] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3224] <= 1'b0;
    end else if(N974) begin
      btb_q[3224] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3223] <= 1'b0;
    end else if(N974) begin
      btb_q[3223] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3222] <= 1'b0;
    end else if(N974) begin
      btb_q[3222] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3221] <= 1'b0;
    end else if(N974) begin
      btb_q[3221] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3220] <= 1'b0;
    end else if(N974) begin
      btb_q[3220] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3219] <= 1'b0;
    end else if(N974) begin
      btb_q[3219] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3218] <= 1'b0;
    end else if(N974) begin
      btb_q[3218] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3217] <= 1'b0;
    end else if(N974) begin
      btb_q[3217] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3216] <= 1'b0;
    end else if(N978) begin
      btb_q[3216] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3215] <= 1'b0;
    end else if(N978) begin
      btb_q[3215] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3214] <= 1'b0;
    end else if(N978) begin
      btb_q[3214] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3213] <= 1'b0;
    end else if(N978) begin
      btb_q[3213] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3212] <= 1'b0;
    end else if(N978) begin
      btb_q[3212] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3211] <= 1'b0;
    end else if(N978) begin
      btb_q[3211] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3210] <= 1'b0;
    end else if(N978) begin
      btb_q[3210] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3209] <= 1'b0;
    end else if(N978) begin
      btb_q[3209] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3208] <= 1'b0;
    end else if(N978) begin
      btb_q[3208] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3207] <= 1'b0;
    end else if(N978) begin
      btb_q[3207] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3206] <= 1'b0;
    end else if(N978) begin
      btb_q[3206] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3205] <= 1'b0;
    end else if(N978) begin
      btb_q[3205] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3204] <= 1'b0;
    end else if(N978) begin
      btb_q[3204] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3203] <= 1'b0;
    end else if(N978) begin
      btb_q[3203] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3202] <= 1'b0;
    end else if(N978) begin
      btb_q[3202] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3201] <= 1'b0;
    end else if(N978) begin
      btb_q[3201] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3200] <= 1'b0;
    end else if(N978) begin
      btb_q[3200] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3199] <= 1'b0;
    end else if(N978) begin
      btb_q[3199] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3198] <= 1'b0;
    end else if(N978) begin
      btb_q[3198] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3197] <= 1'b0;
    end else if(N978) begin
      btb_q[3197] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3196] <= 1'b0;
    end else if(N978) begin
      btb_q[3196] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3195] <= 1'b0;
    end else if(N978) begin
      btb_q[3195] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3194] <= 1'b0;
    end else if(N978) begin
      btb_q[3194] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3193] <= 1'b0;
    end else if(N978) begin
      btb_q[3193] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3192] <= 1'b0;
    end else if(N978) begin
      btb_q[3192] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3191] <= 1'b0;
    end else if(N978) begin
      btb_q[3191] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3190] <= 1'b0;
    end else if(N978) begin
      btb_q[3190] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3189] <= 1'b0;
    end else if(N978) begin
      btb_q[3189] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3188] <= 1'b0;
    end else if(N978) begin
      btb_q[3188] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3187] <= 1'b0;
    end else if(N978) begin
      btb_q[3187] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3186] <= 1'b0;
    end else if(N978) begin
      btb_q[3186] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3185] <= 1'b0;
    end else if(N978) begin
      btb_q[3185] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3184] <= 1'b0;
    end else if(N970) begin
      btb_q[3184] <= N578;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3183] <= 1'b0;
    end else if(N982) begin
      btb_q[3183] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3182] <= 1'b0;
    end else if(N982) begin
      btb_q[3182] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3181] <= 1'b0;
    end else if(N982) begin
      btb_q[3181] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3180] <= 1'b0;
    end else if(N982) begin
      btb_q[3180] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3179] <= 1'b0;
    end else if(N982) begin
      btb_q[3179] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3178] <= 1'b0;
    end else if(N982) begin
      btb_q[3178] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3177] <= 1'b0;
    end else if(N982) begin
      btb_q[3177] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3176] <= 1'b0;
    end else if(N982) begin
      btb_q[3176] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3175] <= 1'b0;
    end else if(N982) begin
      btb_q[3175] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3174] <= 1'b0;
    end else if(N982) begin
      btb_q[3174] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3173] <= 1'b0;
    end else if(N982) begin
      btb_q[3173] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3172] <= 1'b0;
    end else if(N982) begin
      btb_q[3172] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3171] <= 1'b0;
    end else if(N982) begin
      btb_q[3171] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3170] <= 1'b0;
    end else if(N982) begin
      btb_q[3170] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3169] <= 1'b0;
    end else if(N982) begin
      btb_q[3169] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3168] <= 1'b0;
    end else if(N982) begin
      btb_q[3168] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3167] <= 1'b0;
    end else if(N985) begin
      btb_q[3167] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3166] <= 1'b0;
    end else if(N985) begin
      btb_q[3166] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3165] <= 1'b0;
    end else if(N985) begin
      btb_q[3165] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3164] <= 1'b0;
    end else if(N985) begin
      btb_q[3164] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3163] <= 1'b0;
    end else if(N985) begin
      btb_q[3163] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3162] <= 1'b0;
    end else if(N985) begin
      btb_q[3162] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3161] <= 1'b0;
    end else if(N985) begin
      btb_q[3161] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3160] <= 1'b0;
    end else if(N985) begin
      btb_q[3160] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3159] <= 1'b0;
    end else if(N985) begin
      btb_q[3159] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3158] <= 1'b0;
    end else if(N985) begin
      btb_q[3158] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3157] <= 1'b0;
    end else if(N985) begin
      btb_q[3157] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3156] <= 1'b0;
    end else if(N985) begin
      btb_q[3156] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3155] <= 1'b0;
    end else if(N985) begin
      btb_q[3155] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3154] <= 1'b0;
    end else if(N985) begin
      btb_q[3154] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3153] <= 1'b0;
    end else if(N986) begin
      btb_q[3153] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3152] <= 1'b0;
    end else if(N986) begin
      btb_q[3152] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3151] <= 1'b0;
    end else if(N986) begin
      btb_q[3151] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3150] <= 1'b0;
    end else if(N986) begin
      btb_q[3150] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3149] <= 1'b0;
    end else if(N986) begin
      btb_q[3149] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3148] <= 1'b0;
    end else if(N986) begin
      btb_q[3148] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3147] <= 1'b0;
    end else if(N986) begin
      btb_q[3147] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3146] <= 1'b0;
    end else if(N986) begin
      btb_q[3146] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3145] <= 1'b0;
    end else if(N986) begin
      btb_q[3145] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3144] <= 1'b0;
    end else if(N986) begin
      btb_q[3144] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3143] <= 1'b0;
    end else if(N986) begin
      btb_q[3143] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3142] <= 1'b0;
    end else if(N986) begin
      btb_q[3142] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3141] <= 1'b0;
    end else if(N986) begin
      btb_q[3141] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3140] <= 1'b0;
    end else if(N986) begin
      btb_q[3140] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3139] <= 1'b0;
    end else if(N986) begin
      btb_q[3139] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3138] <= 1'b0;
    end else if(N986) begin
      btb_q[3138] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3137] <= 1'b0;
    end else if(N986) begin
      btb_q[3137] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3136] <= 1'b0;
    end else if(N986) begin
      btb_q[3136] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3135] <= 1'b0;
    end else if(N986) begin
      btb_q[3135] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3134] <= 1'b0;
    end else if(N986) begin
      btb_q[3134] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3133] <= 1'b0;
    end else if(N986) begin
      btb_q[3133] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3132] <= 1'b0;
    end else if(N986) begin
      btb_q[3132] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3131] <= 1'b0;
    end else if(N986) begin
      btb_q[3131] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3130] <= 1'b0;
    end else if(N986) begin
      btb_q[3130] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3129] <= 1'b0;
    end else if(N986) begin
      btb_q[3129] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3128] <= 1'b0;
    end else if(N986) begin
      btb_q[3128] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3127] <= 1'b0;
    end else if(N986) begin
      btb_q[3127] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3126] <= 1'b0;
    end else if(N986) begin
      btb_q[3126] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3125] <= 1'b0;
    end else if(N986) begin
      btb_q[3125] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3124] <= 1'b0;
    end else if(N986) begin
      btb_q[3124] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3123] <= 1'b0;
    end else if(N986) begin
      btb_q[3123] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3122] <= 1'b0;
    end else if(N986) begin
      btb_q[3122] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3121] <= 1'b0;
    end else if(N986) begin
      btb_q[3121] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3120] <= 1'b0;
    end else if(N986) begin
      btb_q[3120] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3119] <= 1'b0;
    end else if(N987) begin
      btb_q[3119] <= N577;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3118] <= 1'b0;
    end else if(N991) begin
      btb_q[3118] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3117] <= 1'b0;
    end else if(N991) begin
      btb_q[3117] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3116] <= 1'b0;
    end else if(N991) begin
      btb_q[3116] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3115] <= 1'b0;
    end else if(N995) begin
      btb_q[3115] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3114] <= 1'b0;
    end else if(N995) begin
      btb_q[3114] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3113] <= 1'b0;
    end else if(N995) begin
      btb_q[3113] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3112] <= 1'b0;
    end else if(N995) begin
      btb_q[3112] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3111] <= 1'b0;
    end else if(N995) begin
      btb_q[3111] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3110] <= 1'b0;
    end else if(N995) begin
      btb_q[3110] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3109] <= 1'b0;
    end else if(N995) begin
      btb_q[3109] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3108] <= 1'b0;
    end else if(N995) begin
      btb_q[3108] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3107] <= 1'b0;
    end else if(N995) begin
      btb_q[3107] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3106] <= 1'b0;
    end else if(N995) begin
      btb_q[3106] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3105] <= 1'b0;
    end else if(N995) begin
      btb_q[3105] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3104] <= 1'b0;
    end else if(N995) begin
      btb_q[3104] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3103] <= 1'b0;
    end else if(N995) begin
      btb_q[3103] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3102] <= 1'b0;
    end else if(N995) begin
      btb_q[3102] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3101] <= 1'b0;
    end else if(N995) begin
      btb_q[3101] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3100] <= 1'b0;
    end else if(N995) begin
      btb_q[3100] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3099] <= 1'b0;
    end else if(N995) begin
      btb_q[3099] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3098] <= 1'b0;
    end else if(N995) begin
      btb_q[3098] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3097] <= 1'b0;
    end else if(N995) begin
      btb_q[3097] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3096] <= 1'b0;
    end else if(N995) begin
      btb_q[3096] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3095] <= 1'b0;
    end else if(N995) begin
      btb_q[3095] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3094] <= 1'b0;
    end else if(N995) begin
      btb_q[3094] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3093] <= 1'b0;
    end else if(N995) begin
      btb_q[3093] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3092] <= 1'b0;
    end else if(N995) begin
      btb_q[3092] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3091] <= 1'b0;
    end else if(N995) begin
      btb_q[3091] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3090] <= 1'b0;
    end else if(N995) begin
      btb_q[3090] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3089] <= 1'b0;
    end else if(N995) begin
      btb_q[3089] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3088] <= 1'b0;
    end else if(N995) begin
      btb_q[3088] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3087] <= 1'b0;
    end else if(N995) begin
      btb_q[3087] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3086] <= 1'b0;
    end else if(N995) begin
      btb_q[3086] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3085] <= 1'b0;
    end else if(N995) begin
      btb_q[3085] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3084] <= 1'b0;
    end else if(N995) begin
      btb_q[3084] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3083] <= 1'b0;
    end else if(N995) begin
      btb_q[3083] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3082] <= 1'b0;
    end else if(N995) begin
      btb_q[3082] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3081] <= 1'b0;
    end else if(N995) begin
      btb_q[3081] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3080] <= 1'b0;
    end else if(N995) begin
      btb_q[3080] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3079] <= 1'b0;
    end else if(N995) begin
      btb_q[3079] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3078] <= 1'b0;
    end else if(N995) begin
      btb_q[3078] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3077] <= 1'b0;
    end else if(N995) begin
      btb_q[3077] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3076] <= 1'b0;
    end else if(N995) begin
      btb_q[3076] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3075] <= 1'b0;
    end else if(N995) begin
      btb_q[3075] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3074] <= 1'b0;
    end else if(N995) begin
      btb_q[3074] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3073] <= 1'b0;
    end else if(N995) begin
      btb_q[3073] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3072] <= 1'b0;
    end else if(N995) begin
      btb_q[3072] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3071] <= 1'b0;
    end else if(N995) begin
      btb_q[3071] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3070] <= 1'b0;
    end else if(N995) begin
      btb_q[3070] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3069] <= 1'b0;
    end else if(N995) begin
      btb_q[3069] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3068] <= 1'b0;
    end else if(N998) begin
      btb_q[3068] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3067] <= 1'b0;
    end else if(N998) begin
      btb_q[3067] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3066] <= 1'b0;
    end else if(N998) begin
      btb_q[3066] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3065] <= 1'b0;
    end else if(N998) begin
      btb_q[3065] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3064] <= 1'b0;
    end else if(N998) begin
      btb_q[3064] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3063] <= 1'b0;
    end else if(N998) begin
      btb_q[3063] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3062] <= 1'b0;
    end else if(N998) begin
      btb_q[3062] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3061] <= 1'b0;
    end else if(N998) begin
      btb_q[3061] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3060] <= 1'b0;
    end else if(N998) begin
      btb_q[3060] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3059] <= 1'b0;
    end else if(N998) begin
      btb_q[3059] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3058] <= 1'b0;
    end else if(N998) begin
      btb_q[3058] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3057] <= 1'b0;
    end else if(N998) begin
      btb_q[3057] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3056] <= 1'b0;
    end else if(N998) begin
      btb_q[3056] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3055] <= 1'b0;
    end else if(N998) begin
      btb_q[3055] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3054] <= 1'b0;
    end else if(N999) begin
      btb_q[3054] <= N576;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3053] <= 1'b0;
    end else if(N1003) begin
      btb_q[3053] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3052] <= 1'b0;
    end else if(N1004) begin
      btb_q[3052] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3051] <= 1'b0;
    end else if(N1004) begin
      btb_q[3051] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3050] <= 1'b0;
    end else if(N1004) begin
      btb_q[3050] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3049] <= 1'b0;
    end else if(N1004) begin
      btb_q[3049] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3048] <= 1'b0;
    end else if(N1004) begin
      btb_q[3048] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3047] <= 1'b0;
    end else if(N1004) begin
      btb_q[3047] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3046] <= 1'b0;
    end else if(N1004) begin
      btb_q[3046] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3045] <= 1'b0;
    end else if(N1004) begin
      btb_q[3045] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3044] <= 1'b0;
    end else if(N1004) begin
      btb_q[3044] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3043] <= 1'b0;
    end else if(N1004) begin
      btb_q[3043] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3042] <= 1'b0;
    end else if(N1004) begin
      btb_q[3042] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3041] <= 1'b0;
    end else if(N1004) begin
      btb_q[3041] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3040] <= 1'b0;
    end else if(N1004) begin
      btb_q[3040] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3039] <= 1'b0;
    end else if(N1004) begin
      btb_q[3039] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3038] <= 1'b0;
    end else if(N1004) begin
      btb_q[3038] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3037] <= 1'b0;
    end else if(N1004) begin
      btb_q[3037] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3036] <= 1'b0;
    end else if(N1004) begin
      btb_q[3036] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3035] <= 1'b0;
    end else if(N1004) begin
      btb_q[3035] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3034] <= 1'b0;
    end else if(N1004) begin
      btb_q[3034] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3033] <= 1'b0;
    end else if(N1004) begin
      btb_q[3033] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3032] <= 1'b0;
    end else if(N1004) begin
      btb_q[3032] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3031] <= 1'b0;
    end else if(N1004) begin
      btb_q[3031] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3030] <= 1'b0;
    end else if(N1004) begin
      btb_q[3030] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3029] <= 1'b0;
    end else if(N1004) begin
      btb_q[3029] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3028] <= 1'b0;
    end else if(N1004) begin
      btb_q[3028] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3027] <= 1'b0;
    end else if(N1004) begin
      btb_q[3027] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3026] <= 1'b0;
    end else if(N1004) begin
      btb_q[3026] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3025] <= 1'b0;
    end else if(N1004) begin
      btb_q[3025] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3024] <= 1'b0;
    end else if(N1004) begin
      btb_q[3024] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3023] <= 1'b0;
    end else if(N1004) begin
      btb_q[3023] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3022] <= 1'b0;
    end else if(N1004) begin
      btb_q[3022] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3021] <= 1'b0;
    end else if(N1004) begin
      btb_q[3021] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3020] <= 1'b0;
    end else if(N1004) begin
      btb_q[3020] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3019] <= 1'b0;
    end else if(N1004) begin
      btb_q[3019] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3018] <= 1'b0;
    end else if(N1004) begin
      btb_q[3018] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3017] <= 1'b0;
    end else if(N1004) begin
      btb_q[3017] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3016] <= 1'b0;
    end else if(N1004) begin
      btb_q[3016] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3015] <= 1'b0;
    end else if(N1008) begin
      btb_q[3015] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3014] <= 1'b0;
    end else if(N1008) begin
      btb_q[3014] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3013] <= 1'b0;
    end else if(N1008) begin
      btb_q[3013] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3012] <= 1'b0;
    end else if(N1008) begin
      btb_q[3012] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3011] <= 1'b0;
    end else if(N1008) begin
      btb_q[3011] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3010] <= 1'b0;
    end else if(N1008) begin
      btb_q[3010] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3009] <= 1'b0;
    end else if(N1008) begin
      btb_q[3009] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3008] <= 1'b0;
    end else if(N1008) begin
      btb_q[3008] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3007] <= 1'b0;
    end else if(N1008) begin
      btb_q[3007] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3006] <= 1'b0;
    end else if(N1008) begin
      btb_q[3006] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3005] <= 1'b0;
    end else if(N1008) begin
      btb_q[3005] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3004] <= 1'b0;
    end else if(N1008) begin
      btb_q[3004] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3003] <= 1'b0;
    end else if(N1008) begin
      btb_q[3003] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3002] <= 1'b0;
    end else if(N1008) begin
      btb_q[3002] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3001] <= 1'b0;
    end else if(N1008) begin
      btb_q[3001] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3000] <= 1'b0;
    end else if(N1008) begin
      btb_q[3000] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2999] <= 1'b0;
    end else if(N1008) begin
      btb_q[2999] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2998] <= 1'b0;
    end else if(N1008) begin
      btb_q[2998] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2997] <= 1'b0;
    end else if(N1008) begin
      btb_q[2997] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2996] <= 1'b0;
    end else if(N1008) begin
      btb_q[2996] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2995] <= 1'b0;
    end else if(N1008) begin
      btb_q[2995] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2994] <= 1'b0;
    end else if(N1008) begin
      btb_q[2994] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2993] <= 1'b0;
    end else if(N1008) begin
      btb_q[2993] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2992] <= 1'b0;
    end else if(N1008) begin
      btb_q[2992] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2991] <= 1'b0;
    end else if(N1008) begin
      btb_q[2991] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2990] <= 1'b0;
    end else if(N1008) begin
      btb_q[2990] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2989] <= 1'b0;
    end else if(N999) begin
      btb_q[2989] <= N575;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2988] <= 1'b0;
    end else if(N1012) begin
      btb_q[2988] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2987] <= 1'b0;
    end else if(N1012) begin
      btb_q[2987] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2986] <= 1'b0;
    end else if(N1012) begin
      btb_q[2986] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2985] <= 1'b0;
    end else if(N1012) begin
      btb_q[2985] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2984] <= 1'b0;
    end else if(N1012) begin
      btb_q[2984] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2983] <= 1'b0;
    end else if(N1012) begin
      btb_q[2983] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2982] <= 1'b0;
    end else if(N1012) begin
      btb_q[2982] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2981] <= 1'b0;
    end else if(N1012) begin
      btb_q[2981] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2980] <= 1'b0;
    end else if(N1012) begin
      btb_q[2980] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2979] <= 1'b0;
    end else if(N1012) begin
      btb_q[2979] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2978] <= 1'b0;
    end else if(N1012) begin
      btb_q[2978] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2977] <= 1'b0;
    end else if(N1012) begin
      btb_q[2977] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2976] <= 1'b0;
    end else if(N1012) begin
      btb_q[2976] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2975] <= 1'b0;
    end else if(N1012) begin
      btb_q[2975] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2974] <= 1'b0;
    end else if(N1012) begin
      btb_q[2974] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2973] <= 1'b0;
    end else if(N1012) begin
      btb_q[2973] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2972] <= 1'b0;
    end else if(N1012) begin
      btb_q[2972] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2971] <= 1'b0;
    end else if(N1012) begin
      btb_q[2971] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2970] <= 1'b0;
    end else if(N1012) begin
      btb_q[2970] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2969] <= 1'b0;
    end else if(N1015) begin
      btb_q[2969] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2968] <= 1'b0;
    end else if(N1015) begin
      btb_q[2968] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2967] <= 1'b0;
    end else if(N1015) begin
      btb_q[2967] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2966] <= 1'b0;
    end else if(N1015) begin
      btb_q[2966] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2965] <= 1'b0;
    end else if(N1015) begin
      btb_q[2965] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2964] <= 1'b0;
    end else if(N1015) begin
      btb_q[2964] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2963] <= 1'b0;
    end else if(N1015) begin
      btb_q[2963] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2962] <= 1'b0;
    end else if(N1015) begin
      btb_q[2962] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2961] <= 1'b0;
    end else if(N1015) begin
      btb_q[2961] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2960] <= 1'b0;
    end else if(N1015) begin
      btb_q[2960] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2959] <= 1'b0;
    end else if(N1015) begin
      btb_q[2959] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2958] <= 1'b0;
    end else if(N1015) begin
      btb_q[2958] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2957] <= 1'b0;
    end else if(N1015) begin
      btb_q[2957] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2956] <= 1'b0;
    end else if(N1015) begin
      btb_q[2956] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2955] <= 1'b0;
    end else if(N1015) begin
      btb_q[2955] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2954] <= 1'b0;
    end else if(N1015) begin
      btb_q[2954] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2953] <= 1'b0;
    end else if(N1015) begin
      btb_q[2953] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2952] <= 1'b0;
    end else if(N1016) begin
      btb_q[2952] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2951] <= 1'b0;
    end else if(N1016) begin
      btb_q[2951] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2950] <= 1'b0;
    end else if(N1016) begin
      btb_q[2950] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2949] <= 1'b0;
    end else if(N1016) begin
      btb_q[2949] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2948] <= 1'b0;
    end else if(N1016) begin
      btb_q[2948] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2947] <= 1'b0;
    end else if(N1016) begin
      btb_q[2947] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2946] <= 1'b0;
    end else if(N1016) begin
      btb_q[2946] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2945] <= 1'b0;
    end else if(N1016) begin
      btb_q[2945] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2944] <= 1'b0;
    end else if(N1016) begin
      btb_q[2944] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2943] <= 1'b0;
    end else if(N1016) begin
      btb_q[2943] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2942] <= 1'b0;
    end else if(N1016) begin
      btb_q[2942] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2941] <= 1'b0;
    end else if(N1016) begin
      btb_q[2941] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2940] <= 1'b0;
    end else if(N1016) begin
      btb_q[2940] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2939] <= 1'b0;
    end else if(N1016) begin
      btb_q[2939] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2938] <= 1'b0;
    end else if(N1016) begin
      btb_q[2938] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2937] <= 1'b0;
    end else if(N1016) begin
      btb_q[2937] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2936] <= 1'b0;
    end else if(N1016) begin
      btb_q[2936] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2935] <= 1'b0;
    end else if(N1016) begin
      btb_q[2935] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2934] <= 1'b0;
    end else if(N1016) begin
      btb_q[2934] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2933] <= 1'b0;
    end else if(N1016) begin
      btb_q[2933] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2932] <= 1'b0;
    end else if(N1016) begin
      btb_q[2932] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2931] <= 1'b0;
    end else if(N1016) begin
      btb_q[2931] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2930] <= 1'b0;
    end else if(N1016) begin
      btb_q[2930] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2929] <= 1'b0;
    end else if(N1016) begin
      btb_q[2929] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2928] <= 1'b0;
    end else if(N1016) begin
      btb_q[2928] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2927] <= 1'b0;
    end else if(N1016) begin
      btb_q[2927] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2926] <= 1'b0;
    end else if(N1016) begin
      btb_q[2926] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2925] <= 1'b0;
    end else if(N1016) begin
      btb_q[2925] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2924] <= 1'b0;
    end else if(N1017) begin
      btb_q[2924] <= N574;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2923] <= 1'b0;
    end else if(N1021) begin
      btb_q[2923] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2922] <= 1'b0;
    end else if(N1021) begin
      btb_q[2922] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2921] <= 1'b0;
    end else if(N1021) begin
      btb_q[2921] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2920] <= 1'b0;
    end else if(N1021) begin
      btb_q[2920] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2919] <= 1'b0;
    end else if(N1021) begin
      btb_q[2919] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2918] <= 1'b0;
    end else if(N1021) begin
      btb_q[2918] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2917] <= 1'b0;
    end else if(N1021) begin
      btb_q[2917] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2916] <= 1'b0;
    end else if(N1021) begin
      btb_q[2916] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2915] <= 1'b0;
    end else if(N1021) begin
      btb_q[2915] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2914] <= 1'b0;
    end else if(N1025) begin
      btb_q[2914] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2913] <= 1'b0;
    end else if(N1025) begin
      btb_q[2913] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2912] <= 1'b0;
    end else if(N1025) begin
      btb_q[2912] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2911] <= 1'b0;
    end else if(N1025) begin
      btb_q[2911] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2910] <= 1'b0;
    end else if(N1025) begin
      btb_q[2910] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2909] <= 1'b0;
    end else if(N1025) begin
      btb_q[2909] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2908] <= 1'b0;
    end else if(N1025) begin
      btb_q[2908] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2907] <= 1'b0;
    end else if(N1025) begin
      btb_q[2907] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2906] <= 1'b0;
    end else if(N1025) begin
      btb_q[2906] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2905] <= 1'b0;
    end else if(N1025) begin
      btb_q[2905] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2904] <= 1'b0;
    end else if(N1025) begin
      btb_q[2904] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2903] <= 1'b0;
    end else if(N1025) begin
      btb_q[2903] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2902] <= 1'b0;
    end else if(N1025) begin
      btb_q[2902] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2901] <= 1'b0;
    end else if(N1025) begin
      btb_q[2901] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2900] <= 1'b0;
    end else if(N1025) begin
      btb_q[2900] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2899] <= 1'b0;
    end else if(N1025) begin
      btb_q[2899] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2898] <= 1'b0;
    end else if(N1025) begin
      btb_q[2898] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2897] <= 1'b0;
    end else if(N1025) begin
      btb_q[2897] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2896] <= 1'b0;
    end else if(N1025) begin
      btb_q[2896] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2895] <= 1'b0;
    end else if(N1025) begin
      btb_q[2895] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2894] <= 1'b0;
    end else if(N1025) begin
      btb_q[2894] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2893] <= 1'b0;
    end else if(N1025) begin
      btb_q[2893] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2892] <= 1'b0;
    end else if(N1025) begin
      btb_q[2892] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2891] <= 1'b0;
    end else if(N1025) begin
      btb_q[2891] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2890] <= 1'b0;
    end else if(N1025) begin
      btb_q[2890] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2889] <= 1'b0;
    end else if(N1025) begin
      btb_q[2889] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2888] <= 1'b0;
    end else if(N1025) begin
      btb_q[2888] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2887] <= 1'b0;
    end else if(N1025) begin
      btb_q[2887] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2886] <= 1'b0;
    end else if(N1025) begin
      btb_q[2886] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2885] <= 1'b0;
    end else if(N1025) begin
      btb_q[2885] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2884] <= 1'b0;
    end else if(N1025) begin
      btb_q[2884] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2883] <= 1'b0;
    end else if(N1025) begin
      btb_q[2883] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2882] <= 1'b0;
    end else if(N1025) begin
      btb_q[2882] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2881] <= 1'b0;
    end else if(N1025) begin
      btb_q[2881] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2880] <= 1'b0;
    end else if(N1025) begin
      btb_q[2880] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2879] <= 1'b0;
    end else if(N1025) begin
      btb_q[2879] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2878] <= 1'b0;
    end else if(N1025) begin
      btb_q[2878] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2877] <= 1'b0;
    end else if(N1025) begin
      btb_q[2877] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2876] <= 1'b0;
    end else if(N1025) begin
      btb_q[2876] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2875] <= 1'b0;
    end else if(N1025) begin
      btb_q[2875] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2874] <= 1'b0;
    end else if(N1025) begin
      btb_q[2874] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2873] <= 1'b0;
    end else if(N1025) begin
      btb_q[2873] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2872] <= 1'b0;
    end else if(N1025) begin
      btb_q[2872] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2871] <= 1'b0;
    end else if(N1025) begin
      btb_q[2871] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2870] <= 1'b0;
    end else if(N1028) begin
      btb_q[2870] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2869] <= 1'b0;
    end else if(N1028) begin
      btb_q[2869] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2868] <= 1'b0;
    end else if(N1028) begin
      btb_q[2868] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2867] <= 1'b0;
    end else if(N1028) begin
      btb_q[2867] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2866] <= 1'b0;
    end else if(N1028) begin
      btb_q[2866] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2865] <= 1'b0;
    end else if(N1028) begin
      btb_q[2865] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2864] <= 1'b0;
    end else if(N1028) begin
      btb_q[2864] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2863] <= 1'b0;
    end else if(N1028) begin
      btb_q[2863] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2862] <= 1'b0;
    end else if(N1028) begin
      btb_q[2862] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2861] <= 1'b0;
    end else if(N1028) begin
      btb_q[2861] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2860] <= 1'b0;
    end else if(N1028) begin
      btb_q[2860] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2859] <= 1'b0;
    end else if(N1029) begin
      btb_q[2859] <= N573;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2858] <= 1'b0;
    end else if(N1033) begin
      btb_q[2858] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2857] <= 1'b0;
    end else if(N1033) begin
      btb_q[2857] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2856] <= 1'b0;
    end else if(N1033) begin
      btb_q[2856] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2855] <= 1'b0;
    end else if(N1033) begin
      btb_q[2855] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2854] <= 1'b0;
    end else if(N1033) begin
      btb_q[2854] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2853] <= 1'b0;
    end else if(N1033) begin
      btb_q[2853] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2852] <= 1'b0;
    end else if(N1033) begin
      btb_q[2852] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2851] <= 1'b0;
    end else if(N1034) begin
      btb_q[2851] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2850] <= 1'b0;
    end else if(N1034) begin
      btb_q[2850] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2849] <= 1'b0;
    end else if(N1034) begin
      btb_q[2849] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2848] <= 1'b0;
    end else if(N1034) begin
      btb_q[2848] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2847] <= 1'b0;
    end else if(N1034) begin
      btb_q[2847] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2846] <= 1'b0;
    end else if(N1034) begin
      btb_q[2846] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2845] <= 1'b0;
    end else if(N1034) begin
      btb_q[2845] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2844] <= 1'b0;
    end else if(N1034) begin
      btb_q[2844] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2843] <= 1'b0;
    end else if(N1034) begin
      btb_q[2843] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2842] <= 1'b0;
    end else if(N1034) begin
      btb_q[2842] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2841] <= 1'b0;
    end else if(N1034) begin
      btb_q[2841] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2840] <= 1'b0;
    end else if(N1034) begin
      btb_q[2840] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2839] <= 1'b0;
    end else if(N1034) begin
      btb_q[2839] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2838] <= 1'b0;
    end else if(N1034) begin
      btb_q[2838] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2837] <= 1'b0;
    end else if(N1034) begin
      btb_q[2837] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2836] <= 1'b0;
    end else if(N1034) begin
      btb_q[2836] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2835] <= 1'b0;
    end else if(N1034) begin
      btb_q[2835] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2834] <= 1'b0;
    end else if(N1034) begin
      btb_q[2834] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2833] <= 1'b0;
    end else if(N1034) begin
      btb_q[2833] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2832] <= 1'b0;
    end else if(N1034) begin
      btb_q[2832] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2831] <= 1'b0;
    end else if(N1034) begin
      btb_q[2831] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2830] <= 1'b0;
    end else if(N1034) begin
      btb_q[2830] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2829] <= 1'b0;
    end else if(N1034) begin
      btb_q[2829] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2828] <= 1'b0;
    end else if(N1034) begin
      btb_q[2828] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2827] <= 1'b0;
    end else if(N1034) begin
      btb_q[2827] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2826] <= 1'b0;
    end else if(N1034) begin
      btb_q[2826] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2825] <= 1'b0;
    end else if(N1034) begin
      btb_q[2825] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2824] <= 1'b0;
    end else if(N1034) begin
      btb_q[2824] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2823] <= 1'b0;
    end else if(N1034) begin
      btb_q[2823] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2822] <= 1'b0;
    end else if(N1034) begin
      btb_q[2822] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2821] <= 1'b0;
    end else if(N1034) begin
      btb_q[2821] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2820] <= 1'b0;
    end else if(N1034) begin
      btb_q[2820] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2819] <= 1'b0;
    end else if(N1034) begin
      btb_q[2819] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2818] <= 1'b0;
    end else if(N1034) begin
      btb_q[2818] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2817] <= 1'b0;
    end else if(N1034) begin
      btb_q[2817] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2816] <= 1'b0;
    end else if(N1034) begin
      btb_q[2816] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2815] <= 1'b0;
    end else if(N1034) begin
      btb_q[2815] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2814] <= 1'b0;
    end else if(N1038) begin
      btb_q[2814] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2813] <= 1'b0;
    end else if(N1038) begin
      btb_q[2813] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2812] <= 1'b0;
    end else if(N1038) begin
      btb_q[2812] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2811] <= 1'b0;
    end else if(N1038) begin
      btb_q[2811] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2810] <= 1'b0;
    end else if(N1038) begin
      btb_q[2810] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2809] <= 1'b0;
    end else if(N1038) begin
      btb_q[2809] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2808] <= 1'b0;
    end else if(N1038) begin
      btb_q[2808] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2807] <= 1'b0;
    end else if(N1038) begin
      btb_q[2807] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2806] <= 1'b0;
    end else if(N1038) begin
      btb_q[2806] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2805] <= 1'b0;
    end else if(N1038) begin
      btb_q[2805] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2804] <= 1'b0;
    end else if(N1038) begin
      btb_q[2804] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2803] <= 1'b0;
    end else if(N1038) begin
      btb_q[2803] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2802] <= 1'b0;
    end else if(N1038) begin
      btb_q[2802] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2801] <= 1'b0;
    end else if(N1038) begin
      btb_q[2801] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2800] <= 1'b0;
    end else if(N1038) begin
      btb_q[2800] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2799] <= 1'b0;
    end else if(N1038) begin
      btb_q[2799] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2798] <= 1'b0;
    end else if(N1038) begin
      btb_q[2798] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2797] <= 1'b0;
    end else if(N1038) begin
      btb_q[2797] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2796] <= 1'b0;
    end else if(N1038) begin
      btb_q[2796] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2795] <= 1'b0;
    end else if(N1038) begin
      btb_q[2795] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2794] <= 1'b0;
    end else if(N1029) begin
      btb_q[2794] <= N572;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2793] <= 1'b0;
    end else if(N1042) begin
      btb_q[2793] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2792] <= 1'b0;
    end else if(N1042) begin
      btb_q[2792] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2791] <= 1'b0;
    end else if(N1042) begin
      btb_q[2791] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2790] <= 1'b0;
    end else if(N1042) begin
      btb_q[2790] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2789] <= 1'b0;
    end else if(N1042) begin
      btb_q[2789] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2788] <= 1'b0;
    end else if(N1042) begin
      btb_q[2788] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2787] <= 1'b0;
    end else if(N1042) begin
      btb_q[2787] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2786] <= 1'b0;
    end else if(N1042) begin
      btb_q[2786] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2785] <= 1'b0;
    end else if(N1042) begin
      btb_q[2785] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2784] <= 1'b0;
    end else if(N1042) begin
      btb_q[2784] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2783] <= 1'b0;
    end else if(N1042) begin
      btb_q[2783] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2782] <= 1'b0;
    end else if(N1042) begin
      btb_q[2782] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2781] <= 1'b0;
    end else if(N1042) begin
      btb_q[2781] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2780] <= 1'b0;
    end else if(N1042) begin
      btb_q[2780] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2779] <= 1'b0;
    end else if(N1042) begin
      btb_q[2779] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2778] <= 1'b0;
    end else if(N1042) begin
      btb_q[2778] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2777] <= 1'b0;
    end else if(N1042) begin
      btb_q[2777] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2776] <= 1'b0;
    end else if(N1042) begin
      btb_q[2776] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2775] <= 1'b0;
    end else if(N1042) begin
      btb_q[2775] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2774] <= 1'b0;
    end else if(N1042) begin
      btb_q[2774] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2773] <= 1'b0;
    end else if(N1042) begin
      btb_q[2773] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2772] <= 1'b0;
    end else if(N1042) begin
      btb_q[2772] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2771] <= 1'b0;
    end else if(N1045) begin
      btb_q[2771] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2770] <= 1'b0;
    end else if(N1045) begin
      btb_q[2770] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2769] <= 1'b0;
    end else if(N1045) begin
      btb_q[2769] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2768] <= 1'b0;
    end else if(N1045) begin
      btb_q[2768] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2767] <= 1'b0;
    end else if(N1045) begin
      btb_q[2767] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2766] <= 1'b0;
    end else if(N1045) begin
      btb_q[2766] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2765] <= 1'b0;
    end else if(N1045) begin
      btb_q[2765] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2764] <= 1'b0;
    end else if(N1045) begin
      btb_q[2764] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2763] <= 1'b0;
    end else if(N1045) begin
      btb_q[2763] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2762] <= 1'b0;
    end else if(N1045) begin
      btb_q[2762] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2761] <= 1'b0;
    end else if(N1045) begin
      btb_q[2761] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2760] <= 1'b0;
    end else if(N1045) begin
      btb_q[2760] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2759] <= 1'b0;
    end else if(N1045) begin
      btb_q[2759] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2758] <= 1'b0;
    end else if(N1045) begin
      btb_q[2758] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2757] <= 1'b0;
    end else if(N1045) begin
      btb_q[2757] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2756] <= 1'b0;
    end else if(N1045) begin
      btb_q[2756] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2755] <= 1'b0;
    end else if(N1045) begin
      btb_q[2755] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2754] <= 1'b0;
    end else if(N1045) begin
      btb_q[2754] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2753] <= 1'b0;
    end else if(N1045) begin
      btb_q[2753] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2752] <= 1'b0;
    end else if(N1045) begin
      btb_q[2752] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2751] <= 1'b0;
    end else if(N1046) begin
      btb_q[2751] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2750] <= 1'b0;
    end else if(N1046) begin
      btb_q[2750] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2749] <= 1'b0;
    end else if(N1046) begin
      btb_q[2749] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2748] <= 1'b0;
    end else if(N1046) begin
      btb_q[2748] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2747] <= 1'b0;
    end else if(N1046) begin
      btb_q[2747] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2746] <= 1'b0;
    end else if(N1046) begin
      btb_q[2746] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2745] <= 1'b0;
    end else if(N1046) begin
      btb_q[2745] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2744] <= 1'b0;
    end else if(N1046) begin
      btb_q[2744] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2743] <= 1'b0;
    end else if(N1046) begin
      btb_q[2743] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2742] <= 1'b0;
    end else if(N1046) begin
      btb_q[2742] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2741] <= 1'b0;
    end else if(N1046) begin
      btb_q[2741] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2740] <= 1'b0;
    end else if(N1046) begin
      btb_q[2740] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2739] <= 1'b0;
    end else if(N1046) begin
      btb_q[2739] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2738] <= 1'b0;
    end else if(N1046) begin
      btb_q[2738] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2737] <= 1'b0;
    end else if(N1046) begin
      btb_q[2737] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2736] <= 1'b0;
    end else if(N1046) begin
      btb_q[2736] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2735] <= 1'b0;
    end else if(N1046) begin
      btb_q[2735] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2734] <= 1'b0;
    end else if(N1046) begin
      btb_q[2734] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2733] <= 1'b0;
    end else if(N1046) begin
      btb_q[2733] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2732] <= 1'b0;
    end else if(N1046) begin
      btb_q[2732] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2731] <= 1'b0;
    end else if(N1046) begin
      btb_q[2731] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2730] <= 1'b0;
    end else if(N1046) begin
      btb_q[2730] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2729] <= 1'b0;
    end else if(N1047) begin
      btb_q[2729] <= N571;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2728] <= 1'b0;
    end else if(N1051) begin
      btb_q[2728] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2727] <= 1'b0;
    end else if(N1051) begin
      btb_q[2727] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2726] <= 1'b0;
    end else if(N1051) begin
      btb_q[2726] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2725] <= 1'b0;
    end else if(N1051) begin
      btb_q[2725] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2724] <= 1'b0;
    end else if(N1051) begin
      btb_q[2724] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2723] <= 1'b0;
    end else if(N1051) begin
      btb_q[2723] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2722] <= 1'b0;
    end else if(N1051) begin
      btb_q[2722] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2721] <= 1'b0;
    end else if(N1051) begin
      btb_q[2721] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2720] <= 1'b0;
    end else if(N1051) begin
      btb_q[2720] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2719] <= 1'b0;
    end else if(N1051) begin
      btb_q[2719] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2718] <= 1'b0;
    end else if(N1051) begin
      btb_q[2718] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2717] <= 1'b0;
    end else if(N1051) begin
      btb_q[2717] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2716] <= 1'b0;
    end else if(N1051) begin
      btb_q[2716] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2715] <= 1'b0;
    end else if(N1051) begin
      btb_q[2715] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2714] <= 1'b0;
    end else if(N1051) begin
      btb_q[2714] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2713] <= 1'b0;
    end else if(N1055) begin
      btb_q[2713] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2712] <= 1'b0;
    end else if(N1055) begin
      btb_q[2712] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2711] <= 1'b0;
    end else if(N1055) begin
      btb_q[2711] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2710] <= 1'b0;
    end else if(N1055) begin
      btb_q[2710] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2709] <= 1'b0;
    end else if(N1055) begin
      btb_q[2709] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2708] <= 1'b0;
    end else if(N1055) begin
      btb_q[2708] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2707] <= 1'b0;
    end else if(N1055) begin
      btb_q[2707] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2706] <= 1'b0;
    end else if(N1055) begin
      btb_q[2706] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2705] <= 1'b0;
    end else if(N1055) begin
      btb_q[2705] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2704] <= 1'b0;
    end else if(N1055) begin
      btb_q[2704] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2703] <= 1'b0;
    end else if(N1055) begin
      btb_q[2703] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2702] <= 1'b0;
    end else if(N1055) begin
      btb_q[2702] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2701] <= 1'b0;
    end else if(N1055) begin
      btb_q[2701] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2700] <= 1'b0;
    end else if(N1055) begin
      btb_q[2700] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2699] <= 1'b0;
    end else if(N1055) begin
      btb_q[2699] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2698] <= 1'b0;
    end else if(N1055) begin
      btb_q[2698] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2697] <= 1'b0;
    end else if(N1055) begin
      btb_q[2697] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2696] <= 1'b0;
    end else if(N1055) begin
      btb_q[2696] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2695] <= 1'b0;
    end else if(N1055) begin
      btb_q[2695] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2694] <= 1'b0;
    end else if(N1055) begin
      btb_q[2694] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2693] <= 1'b0;
    end else if(N1055) begin
      btb_q[2693] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2692] <= 1'b0;
    end else if(N1055) begin
      btb_q[2692] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2691] <= 1'b0;
    end else if(N1055) begin
      btb_q[2691] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2690] <= 1'b0;
    end else if(N1055) begin
      btb_q[2690] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2689] <= 1'b0;
    end else if(N1055) begin
      btb_q[2689] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2688] <= 1'b0;
    end else if(N1055) begin
      btb_q[2688] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2687] <= 1'b0;
    end else if(N1055) begin
      btb_q[2687] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2686] <= 1'b0;
    end else if(N1055) begin
      btb_q[2686] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2685] <= 1'b0;
    end else if(N1055) begin
      btb_q[2685] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2684] <= 1'b0;
    end else if(N1055) begin
      btb_q[2684] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2683] <= 1'b0;
    end else if(N1055) begin
      btb_q[2683] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2682] <= 1'b0;
    end else if(N1055) begin
      btb_q[2682] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2681] <= 1'b0;
    end else if(N1055) begin
      btb_q[2681] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2680] <= 1'b0;
    end else if(N1055) begin
      btb_q[2680] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2679] <= 1'b0;
    end else if(N1055) begin
      btb_q[2679] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2678] <= 1'b0;
    end else if(N1055) begin
      btb_q[2678] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2677] <= 1'b0;
    end else if(N1055) begin
      btb_q[2677] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2676] <= 1'b0;
    end else if(N1055) begin
      btb_q[2676] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2675] <= 1'b0;
    end else if(N1055) begin
      btb_q[2675] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2674] <= 1'b0;
    end else if(N1055) begin
      btb_q[2674] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2673] <= 1'b0;
    end else if(N1055) begin
      btb_q[2673] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2672] <= 1'b0;
    end else if(N1058) begin
      btb_q[2672] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2671] <= 1'b0;
    end else if(N1058) begin
      btb_q[2671] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2670] <= 1'b0;
    end else if(N1058) begin
      btb_q[2670] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2669] <= 1'b0;
    end else if(N1058) begin
      btb_q[2669] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2668] <= 1'b0;
    end else if(N1058) begin
      btb_q[2668] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2667] <= 1'b0;
    end else if(N1058) begin
      btb_q[2667] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2666] <= 1'b0;
    end else if(N1058) begin
      btb_q[2666] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2665] <= 1'b0;
    end else if(N1058) begin
      btb_q[2665] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2664] <= 1'b0;
    end else if(N1059) begin
      btb_q[2664] <= N570;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2663] <= 1'b0;
    end else if(N1063) begin
      btb_q[2663] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2662] <= 1'b0;
    end else if(N1063) begin
      btb_q[2662] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2661] <= 1'b0;
    end else if(N1063) begin
      btb_q[2661] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2660] <= 1'b0;
    end else if(N1063) begin
      btb_q[2660] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2659] <= 1'b0;
    end else if(N1063) begin
      btb_q[2659] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2658] <= 1'b0;
    end else if(N1063) begin
      btb_q[2658] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2657] <= 1'b0;
    end else if(N1063) begin
      btb_q[2657] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2656] <= 1'b0;
    end else if(N1063) begin
      btb_q[2656] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2655] <= 1'b0;
    end else if(N1063) begin
      btb_q[2655] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2654] <= 1'b0;
    end else if(N1063) begin
      btb_q[2654] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2653] <= 1'b0;
    end else if(N1063) begin
      btb_q[2653] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2652] <= 1'b0;
    end else if(N1063) begin
      btb_q[2652] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2651] <= 1'b0;
    end else if(N1063) begin
      btb_q[2651] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2650] <= 1'b0;
    end else if(N1064) begin
      btb_q[2650] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2649] <= 1'b0;
    end else if(N1064) begin
      btb_q[2649] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2648] <= 1'b0;
    end else if(N1064) begin
      btb_q[2648] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2647] <= 1'b0;
    end else if(N1064) begin
      btb_q[2647] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2646] <= 1'b0;
    end else if(N1064) begin
      btb_q[2646] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2645] <= 1'b0;
    end else if(N1064) begin
      btb_q[2645] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2644] <= 1'b0;
    end else if(N1064) begin
      btb_q[2644] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2643] <= 1'b0;
    end else if(N1064) begin
      btb_q[2643] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2642] <= 1'b0;
    end else if(N1064) begin
      btb_q[2642] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2641] <= 1'b0;
    end else if(N1064) begin
      btb_q[2641] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2640] <= 1'b0;
    end else if(N1064) begin
      btb_q[2640] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2639] <= 1'b0;
    end else if(N1064) begin
      btb_q[2639] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2638] <= 1'b0;
    end else if(N1064) begin
      btb_q[2638] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2637] <= 1'b0;
    end else if(N1064) begin
      btb_q[2637] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2636] <= 1'b0;
    end else if(N1064) begin
      btb_q[2636] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2635] <= 1'b0;
    end else if(N1064) begin
      btb_q[2635] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2634] <= 1'b0;
    end else if(N1064) begin
      btb_q[2634] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2633] <= 1'b0;
    end else if(N1064) begin
      btb_q[2633] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2632] <= 1'b0;
    end else if(N1064) begin
      btb_q[2632] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2631] <= 1'b0;
    end else if(N1064) begin
      btb_q[2631] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2630] <= 1'b0;
    end else if(N1064) begin
      btb_q[2630] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2629] <= 1'b0;
    end else if(N1064) begin
      btb_q[2629] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2628] <= 1'b0;
    end else if(N1064) begin
      btb_q[2628] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2627] <= 1'b0;
    end else if(N1064) begin
      btb_q[2627] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2626] <= 1'b0;
    end else if(N1064) begin
      btb_q[2626] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2625] <= 1'b0;
    end else if(N1064) begin
      btb_q[2625] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2624] <= 1'b0;
    end else if(N1064) begin
      btb_q[2624] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2623] <= 1'b0;
    end else if(N1064) begin
      btb_q[2623] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2622] <= 1'b0;
    end else if(N1064) begin
      btb_q[2622] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2621] <= 1'b0;
    end else if(N1064) begin
      btb_q[2621] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2620] <= 1'b0;
    end else if(N1064) begin
      btb_q[2620] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2619] <= 1'b0;
    end else if(N1064) begin
      btb_q[2619] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2618] <= 1'b0;
    end else if(N1064) begin
      btb_q[2618] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2617] <= 1'b0;
    end else if(N1064) begin
      btb_q[2617] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2616] <= 1'b0;
    end else if(N1064) begin
      btb_q[2616] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2615] <= 1'b0;
    end else if(N1064) begin
      btb_q[2615] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2614] <= 1'b0;
    end else if(N1064) begin
      btb_q[2614] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2613] <= 1'b0;
    end else if(N1068) begin
      btb_q[2613] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2612] <= 1'b0;
    end else if(N1068) begin
      btb_q[2612] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2611] <= 1'b0;
    end else if(N1068) begin
      btb_q[2611] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2610] <= 1'b0;
    end else if(N1068) begin
      btb_q[2610] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2609] <= 1'b0;
    end else if(N1068) begin
      btb_q[2609] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2608] <= 1'b0;
    end else if(N1068) begin
      btb_q[2608] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2607] <= 1'b0;
    end else if(N1068) begin
      btb_q[2607] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2606] <= 1'b0;
    end else if(N1068) begin
      btb_q[2606] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2605] <= 1'b0;
    end else if(N1068) begin
      btb_q[2605] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2604] <= 1'b0;
    end else if(N1068) begin
      btb_q[2604] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2603] <= 1'b0;
    end else if(N1068) begin
      btb_q[2603] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2602] <= 1'b0;
    end else if(N1068) begin
      btb_q[2602] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2601] <= 1'b0;
    end else if(N1068) begin
      btb_q[2601] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2600] <= 1'b0;
    end else if(N1068) begin
      btb_q[2600] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2599] <= 1'b0;
    end else if(N1059) begin
      btb_q[2599] <= N569;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2598] <= 1'b0;
    end else if(N1072) begin
      btb_q[2598] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2597] <= 1'b0;
    end else if(N1072) begin
      btb_q[2597] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2596] <= 1'b0;
    end else if(N1072) begin
      btb_q[2596] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2595] <= 1'b0;
    end else if(N1072) begin
      btb_q[2595] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2594] <= 1'b0;
    end else if(N1072) begin
      btb_q[2594] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2593] <= 1'b0;
    end else if(N1072) begin
      btb_q[2593] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2592] <= 1'b0;
    end else if(N1072) begin
      btb_q[2592] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2591] <= 1'b0;
    end else if(N1072) begin
      btb_q[2591] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2590] <= 1'b0;
    end else if(N1072) begin
      btb_q[2590] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2589] <= 1'b0;
    end else if(N1072) begin
      btb_q[2589] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2588] <= 1'b0;
    end else if(N1072) begin
      btb_q[2588] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2587] <= 1'b0;
    end else if(N1072) begin
      btb_q[2587] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2586] <= 1'b0;
    end else if(N1072) begin
      btb_q[2586] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2585] <= 1'b0;
    end else if(N1072) begin
      btb_q[2585] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2584] <= 1'b0;
    end else if(N1072) begin
      btb_q[2584] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2583] <= 1'b0;
    end else if(N1072) begin
      btb_q[2583] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2582] <= 1'b0;
    end else if(N1072) begin
      btb_q[2582] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2581] <= 1'b0;
    end else if(N1072) begin
      btb_q[2581] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2580] <= 1'b0;
    end else if(N1072) begin
      btb_q[2580] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2579] <= 1'b0;
    end else if(N1072) begin
      btb_q[2579] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2578] <= 1'b0;
    end else if(N1072) begin
      btb_q[2578] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2577] <= 1'b0;
    end else if(N1072) begin
      btb_q[2577] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2576] <= 1'b0;
    end else if(N1072) begin
      btb_q[2576] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2575] <= 1'b0;
    end else if(N1072) begin
      btb_q[2575] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2574] <= 1'b0;
    end else if(N1072) begin
      btb_q[2574] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2573] <= 1'b0;
    end else if(N1075) begin
      btb_q[2573] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2572] <= 1'b0;
    end else if(N1075) begin
      btb_q[2572] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2571] <= 1'b0;
    end else if(N1075) begin
      btb_q[2571] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2570] <= 1'b0;
    end else if(N1075) begin
      btb_q[2570] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2569] <= 1'b0;
    end else if(N1075) begin
      btb_q[2569] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2568] <= 1'b0;
    end else if(N1075) begin
      btb_q[2568] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2567] <= 1'b0;
    end else if(N1075) begin
      btb_q[2567] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2566] <= 1'b0;
    end else if(N1075) begin
      btb_q[2566] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2565] <= 1'b0;
    end else if(N1075) begin
      btb_q[2565] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2564] <= 1'b0;
    end else if(N1075) begin
      btb_q[2564] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2563] <= 1'b0;
    end else if(N1075) begin
      btb_q[2563] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2562] <= 1'b0;
    end else if(N1075) begin
      btb_q[2562] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2561] <= 1'b0;
    end else if(N1075) begin
      btb_q[2561] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2560] <= 1'b0;
    end else if(N1075) begin
      btb_q[2560] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2559] <= 1'b0;
    end else if(N1075) begin
      btb_q[2559] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2558] <= 1'b0;
    end else if(N1075) begin
      btb_q[2558] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2557] <= 1'b0;
    end else if(N1075) begin
      btb_q[2557] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2556] <= 1'b0;
    end else if(N1075) begin
      btb_q[2556] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2555] <= 1'b0;
    end else if(N1075) begin
      btb_q[2555] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2554] <= 1'b0;
    end else if(N1075) begin
      btb_q[2554] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2553] <= 1'b0;
    end else if(N1075) begin
      btb_q[2553] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2552] <= 1'b0;
    end else if(N1075) begin
      btb_q[2552] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2551] <= 1'b0;
    end else if(N1075) begin
      btb_q[2551] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2550] <= 1'b0;
    end else if(N1076) begin
      btb_q[2550] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2549] <= 1'b0;
    end else if(N1076) begin
      btb_q[2549] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2548] <= 1'b0;
    end else if(N1076) begin
      btb_q[2548] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2547] <= 1'b0;
    end else if(N1076) begin
      btb_q[2547] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2546] <= 1'b0;
    end else if(N1076) begin
      btb_q[2546] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2545] <= 1'b0;
    end else if(N1076) begin
      btb_q[2545] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2544] <= 1'b0;
    end else if(N1076) begin
      btb_q[2544] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2543] <= 1'b0;
    end else if(N1076) begin
      btb_q[2543] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2542] <= 1'b0;
    end else if(N1076) begin
      btb_q[2542] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2541] <= 1'b0;
    end else if(N1076) begin
      btb_q[2541] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2540] <= 1'b0;
    end else if(N1076) begin
      btb_q[2540] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2539] <= 1'b0;
    end else if(N1076) begin
      btb_q[2539] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2538] <= 1'b0;
    end else if(N1076) begin
      btb_q[2538] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2537] <= 1'b0;
    end else if(N1076) begin
      btb_q[2537] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2536] <= 1'b0;
    end else if(N1076) begin
      btb_q[2536] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2535] <= 1'b0;
    end else if(N1076) begin
      btb_q[2535] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2534] <= 1'b0;
    end else if(N1077) begin
      btb_q[2534] <= N568;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2533] <= 1'b0;
    end else if(N1081) begin
      btb_q[2533] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2532] <= 1'b0;
    end else if(N1081) begin
      btb_q[2532] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2531] <= 1'b0;
    end else if(N1081) begin
      btb_q[2531] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2530] <= 1'b0;
    end else if(N1081) begin
      btb_q[2530] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2529] <= 1'b0;
    end else if(N1081) begin
      btb_q[2529] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2528] <= 1'b0;
    end else if(N1081) begin
      btb_q[2528] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2527] <= 1'b0;
    end else if(N1081) begin
      btb_q[2527] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2526] <= 1'b0;
    end else if(N1081) begin
      btb_q[2526] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2525] <= 1'b0;
    end else if(N1081) begin
      btb_q[2525] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2524] <= 1'b0;
    end else if(N1081) begin
      btb_q[2524] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2523] <= 1'b0;
    end else if(N1081) begin
      btb_q[2523] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2522] <= 1'b0;
    end else if(N1081) begin
      btb_q[2522] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2521] <= 1'b0;
    end else if(N1081) begin
      btb_q[2521] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2520] <= 1'b0;
    end else if(N1081) begin
      btb_q[2520] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2519] <= 1'b0;
    end else if(N1081) begin
      btb_q[2519] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2518] <= 1'b0;
    end else if(N1081) begin
      btb_q[2518] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2517] <= 1'b0;
    end else if(N1081) begin
      btb_q[2517] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2516] <= 1'b0;
    end else if(N1081) begin
      btb_q[2516] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2515] <= 1'b0;
    end else if(N1081) begin
      btb_q[2515] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2514] <= 1'b0;
    end else if(N1081) begin
      btb_q[2514] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2513] <= 1'b0;
    end else if(N1081) begin
      btb_q[2513] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2512] <= 1'b0;
    end else if(N1085) begin
      btb_q[2512] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2511] <= 1'b0;
    end else if(N1085) begin
      btb_q[2511] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2510] <= 1'b0;
    end else if(N1085) begin
      btb_q[2510] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2509] <= 1'b0;
    end else if(N1085) begin
      btb_q[2509] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2508] <= 1'b0;
    end else if(N1085) begin
      btb_q[2508] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2507] <= 1'b0;
    end else if(N1085) begin
      btb_q[2507] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2506] <= 1'b0;
    end else if(N1085) begin
      btb_q[2506] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2505] <= 1'b0;
    end else if(N1085) begin
      btb_q[2505] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2504] <= 1'b0;
    end else if(N1085) begin
      btb_q[2504] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2503] <= 1'b0;
    end else if(N1085) begin
      btb_q[2503] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2502] <= 1'b0;
    end else if(N1085) begin
      btb_q[2502] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2501] <= 1'b0;
    end else if(N1085) begin
      btb_q[2501] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2500] <= 1'b0;
    end else if(N1085) begin
      btb_q[2500] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2499] <= 1'b0;
    end else if(N1085) begin
      btb_q[2499] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2498] <= 1'b0;
    end else if(N1085) begin
      btb_q[2498] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2497] <= 1'b0;
    end else if(N1085) begin
      btb_q[2497] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2496] <= 1'b0;
    end else if(N1085) begin
      btb_q[2496] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2495] <= 1'b0;
    end else if(N1085) begin
      btb_q[2495] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2494] <= 1'b0;
    end else if(N1085) begin
      btb_q[2494] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2493] <= 1'b0;
    end else if(N1085) begin
      btb_q[2493] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2492] <= 1'b0;
    end else if(N1085) begin
      btb_q[2492] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2491] <= 1'b0;
    end else if(N1085) begin
      btb_q[2491] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2490] <= 1'b0;
    end else if(N1085) begin
      btb_q[2490] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2489] <= 1'b0;
    end else if(N1085) begin
      btb_q[2489] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2488] <= 1'b0;
    end else if(N1085) begin
      btb_q[2488] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2487] <= 1'b0;
    end else if(N1085) begin
      btb_q[2487] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2486] <= 1'b0;
    end else if(N1085) begin
      btb_q[2486] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2485] <= 1'b0;
    end else if(N1085) begin
      btb_q[2485] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2484] <= 1'b0;
    end else if(N1085) begin
      btb_q[2484] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2483] <= 1'b0;
    end else if(N1085) begin
      btb_q[2483] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2482] <= 1'b0;
    end else if(N1085) begin
      btb_q[2482] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2481] <= 1'b0;
    end else if(N1085) begin
      btb_q[2481] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2480] <= 1'b0;
    end else if(N1085) begin
      btb_q[2480] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2479] <= 1'b0;
    end else if(N1085) begin
      btb_q[2479] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2478] <= 1'b0;
    end else if(N1085) begin
      btb_q[2478] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2477] <= 1'b0;
    end else if(N1085) begin
      btb_q[2477] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2476] <= 1'b0;
    end else if(N1085) begin
      btb_q[2476] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2475] <= 1'b0;
    end else if(N1085) begin
      btb_q[2475] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2474] <= 1'b0;
    end else if(N1088) begin
      btb_q[2474] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2473] <= 1'b0;
    end else if(N1088) begin
      btb_q[2473] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2472] <= 1'b0;
    end else if(N1088) begin
      btb_q[2472] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2471] <= 1'b0;
    end else if(N1088) begin
      btb_q[2471] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2470] <= 1'b0;
    end else if(N1088) begin
      btb_q[2470] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2469] <= 1'b0;
    end else if(N1089) begin
      btb_q[2469] <= N567;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2468] <= 1'b0;
    end else if(N1093) begin
      btb_q[2468] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2467] <= 1'b0;
    end else if(N1093) begin
      btb_q[2467] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2466] <= 1'b0;
    end else if(N1093) begin
      btb_q[2466] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2465] <= 1'b0;
    end else if(N1093) begin
      btb_q[2465] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2464] <= 1'b0;
    end else if(N1093) begin
      btb_q[2464] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2463] <= 1'b0;
    end else if(N1093) begin
      btb_q[2463] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2462] <= 1'b0;
    end else if(N1093) begin
      btb_q[2462] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2461] <= 1'b0;
    end else if(N1093) begin
      btb_q[2461] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2460] <= 1'b0;
    end else if(N1093) begin
      btb_q[2460] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2459] <= 1'b0;
    end else if(N1093) begin
      btb_q[2459] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2458] <= 1'b0;
    end else if(N1093) begin
      btb_q[2458] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2457] <= 1'b0;
    end else if(N1093) begin
      btb_q[2457] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2456] <= 1'b0;
    end else if(N1093) begin
      btb_q[2456] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2455] <= 1'b0;
    end else if(N1093) begin
      btb_q[2455] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2454] <= 1'b0;
    end else if(N1093) begin
      btb_q[2454] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2453] <= 1'b0;
    end else if(N1093) begin
      btb_q[2453] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2452] <= 1'b0;
    end else if(N1093) begin
      btb_q[2452] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2451] <= 1'b0;
    end else if(N1093) begin
      btb_q[2451] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2450] <= 1'b0;
    end else if(N1093) begin
      btb_q[2450] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2449] <= 1'b0;
    end else if(N1094) begin
      btb_q[2449] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2448] <= 1'b0;
    end else if(N1094) begin
      btb_q[2448] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2447] <= 1'b0;
    end else if(N1094) begin
      btb_q[2447] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2446] <= 1'b0;
    end else if(N1094) begin
      btb_q[2446] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2445] <= 1'b0;
    end else if(N1094) begin
      btb_q[2445] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2444] <= 1'b0;
    end else if(N1094) begin
      btb_q[2444] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2443] <= 1'b0;
    end else if(N1094) begin
      btb_q[2443] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2442] <= 1'b0;
    end else if(N1094) begin
      btb_q[2442] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2441] <= 1'b0;
    end else if(N1094) begin
      btb_q[2441] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2440] <= 1'b0;
    end else if(N1094) begin
      btb_q[2440] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2439] <= 1'b0;
    end else if(N1094) begin
      btb_q[2439] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2438] <= 1'b0;
    end else if(N1094) begin
      btb_q[2438] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2437] <= 1'b0;
    end else if(N1094) begin
      btb_q[2437] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2436] <= 1'b0;
    end else if(N1094) begin
      btb_q[2436] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2435] <= 1'b0;
    end else if(N1094) begin
      btb_q[2435] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2434] <= 1'b0;
    end else if(N1094) begin
      btb_q[2434] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2433] <= 1'b0;
    end else if(N1094) begin
      btb_q[2433] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2432] <= 1'b0;
    end else if(N1094) begin
      btb_q[2432] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2431] <= 1'b0;
    end else if(N1094) begin
      btb_q[2431] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2430] <= 1'b0;
    end else if(N1094) begin
      btb_q[2430] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2429] <= 1'b0;
    end else if(N1094) begin
      btb_q[2429] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2428] <= 1'b0;
    end else if(N1094) begin
      btb_q[2428] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2427] <= 1'b0;
    end else if(N1094) begin
      btb_q[2427] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2426] <= 1'b0;
    end else if(N1094) begin
      btb_q[2426] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2425] <= 1'b0;
    end else if(N1094) begin
      btb_q[2425] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2424] <= 1'b0;
    end else if(N1094) begin
      btb_q[2424] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2423] <= 1'b0;
    end else if(N1094) begin
      btb_q[2423] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2422] <= 1'b0;
    end else if(N1094) begin
      btb_q[2422] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2421] <= 1'b0;
    end else if(N1094) begin
      btb_q[2421] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2420] <= 1'b0;
    end else if(N1094) begin
      btb_q[2420] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2419] <= 1'b0;
    end else if(N1094) begin
      btb_q[2419] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2418] <= 1'b0;
    end else if(N1094) begin
      btb_q[2418] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2417] <= 1'b0;
    end else if(N1094) begin
      btb_q[2417] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2416] <= 1'b0;
    end else if(N1094) begin
      btb_q[2416] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2415] <= 1'b0;
    end else if(N1094) begin
      btb_q[2415] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2414] <= 1'b0;
    end else if(N1094) begin
      btb_q[2414] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2413] <= 1'b0;
    end else if(N1094) begin
      btb_q[2413] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2412] <= 1'b0;
    end else if(N1098) begin
      btb_q[2412] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2411] <= 1'b0;
    end else if(N1098) begin
      btb_q[2411] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2410] <= 1'b0;
    end else if(N1098) begin
      btb_q[2410] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2409] <= 1'b0;
    end else if(N1098) begin
      btb_q[2409] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2408] <= 1'b0;
    end else if(N1098) begin
      btb_q[2408] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2407] <= 1'b0;
    end else if(N1098) begin
      btb_q[2407] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2406] <= 1'b0;
    end else if(N1098) begin
      btb_q[2406] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2405] <= 1'b0;
    end else if(N1098) begin
      btb_q[2405] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2404] <= 1'b0;
    end else if(N1089) begin
      btb_q[2404] <= N566;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2403] <= 1'b0;
    end else if(N1102) begin
      btb_q[2403] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2402] <= 1'b0;
    end else if(N1102) begin
      btb_q[2402] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2401] <= 1'b0;
    end else if(N1102) begin
      btb_q[2401] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2400] <= 1'b0;
    end else if(N1102) begin
      btb_q[2400] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2399] <= 1'b0;
    end else if(N1102) begin
      btb_q[2399] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2398] <= 1'b0;
    end else if(N1102) begin
      btb_q[2398] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2397] <= 1'b0;
    end else if(N1102) begin
      btb_q[2397] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2396] <= 1'b0;
    end else if(N1102) begin
      btb_q[2396] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2395] <= 1'b0;
    end else if(N1102) begin
      btb_q[2395] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2394] <= 1'b0;
    end else if(N1102) begin
      btb_q[2394] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2393] <= 1'b0;
    end else if(N1102) begin
      btb_q[2393] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2392] <= 1'b0;
    end else if(N1102) begin
      btb_q[2392] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2391] <= 1'b0;
    end else if(N1102) begin
      btb_q[2391] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2390] <= 1'b0;
    end else if(N1102) begin
      btb_q[2390] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2389] <= 1'b0;
    end else if(N1102) begin
      btb_q[2389] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2388] <= 1'b0;
    end else if(N1102) begin
      btb_q[2388] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2387] <= 1'b0;
    end else if(N1102) begin
      btb_q[2387] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2386] <= 1'b0;
    end else if(N1102) begin
      btb_q[2386] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2385] <= 1'b0;
    end else if(N1102) begin
      btb_q[2385] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2384] <= 1'b0;
    end else if(N1102) begin
      btb_q[2384] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2383] <= 1'b0;
    end else if(N1102) begin
      btb_q[2383] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2382] <= 1'b0;
    end else if(N1102) begin
      btb_q[2382] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2381] <= 1'b0;
    end else if(N1102) begin
      btb_q[2381] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2380] <= 1'b0;
    end else if(N1102) begin
      btb_q[2380] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2379] <= 1'b0;
    end else if(N1102) begin
      btb_q[2379] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2378] <= 1'b0;
    end else if(N1102) begin
      btb_q[2378] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2377] <= 1'b0;
    end else if(N1102) begin
      btb_q[2377] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2376] <= 1'b0;
    end else if(N1102) begin
      btb_q[2376] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2375] <= 1'b0;
    end else if(N1105) begin
      btb_q[2375] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2374] <= 1'b0;
    end else if(N1105) begin
      btb_q[2374] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2373] <= 1'b0;
    end else if(N1105) begin
      btb_q[2373] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2372] <= 1'b0;
    end else if(N1105) begin
      btb_q[2372] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2371] <= 1'b0;
    end else if(N1105) begin
      btb_q[2371] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2370] <= 1'b0;
    end else if(N1105) begin
      btb_q[2370] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2369] <= 1'b0;
    end else if(N1105) begin
      btb_q[2369] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2368] <= 1'b0;
    end else if(N1105) begin
      btb_q[2368] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2367] <= 1'b0;
    end else if(N1105) begin
      btb_q[2367] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2366] <= 1'b0;
    end else if(N1105) begin
      btb_q[2366] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2365] <= 1'b0;
    end else if(N1105) begin
      btb_q[2365] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2364] <= 1'b0;
    end else if(N1105) begin
      btb_q[2364] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2363] <= 1'b0;
    end else if(N1105) begin
      btb_q[2363] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2362] <= 1'b0;
    end else if(N1105) begin
      btb_q[2362] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2361] <= 1'b0;
    end else if(N1105) begin
      btb_q[2361] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2360] <= 1'b0;
    end else if(N1105) begin
      btb_q[2360] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2359] <= 1'b0;
    end else if(N1105) begin
      btb_q[2359] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2358] <= 1'b0;
    end else if(N1105) begin
      btb_q[2358] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2357] <= 1'b0;
    end else if(N1105) begin
      btb_q[2357] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2356] <= 1'b0;
    end else if(N1105) begin
      btb_q[2356] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2355] <= 1'b0;
    end else if(N1105) begin
      btb_q[2355] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2354] <= 1'b0;
    end else if(N1105) begin
      btb_q[2354] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2353] <= 1'b0;
    end else if(N1105) begin
      btb_q[2353] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2352] <= 1'b0;
    end else if(N1105) begin
      btb_q[2352] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2351] <= 1'b0;
    end else if(N1105) begin
      btb_q[2351] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2350] <= 1'b0;
    end else if(N1105) begin
      btb_q[2350] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2349] <= 1'b0;
    end else if(N1106) begin
      btb_q[2349] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2348] <= 1'b0;
    end else if(N1106) begin
      btb_q[2348] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2347] <= 1'b0;
    end else if(N1106) begin
      btb_q[2347] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2346] <= 1'b0;
    end else if(N1106) begin
      btb_q[2346] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2345] <= 1'b0;
    end else if(N1106) begin
      btb_q[2345] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2344] <= 1'b0;
    end else if(N1106) begin
      btb_q[2344] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2343] <= 1'b0;
    end else if(N1106) begin
      btb_q[2343] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2342] <= 1'b0;
    end else if(N1106) begin
      btb_q[2342] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2341] <= 1'b0;
    end else if(N1106) begin
      btb_q[2341] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2340] <= 1'b0;
    end else if(N1106) begin
      btb_q[2340] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2339] <= 1'b0;
    end else if(N1107) begin
      btb_q[2339] <= N565;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2338] <= 1'b0;
    end else if(N1111) begin
      btb_q[2338] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2337] <= 1'b0;
    end else if(N1111) begin
      btb_q[2337] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2336] <= 1'b0;
    end else if(N1111) begin
      btb_q[2336] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2335] <= 1'b0;
    end else if(N1111) begin
      btb_q[2335] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2334] <= 1'b0;
    end else if(N1111) begin
      btb_q[2334] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2333] <= 1'b0;
    end else if(N1111) begin
      btb_q[2333] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2332] <= 1'b0;
    end else if(N1111) begin
      btb_q[2332] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2331] <= 1'b0;
    end else if(N1111) begin
      btb_q[2331] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2330] <= 1'b0;
    end else if(N1111) begin
      btb_q[2330] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2329] <= 1'b0;
    end else if(N1111) begin
      btb_q[2329] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2328] <= 1'b0;
    end else if(N1111) begin
      btb_q[2328] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2327] <= 1'b0;
    end else if(N1111) begin
      btb_q[2327] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2326] <= 1'b0;
    end else if(N1111) begin
      btb_q[2326] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2325] <= 1'b0;
    end else if(N1111) begin
      btb_q[2325] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2324] <= 1'b0;
    end else if(N1111) begin
      btb_q[2324] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2323] <= 1'b0;
    end else if(N1111) begin
      btb_q[2323] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2322] <= 1'b0;
    end else if(N1111) begin
      btb_q[2322] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2321] <= 1'b0;
    end else if(N1111) begin
      btb_q[2321] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2320] <= 1'b0;
    end else if(N1111) begin
      btb_q[2320] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2319] <= 1'b0;
    end else if(N1111) begin
      btb_q[2319] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2318] <= 1'b0;
    end else if(N1111) begin
      btb_q[2318] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2317] <= 1'b0;
    end else if(N1111) begin
      btb_q[2317] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2316] <= 1'b0;
    end else if(N1111) begin
      btb_q[2316] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2315] <= 1'b0;
    end else if(N1111) begin
      btb_q[2315] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2314] <= 1'b0;
    end else if(N1111) begin
      btb_q[2314] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2313] <= 1'b0;
    end else if(N1111) begin
      btb_q[2313] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2312] <= 1'b0;
    end else if(N1111) begin
      btb_q[2312] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2311] <= 1'b0;
    end else if(N1115) begin
      btb_q[2311] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2310] <= 1'b0;
    end else if(N1115) begin
      btb_q[2310] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2309] <= 1'b0;
    end else if(N1115) begin
      btb_q[2309] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2308] <= 1'b0;
    end else if(N1115) begin
      btb_q[2308] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2307] <= 1'b0;
    end else if(N1115) begin
      btb_q[2307] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2306] <= 1'b0;
    end else if(N1115) begin
      btb_q[2306] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2305] <= 1'b0;
    end else if(N1115) begin
      btb_q[2305] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2304] <= 1'b0;
    end else if(N1115) begin
      btb_q[2304] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2303] <= 1'b0;
    end else if(N1115) begin
      btb_q[2303] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2302] <= 1'b0;
    end else if(N1115) begin
      btb_q[2302] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2301] <= 1'b0;
    end else if(N1115) begin
      btb_q[2301] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2300] <= 1'b0;
    end else if(N1115) begin
      btb_q[2300] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2299] <= 1'b0;
    end else if(N1115) begin
      btb_q[2299] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2298] <= 1'b0;
    end else if(N1115) begin
      btb_q[2298] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2297] <= 1'b0;
    end else if(N1115) begin
      btb_q[2297] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2296] <= 1'b0;
    end else if(N1115) begin
      btb_q[2296] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2295] <= 1'b0;
    end else if(N1115) begin
      btb_q[2295] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2294] <= 1'b0;
    end else if(N1115) begin
      btb_q[2294] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2293] <= 1'b0;
    end else if(N1115) begin
      btb_q[2293] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2292] <= 1'b0;
    end else if(N1115) begin
      btb_q[2292] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2291] <= 1'b0;
    end else if(N1115) begin
      btb_q[2291] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2290] <= 1'b0;
    end else if(N1115) begin
      btb_q[2290] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2289] <= 1'b0;
    end else if(N1115) begin
      btb_q[2289] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2288] <= 1'b0;
    end else if(N1115) begin
      btb_q[2288] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2287] <= 1'b0;
    end else if(N1115) begin
      btb_q[2287] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2286] <= 1'b0;
    end else if(N1115) begin
      btb_q[2286] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2285] <= 1'b0;
    end else if(N1115) begin
      btb_q[2285] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2284] <= 1'b0;
    end else if(N1115) begin
      btb_q[2284] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2283] <= 1'b0;
    end else if(N1115) begin
      btb_q[2283] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2282] <= 1'b0;
    end else if(N1115) begin
      btb_q[2282] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2281] <= 1'b0;
    end else if(N1115) begin
      btb_q[2281] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2280] <= 1'b0;
    end else if(N1115) begin
      btb_q[2280] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2279] <= 1'b0;
    end else if(N1115) begin
      btb_q[2279] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2278] <= 1'b0;
    end else if(N1115) begin
      btb_q[2278] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2277] <= 1'b0;
    end else if(N1115) begin
      btb_q[2277] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2276] <= 1'b0;
    end else if(N1118) begin
      btb_q[2276] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2275] <= 1'b0;
    end else if(N1118) begin
      btb_q[2275] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2274] <= 1'b0;
    end else if(N1119) begin
      btb_q[2274] <= N564;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2273] <= 1'b0;
    end else if(N1123) begin
      btb_q[2273] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2272] <= 1'b0;
    end else if(N1123) begin
      btb_q[2272] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2271] <= 1'b0;
    end else if(N1123) begin
      btb_q[2271] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2270] <= 1'b0;
    end else if(N1123) begin
      btb_q[2270] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2269] <= 1'b0;
    end else if(N1123) begin
      btb_q[2269] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2268] <= 1'b0;
    end else if(N1123) begin
      btb_q[2268] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2267] <= 1'b0;
    end else if(N1123) begin
      btb_q[2267] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2266] <= 1'b0;
    end else if(N1123) begin
      btb_q[2266] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2265] <= 1'b0;
    end else if(N1123) begin
      btb_q[2265] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2264] <= 1'b0;
    end else if(N1123) begin
      btb_q[2264] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2263] <= 1'b0;
    end else if(N1123) begin
      btb_q[2263] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2262] <= 1'b0;
    end else if(N1123) begin
      btb_q[2262] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2261] <= 1'b0;
    end else if(N1123) begin
      btb_q[2261] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2260] <= 1'b0;
    end else if(N1123) begin
      btb_q[2260] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2259] <= 1'b0;
    end else if(N1123) begin
      btb_q[2259] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2258] <= 1'b0;
    end else if(N1123) begin
      btb_q[2258] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2257] <= 1'b0;
    end else if(N1123) begin
      btb_q[2257] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2256] <= 1'b0;
    end else if(N1123) begin
      btb_q[2256] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2255] <= 1'b0;
    end else if(N1123) begin
      btb_q[2255] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2254] <= 1'b0;
    end else if(N1123) begin
      btb_q[2254] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2253] <= 1'b0;
    end else if(N1123) begin
      btb_q[2253] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2252] <= 1'b0;
    end else if(N1123) begin
      btb_q[2252] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2251] <= 1'b0;
    end else if(N1123) begin
      btb_q[2251] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2250] <= 1'b0;
    end else if(N1123) begin
      btb_q[2250] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2249] <= 1'b0;
    end else if(N1123) begin
      btb_q[2249] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2248] <= 1'b0;
    end else if(N1124) begin
      btb_q[2248] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2247] <= 1'b0;
    end else if(N1124) begin
      btb_q[2247] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2246] <= 1'b0;
    end else if(N1124) begin
      btb_q[2246] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2245] <= 1'b0;
    end else if(N1124) begin
      btb_q[2245] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2244] <= 1'b0;
    end else if(N1124) begin
      btb_q[2244] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2243] <= 1'b0;
    end else if(N1124) begin
      btb_q[2243] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2242] <= 1'b0;
    end else if(N1124) begin
      btb_q[2242] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2241] <= 1'b0;
    end else if(N1124) begin
      btb_q[2241] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2240] <= 1'b0;
    end else if(N1124) begin
      btb_q[2240] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2239] <= 1'b0;
    end else if(N1124) begin
      btb_q[2239] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2238] <= 1'b0;
    end else if(N1124) begin
      btb_q[2238] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2237] <= 1'b0;
    end else if(N1124) begin
      btb_q[2237] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2236] <= 1'b0;
    end else if(N1124) begin
      btb_q[2236] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2235] <= 1'b0;
    end else if(N1124) begin
      btb_q[2235] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2234] <= 1'b0;
    end else if(N1124) begin
      btb_q[2234] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2233] <= 1'b0;
    end else if(N1124) begin
      btb_q[2233] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2232] <= 1'b0;
    end else if(N1124) begin
      btb_q[2232] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2231] <= 1'b0;
    end else if(N1124) begin
      btb_q[2231] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2230] <= 1'b0;
    end else if(N1124) begin
      btb_q[2230] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2229] <= 1'b0;
    end else if(N1124) begin
      btb_q[2229] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2228] <= 1'b0;
    end else if(N1124) begin
      btb_q[2228] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2227] <= 1'b0;
    end else if(N1124) begin
      btb_q[2227] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2226] <= 1'b0;
    end else if(N1124) begin
      btb_q[2226] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2225] <= 1'b0;
    end else if(N1124) begin
      btb_q[2225] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2224] <= 1'b0;
    end else if(N1124) begin
      btb_q[2224] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2223] <= 1'b0;
    end else if(N1124) begin
      btb_q[2223] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2222] <= 1'b0;
    end else if(N1124) begin
      btb_q[2222] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2221] <= 1'b0;
    end else if(N1124) begin
      btb_q[2221] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2220] <= 1'b0;
    end else if(N1124) begin
      btb_q[2220] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2219] <= 1'b0;
    end else if(N1124) begin
      btb_q[2219] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2218] <= 1'b0;
    end else if(N1124) begin
      btb_q[2218] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2217] <= 1'b0;
    end else if(N1124) begin
      btb_q[2217] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2216] <= 1'b0;
    end else if(N1124) begin
      btb_q[2216] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2215] <= 1'b0;
    end else if(N1124) begin
      btb_q[2215] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2214] <= 1'b0;
    end else if(N1124) begin
      btb_q[2214] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2213] <= 1'b0;
    end else if(N1124) begin
      btb_q[2213] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2212] <= 1'b0;
    end else if(N1124) begin
      btb_q[2212] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2211] <= 1'b0;
    end else if(N1128) begin
      btb_q[2211] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2210] <= 1'b0;
    end else if(N1128) begin
      btb_q[2210] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2209] <= 1'b0;
    end else if(N1119) begin
      btb_q[2209] <= N563;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2208] <= 1'b0;
    end else if(N1132) begin
      btb_q[2208] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2207] <= 1'b0;
    end else if(N1132) begin
      btb_q[2207] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2206] <= 1'b0;
    end else if(N1132) begin
      btb_q[2206] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2205] <= 1'b0;
    end else if(N1132) begin
      btb_q[2205] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2204] <= 1'b0;
    end else if(N1132) begin
      btb_q[2204] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2203] <= 1'b0;
    end else if(N1132) begin
      btb_q[2203] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2202] <= 1'b0;
    end else if(N1132) begin
      btb_q[2202] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2201] <= 1'b0;
    end else if(N1132) begin
      btb_q[2201] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2200] <= 1'b0;
    end else if(N1132) begin
      btb_q[2200] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2199] <= 1'b0;
    end else if(N1132) begin
      btb_q[2199] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2198] <= 1'b0;
    end else if(N1132) begin
      btb_q[2198] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2197] <= 1'b0;
    end else if(N1132) begin
      btb_q[2197] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2196] <= 1'b0;
    end else if(N1132) begin
      btb_q[2196] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2195] <= 1'b0;
    end else if(N1132) begin
      btb_q[2195] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2194] <= 1'b0;
    end else if(N1132) begin
      btb_q[2194] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2193] <= 1'b0;
    end else if(N1132) begin
      btb_q[2193] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2192] <= 1'b0;
    end else if(N1132) begin
      btb_q[2192] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2191] <= 1'b0;
    end else if(N1132) begin
      btb_q[2191] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2190] <= 1'b0;
    end else if(N1132) begin
      btb_q[2190] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2189] <= 1'b0;
    end else if(N1132) begin
      btb_q[2189] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2188] <= 1'b0;
    end else if(N1132) begin
      btb_q[2188] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2187] <= 1'b0;
    end else if(N1132) begin
      btb_q[2187] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2186] <= 1'b0;
    end else if(N1132) begin
      btb_q[2186] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2185] <= 1'b0;
    end else if(N1132) begin
      btb_q[2185] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2184] <= 1'b0;
    end else if(N1132) begin
      btb_q[2184] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2183] <= 1'b0;
    end else if(N1132) begin
      btb_q[2183] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2182] <= 1'b0;
    end else if(N1132) begin
      btb_q[2182] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2181] <= 1'b0;
    end else if(N1132) begin
      btb_q[2181] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2180] <= 1'b0;
    end else if(N1132) begin
      btb_q[2180] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2179] <= 1'b0;
    end else if(N1132) begin
      btb_q[2179] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2178] <= 1'b0;
    end else if(N1132) begin
      btb_q[2178] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2177] <= 1'b0;
    end else if(N1135) begin
      btb_q[2177] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2176] <= 1'b0;
    end else if(N1135) begin
      btb_q[2176] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2175] <= 1'b0;
    end else if(N1135) begin
      btb_q[2175] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2174] <= 1'b0;
    end else if(N1135) begin
      btb_q[2174] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2173] <= 1'b0;
    end else if(N1135) begin
      btb_q[2173] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2172] <= 1'b0;
    end else if(N1135) begin
      btb_q[2172] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2171] <= 1'b0;
    end else if(N1135) begin
      btb_q[2171] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2170] <= 1'b0;
    end else if(N1135) begin
      btb_q[2170] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2169] <= 1'b0;
    end else if(N1135) begin
      btb_q[2169] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2168] <= 1'b0;
    end else if(N1135) begin
      btb_q[2168] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2167] <= 1'b0;
    end else if(N1135) begin
      btb_q[2167] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2166] <= 1'b0;
    end else if(N1135) begin
      btb_q[2166] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2165] <= 1'b0;
    end else if(N1135) begin
      btb_q[2165] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2164] <= 1'b0;
    end else if(N1135) begin
      btb_q[2164] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2163] <= 1'b0;
    end else if(N1135) begin
      btb_q[2163] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2162] <= 1'b0;
    end else if(N1135) begin
      btb_q[2162] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2161] <= 1'b0;
    end else if(N1135) begin
      btb_q[2161] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2160] <= 1'b0;
    end else if(N1135) begin
      btb_q[2160] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2159] <= 1'b0;
    end else if(N1135) begin
      btb_q[2159] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2158] <= 1'b0;
    end else if(N1135) begin
      btb_q[2158] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2157] <= 1'b0;
    end else if(N1135) begin
      btb_q[2157] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2156] <= 1'b0;
    end else if(N1135) begin
      btb_q[2156] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2155] <= 1'b0;
    end else if(N1135) begin
      btb_q[2155] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2154] <= 1'b0;
    end else if(N1135) begin
      btb_q[2154] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2153] <= 1'b0;
    end else if(N1135) begin
      btb_q[2153] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2152] <= 1'b0;
    end else if(N1135) begin
      btb_q[2152] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2151] <= 1'b0;
    end else if(N1135) begin
      btb_q[2151] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2150] <= 1'b0;
    end else if(N1135) begin
      btb_q[2150] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2149] <= 1'b0;
    end else if(N1135) begin
      btb_q[2149] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2148] <= 1'b0;
    end else if(N1136) begin
      btb_q[2148] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2147] <= 1'b0;
    end else if(N1136) begin
      btb_q[2147] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2146] <= 1'b0;
    end else if(N1136) begin
      btb_q[2146] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2145] <= 1'b0;
    end else if(N1136) begin
      btb_q[2145] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2144] <= 1'b0;
    end else if(N1137) begin
      btb_q[2144] <= N562;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2143] <= 1'b0;
    end else if(N1141) begin
      btb_q[2143] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2142] <= 1'b0;
    end else if(N1141) begin
      btb_q[2142] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2141] <= 1'b0;
    end else if(N1141) begin
      btb_q[2141] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2140] <= 1'b0;
    end else if(N1141) begin
      btb_q[2140] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2139] <= 1'b0;
    end else if(N1141) begin
      btb_q[2139] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2138] <= 1'b0;
    end else if(N1141) begin
      btb_q[2138] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2137] <= 1'b0;
    end else if(N1141) begin
      btb_q[2137] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2136] <= 1'b0;
    end else if(N1141) begin
      btb_q[2136] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2135] <= 1'b0;
    end else if(N1141) begin
      btb_q[2135] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2134] <= 1'b0;
    end else if(N1141) begin
      btb_q[2134] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2133] <= 1'b0;
    end else if(N1141) begin
      btb_q[2133] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2132] <= 1'b0;
    end else if(N1141) begin
      btb_q[2132] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2131] <= 1'b0;
    end else if(N1141) begin
      btb_q[2131] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2130] <= 1'b0;
    end else if(N1141) begin
      btb_q[2130] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2129] <= 1'b0;
    end else if(N1141) begin
      btb_q[2129] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2128] <= 1'b0;
    end else if(N1141) begin
      btb_q[2128] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2127] <= 1'b0;
    end else if(N1141) begin
      btb_q[2127] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2126] <= 1'b0;
    end else if(N1141) begin
      btb_q[2126] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2125] <= 1'b0;
    end else if(N1141) begin
      btb_q[2125] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2124] <= 1'b0;
    end else if(N1141) begin
      btb_q[2124] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2123] <= 1'b0;
    end else if(N1141) begin
      btb_q[2123] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2122] <= 1'b0;
    end else if(N1141) begin
      btb_q[2122] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2121] <= 1'b0;
    end else if(N1141) begin
      btb_q[2121] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2120] <= 1'b0;
    end else if(N1141) begin
      btb_q[2120] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2119] <= 1'b0;
    end else if(N1141) begin
      btb_q[2119] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2118] <= 1'b0;
    end else if(N1141) begin
      btb_q[2118] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2117] <= 1'b0;
    end else if(N1141) begin
      btb_q[2117] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2116] <= 1'b0;
    end else if(N1141) begin
      btb_q[2116] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2115] <= 1'b0;
    end else if(N1141) begin
      btb_q[2115] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2114] <= 1'b0;
    end else if(N1141) begin
      btb_q[2114] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2113] <= 1'b0;
    end else if(N1141) begin
      btb_q[2113] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2112] <= 1'b0;
    end else if(N1141) begin
      btb_q[2112] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2111] <= 1'b0;
    end else if(N1141) begin
      btb_q[2111] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2110] <= 1'b0;
    end else if(N1145) begin
      btb_q[2110] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2109] <= 1'b0;
    end else if(N1145) begin
      btb_q[2109] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2108] <= 1'b0;
    end else if(N1145) begin
      btb_q[2108] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2107] <= 1'b0;
    end else if(N1145) begin
      btb_q[2107] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2106] <= 1'b0;
    end else if(N1145) begin
      btb_q[2106] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2105] <= 1'b0;
    end else if(N1145) begin
      btb_q[2105] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2104] <= 1'b0;
    end else if(N1145) begin
      btb_q[2104] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2103] <= 1'b0;
    end else if(N1145) begin
      btb_q[2103] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2102] <= 1'b0;
    end else if(N1145) begin
      btb_q[2102] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2101] <= 1'b0;
    end else if(N1145) begin
      btb_q[2101] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2100] <= 1'b0;
    end else if(N1145) begin
      btb_q[2100] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2099] <= 1'b0;
    end else if(N1145) begin
      btb_q[2099] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2098] <= 1'b0;
    end else if(N1145) begin
      btb_q[2098] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2097] <= 1'b0;
    end else if(N1145) begin
      btb_q[2097] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2096] <= 1'b0;
    end else if(N1145) begin
      btb_q[2096] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2095] <= 1'b0;
    end else if(N1145) begin
      btb_q[2095] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2094] <= 1'b0;
    end else if(N1145) begin
      btb_q[2094] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2093] <= 1'b0;
    end else if(N1145) begin
      btb_q[2093] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2092] <= 1'b0;
    end else if(N1145) begin
      btb_q[2092] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2091] <= 1'b0;
    end else if(N1145) begin
      btb_q[2091] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2090] <= 1'b0;
    end else if(N1145) begin
      btb_q[2090] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2089] <= 1'b0;
    end else if(N1145) begin
      btb_q[2089] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2088] <= 1'b0;
    end else if(N1145) begin
      btb_q[2088] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2087] <= 1'b0;
    end else if(N1145) begin
      btb_q[2087] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2086] <= 1'b0;
    end else if(N1145) begin
      btb_q[2086] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2085] <= 1'b0;
    end else if(N1145) begin
      btb_q[2085] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2084] <= 1'b0;
    end else if(N1145) begin
      btb_q[2084] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2083] <= 1'b0;
    end else if(N1145) begin
      btb_q[2083] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2082] <= 1'b0;
    end else if(N1145) begin
      btb_q[2082] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2081] <= 1'b0;
    end else if(N1145) begin
      btb_q[2081] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2080] <= 1'b0;
    end else if(N1145) begin
      btb_q[2080] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2079] <= 1'b0;
    end else if(N1137) begin
      btb_q[2079] <= N561;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2078] <= 1'b0;
    end else if(N1149) begin
      btb_q[2078] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2077] <= 1'b0;
    end else if(N1149) begin
      btb_q[2077] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2076] <= 1'b0;
    end else if(N1149) begin
      btb_q[2076] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2075] <= 1'b0;
    end else if(N1149) begin
      btb_q[2075] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2074] <= 1'b0;
    end else if(N1149) begin
      btb_q[2074] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2073] <= 1'b0;
    end else if(N1149) begin
      btb_q[2073] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2072] <= 1'b0;
    end else if(N1149) begin
      btb_q[2072] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2071] <= 1'b0;
    end else if(N1149) begin
      btb_q[2071] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2070] <= 1'b0;
    end else if(N1149) begin
      btb_q[2070] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2069] <= 1'b0;
    end else if(N1149) begin
      btb_q[2069] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2068] <= 1'b0;
    end else if(N1149) begin
      btb_q[2068] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2067] <= 1'b0;
    end else if(N1149) begin
      btb_q[2067] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2066] <= 1'b0;
    end else if(N1149) begin
      btb_q[2066] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2065] <= 1'b0;
    end else if(N1149) begin
      btb_q[2065] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2064] <= 1'b0;
    end else if(N1149) begin
      btb_q[2064] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2063] <= 1'b0;
    end else if(N1149) begin
      btb_q[2063] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2062] <= 1'b0;
    end else if(N1149) begin
      btb_q[2062] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2061] <= 1'b0;
    end else if(N1149) begin
      btb_q[2061] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2060] <= 1'b0;
    end else if(N1149) begin
      btb_q[2060] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2059] <= 1'b0;
    end else if(N1149) begin
      btb_q[2059] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2058] <= 1'b0;
    end else if(N1149) begin
      btb_q[2058] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2057] <= 1'b0;
    end else if(N1149) begin
      btb_q[2057] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2056] <= 1'b0;
    end else if(N1149) begin
      btb_q[2056] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2055] <= 1'b0;
    end else if(N1149) begin
      btb_q[2055] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2054] <= 1'b0;
    end else if(N1149) begin
      btb_q[2054] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2053] <= 1'b0;
    end else if(N1149) begin
      btb_q[2053] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2052] <= 1'b0;
    end else if(N1149) begin
      btb_q[2052] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2051] <= 1'b0;
    end else if(N1149) begin
      btb_q[2051] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2050] <= 1'b0;
    end else if(N1149) begin
      btb_q[2050] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2049] <= 1'b0;
    end else if(N1149) begin
      btb_q[2049] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2048] <= 1'b0;
    end else if(N1149) begin
      btb_q[2048] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2047] <= 1'b0;
    end else if(N1150) begin
      btb_q[2047] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2046] <= 1'b0;
    end else if(N1150) begin
      btb_q[2046] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2045] <= 1'b0;
    end else if(N1150) begin
      btb_q[2045] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2044] <= 1'b0;
    end else if(N1150) begin
      btb_q[2044] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2043] <= 1'b0;
    end else if(N1150) begin
      btb_q[2043] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2042] <= 1'b0;
    end else if(N1150) begin
      btb_q[2042] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2041] <= 1'b0;
    end else if(N1150) begin
      btb_q[2041] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2040] <= 1'b0;
    end else if(N1150) begin
      btb_q[2040] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2039] <= 1'b0;
    end else if(N1150) begin
      btb_q[2039] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2038] <= 1'b0;
    end else if(N1150) begin
      btb_q[2038] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2037] <= 1'b0;
    end else if(N1150) begin
      btb_q[2037] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2036] <= 1'b0;
    end else if(N1150) begin
      btb_q[2036] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2035] <= 1'b0;
    end else if(N1150) begin
      btb_q[2035] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2034] <= 1'b0;
    end else if(N1150) begin
      btb_q[2034] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2033] <= 1'b0;
    end else if(N1150) begin
      btb_q[2033] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2032] <= 1'b0;
    end else if(N1150) begin
      btb_q[2032] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2031] <= 1'b0;
    end else if(N1150) begin
      btb_q[2031] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2030] <= 1'b0;
    end else if(N1150) begin
      btb_q[2030] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2029] <= 1'b0;
    end else if(N1150) begin
      btb_q[2029] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2028] <= 1'b0;
    end else if(N1150) begin
      btb_q[2028] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2027] <= 1'b0;
    end else if(N1150) begin
      btb_q[2027] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2026] <= 1'b0;
    end else if(N1150) begin
      btb_q[2026] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2025] <= 1'b0;
    end else if(N1150) begin
      btb_q[2025] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2024] <= 1'b0;
    end else if(N1150) begin
      btb_q[2024] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2023] <= 1'b0;
    end else if(N1150) begin
      btb_q[2023] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2022] <= 1'b0;
    end else if(N1150) begin
      btb_q[2022] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2021] <= 1'b0;
    end else if(N1150) begin
      btb_q[2021] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2020] <= 1'b0;
    end else if(N1150) begin
      btb_q[2020] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2019] <= 1'b0;
    end else if(N1150) begin
      btb_q[2019] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2018] <= 1'b0;
    end else if(N1150) begin
      btb_q[2018] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2017] <= 1'b0;
    end else if(N1150) begin
      btb_q[2017] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2016] <= 1'b0;
    end else if(N1150) begin
      btb_q[2016] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2015] <= 1'b0;
    end else if(N1150) begin
      btb_q[2015] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2014] <= 1'b0;
    end else if(N1151) begin
      btb_q[2014] <= N560;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2013] <= 1'b0;
    end else if(N1155) begin
      btb_q[2013] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2012] <= 1'b0;
    end else if(N1155) begin
      btb_q[2012] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2011] <= 1'b0;
    end else if(N1155) begin
      btb_q[2011] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2010] <= 1'b0;
    end else if(N1155) begin
      btb_q[2010] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2009] <= 1'b0;
    end else if(N1159) begin
      btb_q[2009] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2008] <= 1'b0;
    end else if(N1159) begin
      btb_q[2008] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2007] <= 1'b0;
    end else if(N1159) begin
      btb_q[2007] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2006] <= 1'b0;
    end else if(N1159) begin
      btb_q[2006] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2005] <= 1'b0;
    end else if(N1159) begin
      btb_q[2005] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2004] <= 1'b0;
    end else if(N1159) begin
      btb_q[2004] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2003] <= 1'b0;
    end else if(N1159) begin
      btb_q[2003] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2002] <= 1'b0;
    end else if(N1159) begin
      btb_q[2002] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2001] <= 1'b0;
    end else if(N1159) begin
      btb_q[2001] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2000] <= 1'b0;
    end else if(N1159) begin
      btb_q[2000] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1999] <= 1'b0;
    end else if(N1159) begin
      btb_q[1999] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1998] <= 1'b0;
    end else if(N1159) begin
      btb_q[1998] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1997] <= 1'b0;
    end else if(N1159) begin
      btb_q[1997] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1996] <= 1'b0;
    end else if(N1159) begin
      btb_q[1996] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1995] <= 1'b0;
    end else if(N1159) begin
      btb_q[1995] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1994] <= 1'b0;
    end else if(N1159) begin
      btb_q[1994] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1993] <= 1'b0;
    end else if(N1159) begin
      btb_q[1993] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1992] <= 1'b0;
    end else if(N1159) begin
      btb_q[1992] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1991] <= 1'b0;
    end else if(N1159) begin
      btb_q[1991] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1990] <= 1'b0;
    end else if(N1159) begin
      btb_q[1990] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1989] <= 1'b0;
    end else if(N1159) begin
      btb_q[1989] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1988] <= 1'b0;
    end else if(N1159) begin
      btb_q[1988] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1987] <= 1'b0;
    end else if(N1159) begin
      btb_q[1987] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1986] <= 1'b0;
    end else if(N1159) begin
      btb_q[1986] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1985] <= 1'b0;
    end else if(N1159) begin
      btb_q[1985] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1984] <= 1'b0;
    end else if(N1159) begin
      btb_q[1984] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1983] <= 1'b0;
    end else if(N1159) begin
      btb_q[1983] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1982] <= 1'b0;
    end else if(N1159) begin
      btb_q[1982] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1981] <= 1'b0;
    end else if(N1159) begin
      btb_q[1981] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1980] <= 1'b0;
    end else if(N1159) begin
      btb_q[1980] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1979] <= 1'b0;
    end else if(N1162) begin
      btb_q[1979] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1978] <= 1'b0;
    end else if(N1162) begin
      btb_q[1978] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1977] <= 1'b0;
    end else if(N1162) begin
      btb_q[1977] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1976] <= 1'b0;
    end else if(N1162) begin
      btb_q[1976] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1975] <= 1'b0;
    end else if(N1162) begin
      btb_q[1975] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1974] <= 1'b0;
    end else if(N1162) begin
      btb_q[1974] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1973] <= 1'b0;
    end else if(N1162) begin
      btb_q[1973] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1972] <= 1'b0;
    end else if(N1162) begin
      btb_q[1972] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1971] <= 1'b0;
    end else if(N1162) begin
      btb_q[1971] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1970] <= 1'b0;
    end else if(N1162) begin
      btb_q[1970] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1969] <= 1'b0;
    end else if(N1162) begin
      btb_q[1969] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1968] <= 1'b0;
    end else if(N1162) begin
      btb_q[1968] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1967] <= 1'b0;
    end else if(N1162) begin
      btb_q[1967] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1966] <= 1'b0;
    end else if(N1162) begin
      btb_q[1966] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1965] <= 1'b0;
    end else if(N1162) begin
      btb_q[1965] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1964] <= 1'b0;
    end else if(N1162) begin
      btb_q[1964] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1963] <= 1'b0;
    end else if(N1162) begin
      btb_q[1963] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1962] <= 1'b0;
    end else if(N1162) begin
      btb_q[1962] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1961] <= 1'b0;
    end else if(N1162) begin
      btb_q[1961] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1960] <= 1'b0;
    end else if(N1162) begin
      btb_q[1960] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1959] <= 1'b0;
    end else if(N1162) begin
      btb_q[1959] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1958] <= 1'b0;
    end else if(N1162) begin
      btb_q[1958] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1957] <= 1'b0;
    end else if(N1162) begin
      btb_q[1957] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1956] <= 1'b0;
    end else if(N1162) begin
      btb_q[1956] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1955] <= 1'b0;
    end else if(N1162) begin
      btb_q[1955] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1954] <= 1'b0;
    end else if(N1162) begin
      btb_q[1954] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1953] <= 1'b0;
    end else if(N1162) begin
      btb_q[1953] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1952] <= 1'b0;
    end else if(N1162) begin
      btb_q[1952] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1951] <= 1'b0;
    end else if(N1162) begin
      btb_q[1951] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1950] <= 1'b0;
    end else if(N1162) begin
      btb_q[1950] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1949] <= 1'b0;
    end else if(N1163) begin
      btb_q[1949] <= N559;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1948] <= 1'b0;
    end else if(N1167) begin
      btb_q[1948] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1947] <= 1'b0;
    end else if(N1167) begin
      btb_q[1947] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1946] <= 1'b0;
    end else if(N1168) begin
      btb_q[1946] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1945] <= 1'b0;
    end else if(N1168) begin
      btb_q[1945] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1944] <= 1'b0;
    end else if(N1168) begin
      btb_q[1944] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1943] <= 1'b0;
    end else if(N1168) begin
      btb_q[1943] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1942] <= 1'b0;
    end else if(N1168) begin
      btb_q[1942] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1941] <= 1'b0;
    end else if(N1168) begin
      btb_q[1941] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1940] <= 1'b0;
    end else if(N1168) begin
      btb_q[1940] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1939] <= 1'b0;
    end else if(N1168) begin
      btb_q[1939] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1938] <= 1'b0;
    end else if(N1168) begin
      btb_q[1938] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1937] <= 1'b0;
    end else if(N1168) begin
      btb_q[1937] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1936] <= 1'b0;
    end else if(N1168) begin
      btb_q[1936] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1935] <= 1'b0;
    end else if(N1168) begin
      btb_q[1935] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1934] <= 1'b0;
    end else if(N1168) begin
      btb_q[1934] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1933] <= 1'b0;
    end else if(N1168) begin
      btb_q[1933] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1932] <= 1'b0;
    end else if(N1168) begin
      btb_q[1932] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1931] <= 1'b0;
    end else if(N1168) begin
      btb_q[1931] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1930] <= 1'b0;
    end else if(N1168) begin
      btb_q[1930] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1929] <= 1'b0;
    end else if(N1168) begin
      btb_q[1929] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1928] <= 1'b0;
    end else if(N1168) begin
      btb_q[1928] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1927] <= 1'b0;
    end else if(N1168) begin
      btb_q[1927] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1926] <= 1'b0;
    end else if(N1168) begin
      btb_q[1926] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1925] <= 1'b0;
    end else if(N1168) begin
      btb_q[1925] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1924] <= 1'b0;
    end else if(N1168) begin
      btb_q[1924] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1923] <= 1'b0;
    end else if(N1168) begin
      btb_q[1923] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1922] <= 1'b0;
    end else if(N1168) begin
      btb_q[1922] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1921] <= 1'b0;
    end else if(N1168) begin
      btb_q[1921] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1920] <= 1'b0;
    end else if(N1168) begin
      btb_q[1920] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1919] <= 1'b0;
    end else if(N1168) begin
      btb_q[1919] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1918] <= 1'b0;
    end else if(N1168) begin
      btb_q[1918] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1917] <= 1'b0;
    end else if(N1168) begin
      btb_q[1917] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1916] <= 1'b0;
    end else if(N1168) begin
      btb_q[1916] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1915] <= 1'b0;
    end else if(N1168) begin
      btb_q[1915] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1914] <= 1'b0;
    end else if(N1168) begin
      btb_q[1914] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1913] <= 1'b0;
    end else if(N1168) begin
      btb_q[1913] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1912] <= 1'b0;
    end else if(N1168) begin
      btb_q[1912] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1911] <= 1'b0;
    end else if(N1168) begin
      btb_q[1911] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1910] <= 1'b0;
    end else if(N1168) begin
      btb_q[1910] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1909] <= 1'b0;
    end else if(N1172) begin
      btb_q[1909] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1908] <= 1'b0;
    end else if(N1172) begin
      btb_q[1908] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1907] <= 1'b0;
    end else if(N1172) begin
      btb_q[1907] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1906] <= 1'b0;
    end else if(N1172) begin
      btb_q[1906] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1905] <= 1'b0;
    end else if(N1172) begin
      btb_q[1905] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1904] <= 1'b0;
    end else if(N1172) begin
      btb_q[1904] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1903] <= 1'b0;
    end else if(N1172) begin
      btb_q[1903] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1902] <= 1'b0;
    end else if(N1172) begin
      btb_q[1902] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1901] <= 1'b0;
    end else if(N1172) begin
      btb_q[1901] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1900] <= 1'b0;
    end else if(N1172) begin
      btb_q[1900] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1899] <= 1'b0;
    end else if(N1172) begin
      btb_q[1899] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1898] <= 1'b0;
    end else if(N1172) begin
      btb_q[1898] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1897] <= 1'b0;
    end else if(N1172) begin
      btb_q[1897] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1896] <= 1'b0;
    end else if(N1172) begin
      btb_q[1896] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1895] <= 1'b0;
    end else if(N1172) begin
      btb_q[1895] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1894] <= 1'b0;
    end else if(N1172) begin
      btb_q[1894] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1893] <= 1'b0;
    end else if(N1172) begin
      btb_q[1893] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1892] <= 1'b0;
    end else if(N1172) begin
      btb_q[1892] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1891] <= 1'b0;
    end else if(N1172) begin
      btb_q[1891] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1890] <= 1'b0;
    end else if(N1172) begin
      btb_q[1890] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1889] <= 1'b0;
    end else if(N1172) begin
      btb_q[1889] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1888] <= 1'b0;
    end else if(N1172) begin
      btb_q[1888] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1887] <= 1'b0;
    end else if(N1172) begin
      btb_q[1887] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1886] <= 1'b0;
    end else if(N1172) begin
      btb_q[1886] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1885] <= 1'b0;
    end else if(N1172) begin
      btb_q[1885] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1884] <= 1'b0;
    end else if(N1163) begin
      btb_q[1884] <= N558;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1883] <= 1'b0;
    end else if(N1176) begin
      btb_q[1883] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1882] <= 1'b0;
    end else if(N1176) begin
      btb_q[1882] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1881] <= 1'b0;
    end else if(N1176) begin
      btb_q[1881] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1880] <= 1'b0;
    end else if(N1179) begin
      btb_q[1880] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1879] <= 1'b0;
    end else if(N1179) begin
      btb_q[1879] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1878] <= 1'b0;
    end else if(N1179) begin
      btb_q[1878] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1877] <= 1'b0;
    end else if(N1179) begin
      btb_q[1877] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1876] <= 1'b0;
    end else if(N1179) begin
      btb_q[1876] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1875] <= 1'b0;
    end else if(N1179) begin
      btb_q[1875] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1874] <= 1'b0;
    end else if(N1179) begin
      btb_q[1874] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1873] <= 1'b0;
    end else if(N1179) begin
      btb_q[1873] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1872] <= 1'b0;
    end else if(N1179) begin
      btb_q[1872] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1871] <= 1'b0;
    end else if(N1179) begin
      btb_q[1871] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1870] <= 1'b0;
    end else if(N1179) begin
      btb_q[1870] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1869] <= 1'b0;
    end else if(N1179) begin
      btb_q[1869] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1868] <= 1'b0;
    end else if(N1179) begin
      btb_q[1868] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1867] <= 1'b0;
    end else if(N1179) begin
      btb_q[1867] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1866] <= 1'b0;
    end else if(N1179) begin
      btb_q[1866] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1865] <= 1'b0;
    end else if(N1179) begin
      btb_q[1865] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1864] <= 1'b0;
    end else if(N1179) begin
      btb_q[1864] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1863] <= 1'b0;
    end else if(N1179) begin
      btb_q[1863] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1862] <= 1'b0;
    end else if(N1179) begin
      btb_q[1862] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1861] <= 1'b0;
    end else if(N1179) begin
      btb_q[1861] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1860] <= 1'b0;
    end else if(N1179) begin
      btb_q[1860] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1859] <= 1'b0;
    end else if(N1179) begin
      btb_q[1859] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1858] <= 1'b0;
    end else if(N1179) begin
      btb_q[1858] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1857] <= 1'b0;
    end else if(N1179) begin
      btb_q[1857] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1856] <= 1'b0;
    end else if(N1179) begin
      btb_q[1856] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1855] <= 1'b0;
    end else if(N1179) begin
      btb_q[1855] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1854] <= 1'b0;
    end else if(N1179) begin
      btb_q[1854] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1853] <= 1'b0;
    end else if(N1179) begin
      btb_q[1853] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1852] <= 1'b0;
    end else if(N1179) begin
      btb_q[1852] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1851] <= 1'b0;
    end else if(N1179) begin
      btb_q[1851] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1850] <= 1'b0;
    end else if(N1179) begin
      btb_q[1850] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1849] <= 1'b0;
    end else if(N1179) begin
      btb_q[1849] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1848] <= 1'b0;
    end else if(N1179) begin
      btb_q[1848] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1847] <= 1'b0;
    end else if(N1179) begin
      btb_q[1847] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1846] <= 1'b0;
    end else if(N1180) begin
      btb_q[1846] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1845] <= 1'b0;
    end else if(N1180) begin
      btb_q[1845] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1844] <= 1'b0;
    end else if(N1180) begin
      btb_q[1844] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1843] <= 1'b0;
    end else if(N1180) begin
      btb_q[1843] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1842] <= 1'b0;
    end else if(N1180) begin
      btb_q[1842] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1841] <= 1'b0;
    end else if(N1180) begin
      btb_q[1841] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1840] <= 1'b0;
    end else if(N1180) begin
      btb_q[1840] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1839] <= 1'b0;
    end else if(N1180) begin
      btb_q[1839] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1838] <= 1'b0;
    end else if(N1180) begin
      btb_q[1838] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1837] <= 1'b0;
    end else if(N1180) begin
      btb_q[1837] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1836] <= 1'b0;
    end else if(N1180) begin
      btb_q[1836] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1835] <= 1'b0;
    end else if(N1180) begin
      btb_q[1835] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1834] <= 1'b0;
    end else if(N1180) begin
      btb_q[1834] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1833] <= 1'b0;
    end else if(N1180) begin
      btb_q[1833] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1832] <= 1'b0;
    end else if(N1180) begin
      btb_q[1832] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1831] <= 1'b0;
    end else if(N1180) begin
      btb_q[1831] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1830] <= 1'b0;
    end else if(N1180) begin
      btb_q[1830] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1829] <= 1'b0;
    end else if(N1180) begin
      btb_q[1829] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1828] <= 1'b0;
    end else if(N1180) begin
      btb_q[1828] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1827] <= 1'b0;
    end else if(N1180) begin
      btb_q[1827] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1826] <= 1'b0;
    end else if(N1180) begin
      btb_q[1826] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1825] <= 1'b0;
    end else if(N1180) begin
      btb_q[1825] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1824] <= 1'b0;
    end else if(N1180) begin
      btb_q[1824] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1823] <= 1'b0;
    end else if(N1180) begin
      btb_q[1823] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1822] <= 1'b0;
    end else if(N1180) begin
      btb_q[1822] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1821] <= 1'b0;
    end else if(N1180) begin
      btb_q[1821] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1820] <= 1'b0;
    end else if(N1180) begin
      btb_q[1820] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1819] <= 1'b0;
    end else if(N1181) begin
      btb_q[1819] <= N557;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1818] <= 1'b0;
    end else if(N1185) begin
      btb_q[1818] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1817] <= 1'b0;
    end else if(N1185) begin
      btb_q[1817] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1816] <= 1'b0;
    end else if(N1185) begin
      btb_q[1816] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1815] <= 1'b0;
    end else if(N1185) begin
      btb_q[1815] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1814] <= 1'b0;
    end else if(N1185) begin
      btb_q[1814] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1813] <= 1'b0;
    end else if(N1185) begin
      btb_q[1813] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1812] <= 1'b0;
    end else if(N1185) begin
      btb_q[1812] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1811] <= 1'b0;
    end else if(N1185) begin
      btb_q[1811] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1810] <= 1'b0;
    end else if(N1185) begin
      btb_q[1810] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1809] <= 1'b0;
    end else if(N1185) begin
      btb_q[1809] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1808] <= 1'b0;
    end else if(N1189) begin
      btb_q[1808] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1807] <= 1'b0;
    end else if(N1189) begin
      btb_q[1807] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1806] <= 1'b0;
    end else if(N1189) begin
      btb_q[1806] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1805] <= 1'b0;
    end else if(N1189) begin
      btb_q[1805] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1804] <= 1'b0;
    end else if(N1189) begin
      btb_q[1804] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1803] <= 1'b0;
    end else if(N1189) begin
      btb_q[1803] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1802] <= 1'b0;
    end else if(N1189) begin
      btb_q[1802] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1801] <= 1'b0;
    end else if(N1189) begin
      btb_q[1801] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1800] <= 1'b0;
    end else if(N1189) begin
      btb_q[1800] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1799] <= 1'b0;
    end else if(N1189) begin
      btb_q[1799] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1798] <= 1'b0;
    end else if(N1189) begin
      btb_q[1798] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1797] <= 1'b0;
    end else if(N1189) begin
      btb_q[1797] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1796] <= 1'b0;
    end else if(N1189) begin
      btb_q[1796] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1795] <= 1'b0;
    end else if(N1189) begin
      btb_q[1795] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1794] <= 1'b0;
    end else if(N1189) begin
      btb_q[1794] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1793] <= 1'b0;
    end else if(N1189) begin
      btb_q[1793] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1792] <= 1'b0;
    end else if(N1189) begin
      btb_q[1792] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1791] <= 1'b0;
    end else if(N1189) begin
      btb_q[1791] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1790] <= 1'b0;
    end else if(N1189) begin
      btb_q[1790] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1789] <= 1'b0;
    end else if(N1189) begin
      btb_q[1789] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1788] <= 1'b0;
    end else if(N1189) begin
      btb_q[1788] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1787] <= 1'b0;
    end else if(N1189) begin
      btb_q[1787] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1786] <= 1'b0;
    end else if(N1189) begin
      btb_q[1786] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1785] <= 1'b0;
    end else if(N1189) begin
      btb_q[1785] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1784] <= 1'b0;
    end else if(N1189) begin
      btb_q[1784] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1783] <= 1'b0;
    end else if(N1189) begin
      btb_q[1783] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1782] <= 1'b0;
    end else if(N1189) begin
      btb_q[1782] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1781] <= 1'b0;
    end else if(N1192) begin
      btb_q[1781] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1780] <= 1'b0;
    end else if(N1192) begin
      btb_q[1780] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1779] <= 1'b0;
    end else if(N1192) begin
      btb_q[1779] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1778] <= 1'b0;
    end else if(N1192) begin
      btb_q[1778] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1777] <= 1'b0;
    end else if(N1192) begin
      btb_q[1777] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1776] <= 1'b0;
    end else if(N1192) begin
      btb_q[1776] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1775] <= 1'b0;
    end else if(N1192) begin
      btb_q[1775] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1774] <= 1'b0;
    end else if(N1192) begin
      btb_q[1774] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1773] <= 1'b0;
    end else if(N1192) begin
      btb_q[1773] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1772] <= 1'b0;
    end else if(N1192) begin
      btb_q[1772] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1771] <= 1'b0;
    end else if(N1192) begin
      btb_q[1771] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1770] <= 1'b0;
    end else if(N1192) begin
      btb_q[1770] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1769] <= 1'b0;
    end else if(N1192) begin
      btb_q[1769] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1768] <= 1'b0;
    end else if(N1192) begin
      btb_q[1768] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1767] <= 1'b0;
    end else if(N1192) begin
      btb_q[1767] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1766] <= 1'b0;
    end else if(N1192) begin
      btb_q[1766] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1765] <= 1'b0;
    end else if(N1192) begin
      btb_q[1765] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1764] <= 1'b0;
    end else if(N1192) begin
      btb_q[1764] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1763] <= 1'b0;
    end else if(N1192) begin
      btb_q[1763] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1762] <= 1'b0;
    end else if(N1192) begin
      btb_q[1762] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1761] <= 1'b0;
    end else if(N1192) begin
      btb_q[1761] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1760] <= 1'b0;
    end else if(N1192) begin
      btb_q[1760] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1759] <= 1'b0;
    end else if(N1192) begin
      btb_q[1759] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1758] <= 1'b0;
    end else if(N1192) begin
      btb_q[1758] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1757] <= 1'b0;
    end else if(N1192) begin
      btb_q[1757] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1756] <= 1'b0;
    end else if(N1192) begin
      btb_q[1756] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1755] <= 1'b0;
    end else if(N1192) begin
      btb_q[1755] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1754] <= 1'b0;
    end else if(N1193) begin
      btb_q[1754] <= N556;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1753] <= 1'b0;
    end else if(N1197) begin
      btb_q[1753] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1752] <= 1'b0;
    end else if(N1197) begin
      btb_q[1752] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1751] <= 1'b0;
    end else if(N1197) begin
      btb_q[1751] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1750] <= 1'b0;
    end else if(N1197) begin
      btb_q[1750] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1749] <= 1'b0;
    end else if(N1197) begin
      btb_q[1749] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1748] <= 1'b0;
    end else if(N1197) begin
      btb_q[1748] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1747] <= 1'b0;
    end else if(N1197) begin
      btb_q[1747] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1746] <= 1'b0;
    end else if(N1197) begin
      btb_q[1746] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1745] <= 1'b0;
    end else if(N1198) begin
      btb_q[1745] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1744] <= 1'b0;
    end else if(N1198) begin
      btb_q[1744] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1743] <= 1'b0;
    end else if(N1198) begin
      btb_q[1743] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1742] <= 1'b0;
    end else if(N1198) begin
      btb_q[1742] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1741] <= 1'b0;
    end else if(N1198) begin
      btb_q[1741] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1740] <= 1'b0;
    end else if(N1198) begin
      btb_q[1740] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1739] <= 1'b0;
    end else if(N1198) begin
      btb_q[1739] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1738] <= 1'b0;
    end else if(N1198) begin
      btb_q[1738] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1737] <= 1'b0;
    end else if(N1198) begin
      btb_q[1737] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1736] <= 1'b0;
    end else if(N1198) begin
      btb_q[1736] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1735] <= 1'b0;
    end else if(N1198) begin
      btb_q[1735] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1734] <= 1'b0;
    end else if(N1198) begin
      btb_q[1734] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1733] <= 1'b0;
    end else if(N1198) begin
      btb_q[1733] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1732] <= 1'b0;
    end else if(N1198) begin
      btb_q[1732] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1731] <= 1'b0;
    end else if(N1198) begin
      btb_q[1731] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1730] <= 1'b0;
    end else if(N1198) begin
      btb_q[1730] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1729] <= 1'b0;
    end else if(N1198) begin
      btb_q[1729] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1728] <= 1'b0;
    end else if(N1198) begin
      btb_q[1728] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1727] <= 1'b0;
    end else if(N1198) begin
      btb_q[1727] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1726] <= 1'b0;
    end else if(N1198) begin
      btb_q[1726] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1725] <= 1'b0;
    end else if(N1198) begin
      btb_q[1725] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1724] <= 1'b0;
    end else if(N1198) begin
      btb_q[1724] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1723] <= 1'b0;
    end else if(N1198) begin
      btb_q[1723] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1722] <= 1'b0;
    end else if(N1198) begin
      btb_q[1722] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1721] <= 1'b0;
    end else if(N1198) begin
      btb_q[1721] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1720] <= 1'b0;
    end else if(N1198) begin
      btb_q[1720] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1719] <= 1'b0;
    end else if(N1198) begin
      btb_q[1719] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1718] <= 1'b0;
    end else if(N1198) begin
      btb_q[1718] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1717] <= 1'b0;
    end else if(N1198) begin
      btb_q[1717] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1716] <= 1'b0;
    end else if(N1198) begin
      btb_q[1716] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1715] <= 1'b0;
    end else if(N1198) begin
      btb_q[1715] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1714] <= 1'b0;
    end else if(N1198) begin
      btb_q[1714] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1713] <= 1'b0;
    end else if(N1198) begin
      btb_q[1713] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1712] <= 1'b0;
    end else if(N1198) begin
      btb_q[1712] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1711] <= 1'b0;
    end else if(N1198) begin
      btb_q[1711] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1710] <= 1'b0;
    end else if(N1198) begin
      btb_q[1710] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1709] <= 1'b0;
    end else if(N1198) begin
      btb_q[1709] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1708] <= 1'b0;
    end else if(N1202) begin
      btb_q[1708] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1707] <= 1'b0;
    end else if(N1202) begin
      btb_q[1707] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1706] <= 1'b0;
    end else if(N1202) begin
      btb_q[1706] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1705] <= 1'b0;
    end else if(N1202) begin
      btb_q[1705] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1704] <= 1'b0;
    end else if(N1202) begin
      btb_q[1704] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1703] <= 1'b0;
    end else if(N1202) begin
      btb_q[1703] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1702] <= 1'b0;
    end else if(N1202) begin
      btb_q[1702] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1701] <= 1'b0;
    end else if(N1202) begin
      btb_q[1701] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1700] <= 1'b0;
    end else if(N1202) begin
      btb_q[1700] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1699] <= 1'b0;
    end else if(N1202) begin
      btb_q[1699] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1698] <= 1'b0;
    end else if(N1202) begin
      btb_q[1698] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1697] <= 1'b0;
    end else if(N1202) begin
      btb_q[1697] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1696] <= 1'b0;
    end else if(N1202) begin
      btb_q[1696] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1695] <= 1'b0;
    end else if(N1202) begin
      btb_q[1695] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1694] <= 1'b0;
    end else if(N1202) begin
      btb_q[1694] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1693] <= 1'b0;
    end else if(N1202) begin
      btb_q[1693] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1692] <= 1'b0;
    end else if(N1202) begin
      btb_q[1692] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1691] <= 1'b0;
    end else if(N1202) begin
      btb_q[1691] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1690] <= 1'b0;
    end else if(N1202) begin
      btb_q[1690] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1689] <= 1'b0;
    end else if(N1193) begin
      btb_q[1689] <= N555;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1688] <= 1'b0;
    end else if(N1206) begin
      btb_q[1688] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1687] <= 1'b0;
    end else if(N1206) begin
      btb_q[1687] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1686] <= 1'b0;
    end else if(N1206) begin
      btb_q[1686] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1685] <= 1'b0;
    end else if(N1206) begin
      btb_q[1685] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1684] <= 1'b0;
    end else if(N1206) begin
      btb_q[1684] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1683] <= 1'b0;
    end else if(N1206) begin
      btb_q[1683] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1682] <= 1'b0;
    end else if(N1209) begin
      btb_q[1682] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1681] <= 1'b0;
    end else if(N1209) begin
      btb_q[1681] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1680] <= 1'b0;
    end else if(N1209) begin
      btb_q[1680] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1679] <= 1'b0;
    end else if(N1209) begin
      btb_q[1679] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1678] <= 1'b0;
    end else if(N1209) begin
      btb_q[1678] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1677] <= 1'b0;
    end else if(N1209) begin
      btb_q[1677] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1676] <= 1'b0;
    end else if(N1209) begin
      btb_q[1676] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1675] <= 1'b0;
    end else if(N1209) begin
      btb_q[1675] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1674] <= 1'b0;
    end else if(N1209) begin
      btb_q[1674] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1673] <= 1'b0;
    end else if(N1209) begin
      btb_q[1673] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1672] <= 1'b0;
    end else if(N1209) begin
      btb_q[1672] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1671] <= 1'b0;
    end else if(N1209) begin
      btb_q[1671] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1670] <= 1'b0;
    end else if(N1209) begin
      btb_q[1670] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1669] <= 1'b0;
    end else if(N1209) begin
      btb_q[1669] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1668] <= 1'b0;
    end else if(N1209) begin
      btb_q[1668] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1667] <= 1'b0;
    end else if(N1209) begin
      btb_q[1667] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1666] <= 1'b0;
    end else if(N1209) begin
      btb_q[1666] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1665] <= 1'b0;
    end else if(N1209) begin
      btb_q[1665] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1664] <= 1'b0;
    end else if(N1209) begin
      btb_q[1664] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1663] <= 1'b0;
    end else if(N1209) begin
      btb_q[1663] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1662] <= 1'b0;
    end else if(N1209) begin
      btb_q[1662] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1661] <= 1'b0;
    end else if(N1209) begin
      btb_q[1661] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1660] <= 1'b0;
    end else if(N1209) begin
      btb_q[1660] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1659] <= 1'b0;
    end else if(N1209) begin
      btb_q[1659] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1658] <= 1'b0;
    end else if(N1209) begin
      btb_q[1658] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1657] <= 1'b0;
    end else if(N1209) begin
      btb_q[1657] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1656] <= 1'b0;
    end else if(N1209) begin
      btb_q[1656] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1655] <= 1'b0;
    end else if(N1209) begin
      btb_q[1655] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1654] <= 1'b0;
    end else if(N1209) begin
      btb_q[1654] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1653] <= 1'b0;
    end else if(N1209) begin
      btb_q[1653] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1652] <= 1'b0;
    end else if(N1209) begin
      btb_q[1652] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1651] <= 1'b0;
    end else if(N1209) begin
      btb_q[1651] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1650] <= 1'b0;
    end else if(N1209) begin
      btb_q[1650] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1649] <= 1'b0;
    end else if(N1209) begin
      btb_q[1649] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1648] <= 1'b0;
    end else if(N1209) begin
      btb_q[1648] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1647] <= 1'b0;
    end else if(N1209) begin
      btb_q[1647] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1646] <= 1'b0;
    end else if(N1209) begin
      btb_q[1646] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1645] <= 1'b0;
    end else if(N1210) begin
      btb_q[1645] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1644] <= 1'b0;
    end else if(N1210) begin
      btb_q[1644] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1643] <= 1'b0;
    end else if(N1210) begin
      btb_q[1643] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1642] <= 1'b0;
    end else if(N1210) begin
      btb_q[1642] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1641] <= 1'b0;
    end else if(N1210) begin
      btb_q[1641] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1640] <= 1'b0;
    end else if(N1210) begin
      btb_q[1640] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1639] <= 1'b0;
    end else if(N1210) begin
      btb_q[1639] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1638] <= 1'b0;
    end else if(N1210) begin
      btb_q[1638] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1637] <= 1'b0;
    end else if(N1210) begin
      btb_q[1637] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1636] <= 1'b0;
    end else if(N1210) begin
      btb_q[1636] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1635] <= 1'b0;
    end else if(N1210) begin
      btb_q[1635] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1634] <= 1'b0;
    end else if(N1210) begin
      btb_q[1634] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1633] <= 1'b0;
    end else if(N1210) begin
      btb_q[1633] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1632] <= 1'b0;
    end else if(N1210) begin
      btb_q[1632] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1631] <= 1'b0;
    end else if(N1210) begin
      btb_q[1631] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1630] <= 1'b0;
    end else if(N1210) begin
      btb_q[1630] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1629] <= 1'b0;
    end else if(N1210) begin
      btb_q[1629] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1628] <= 1'b0;
    end else if(N1210) begin
      btb_q[1628] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1627] <= 1'b0;
    end else if(N1210) begin
      btb_q[1627] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1626] <= 1'b0;
    end else if(N1210) begin
      btb_q[1626] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1625] <= 1'b0;
    end else if(N1210) begin
      btb_q[1625] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1624] <= 1'b0;
    end else if(N1211) begin
      btb_q[1624] <= N554;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1623] <= 1'b0;
    end else if(N1215) begin
      btb_q[1623] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1622] <= 1'b0;
    end else if(N1215) begin
      btb_q[1622] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1621] <= 1'b0;
    end else if(N1215) begin
      btb_q[1621] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1620] <= 1'b0;
    end else if(N1215) begin
      btb_q[1620] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1619] <= 1'b0;
    end else if(N1215) begin
      btb_q[1619] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1618] <= 1'b0;
    end else if(N1215) begin
      btb_q[1618] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1617] <= 1'b0;
    end else if(N1215) begin
      btb_q[1617] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1616] <= 1'b0;
    end else if(N1215) begin
      btb_q[1616] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1615] <= 1'b0;
    end else if(N1215) begin
      btb_q[1615] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1614] <= 1'b0;
    end else if(N1215) begin
      btb_q[1614] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1613] <= 1'b0;
    end else if(N1215) begin
      btb_q[1613] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1612] <= 1'b0;
    end else if(N1215) begin
      btb_q[1612] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1611] <= 1'b0;
    end else if(N1215) begin
      btb_q[1611] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1610] <= 1'b0;
    end else if(N1215) begin
      btb_q[1610] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1609] <= 1'b0;
    end else if(N1215) begin
      btb_q[1609] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1608] <= 1'b0;
    end else if(N1215) begin
      btb_q[1608] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1607] <= 1'b0;
    end else if(N1219) begin
      btb_q[1607] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1606] <= 1'b0;
    end else if(N1219) begin
      btb_q[1606] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1605] <= 1'b0;
    end else if(N1219) begin
      btb_q[1605] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1604] <= 1'b0;
    end else if(N1219) begin
      btb_q[1604] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1603] <= 1'b0;
    end else if(N1219) begin
      btb_q[1603] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1602] <= 1'b0;
    end else if(N1219) begin
      btb_q[1602] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1601] <= 1'b0;
    end else if(N1219) begin
      btb_q[1601] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1600] <= 1'b0;
    end else if(N1219) begin
      btb_q[1600] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1599] <= 1'b0;
    end else if(N1219) begin
      btb_q[1599] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1598] <= 1'b0;
    end else if(N1219) begin
      btb_q[1598] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1597] <= 1'b0;
    end else if(N1219) begin
      btb_q[1597] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1596] <= 1'b0;
    end else if(N1219) begin
      btb_q[1596] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1595] <= 1'b0;
    end else if(N1219) begin
      btb_q[1595] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1594] <= 1'b0;
    end else if(N1219) begin
      btb_q[1594] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1593] <= 1'b0;
    end else if(N1219) begin
      btb_q[1593] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1592] <= 1'b0;
    end else if(N1219) begin
      btb_q[1592] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1591] <= 1'b0;
    end else if(N1219) begin
      btb_q[1591] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1590] <= 1'b0;
    end else if(N1219) begin
      btb_q[1590] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1589] <= 1'b0;
    end else if(N1219) begin
      btb_q[1589] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1588] <= 1'b0;
    end else if(N1219) begin
      btb_q[1588] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1587] <= 1'b0;
    end else if(N1219) begin
      btb_q[1587] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1586] <= 1'b0;
    end else if(N1219) begin
      btb_q[1586] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1585] <= 1'b0;
    end else if(N1219) begin
      btb_q[1585] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1584] <= 1'b0;
    end else if(N1219) begin
      btb_q[1584] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1583] <= 1'b0;
    end else if(N1222) begin
      btb_q[1583] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1582] <= 1'b0;
    end else if(N1222) begin
      btb_q[1582] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1581] <= 1'b0;
    end else if(N1222) begin
      btb_q[1581] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1580] <= 1'b0;
    end else if(N1222) begin
      btb_q[1580] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1579] <= 1'b0;
    end else if(N1222) begin
      btb_q[1579] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1578] <= 1'b0;
    end else if(N1222) begin
      btb_q[1578] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1577] <= 1'b0;
    end else if(N1222) begin
      btb_q[1577] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1576] <= 1'b0;
    end else if(N1222) begin
      btb_q[1576] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1575] <= 1'b0;
    end else if(N1222) begin
      btb_q[1575] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1574] <= 1'b0;
    end else if(N1222) begin
      btb_q[1574] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1573] <= 1'b0;
    end else if(N1222) begin
      btb_q[1573] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1572] <= 1'b0;
    end else if(N1222) begin
      btb_q[1572] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1571] <= 1'b0;
    end else if(N1222) begin
      btb_q[1571] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1570] <= 1'b0;
    end else if(N1222) begin
      btb_q[1570] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1569] <= 1'b0;
    end else if(N1222) begin
      btb_q[1569] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1568] <= 1'b0;
    end else if(N1222) begin
      btb_q[1568] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1567] <= 1'b0;
    end else if(N1222) begin
      btb_q[1567] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1566] <= 1'b0;
    end else if(N1222) begin
      btb_q[1566] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1565] <= 1'b0;
    end else if(N1222) begin
      btb_q[1565] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1564] <= 1'b0;
    end else if(N1222) begin
      btb_q[1564] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1563] <= 1'b0;
    end else if(N1222) begin
      btb_q[1563] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1562] <= 1'b0;
    end else if(N1222) begin
      btb_q[1562] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1561] <= 1'b0;
    end else if(N1222) begin
      btb_q[1561] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1560] <= 1'b0;
    end else if(N1222) begin
      btb_q[1560] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1559] <= 1'b0;
    end else if(N1223) begin
      btb_q[1559] <= N553;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1558] <= 1'b0;
    end else if(N1227) begin
      btb_q[1558] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1557] <= 1'b0;
    end else if(N1227) begin
      btb_q[1557] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1556] <= 1'b0;
    end else if(N1227) begin
      btb_q[1556] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1555] <= 1'b0;
    end else if(N1227) begin
      btb_q[1555] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1554] <= 1'b0;
    end else if(N1227) begin
      btb_q[1554] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1553] <= 1'b0;
    end else if(N1227) begin
      btb_q[1553] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1552] <= 1'b0;
    end else if(N1227) begin
      btb_q[1552] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1551] <= 1'b0;
    end else if(N1227) begin
      btb_q[1551] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1550] <= 1'b0;
    end else if(N1227) begin
      btb_q[1550] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1549] <= 1'b0;
    end else if(N1227) begin
      btb_q[1549] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1548] <= 1'b0;
    end else if(N1227) begin
      btb_q[1548] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1547] <= 1'b0;
    end else if(N1227) begin
      btb_q[1547] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1546] <= 1'b0;
    end else if(N1227) begin
      btb_q[1546] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1545] <= 1'b0;
    end else if(N1227) begin
      btb_q[1545] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1544] <= 1'b0;
    end else if(N1228) begin
      btb_q[1544] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1543] <= 1'b0;
    end else if(N1228) begin
      btb_q[1543] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1542] <= 1'b0;
    end else if(N1228) begin
      btb_q[1542] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1541] <= 1'b0;
    end else if(N1228) begin
      btb_q[1541] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1540] <= 1'b0;
    end else if(N1228) begin
      btb_q[1540] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1539] <= 1'b0;
    end else if(N1228) begin
      btb_q[1539] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1538] <= 1'b0;
    end else if(N1228) begin
      btb_q[1538] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1537] <= 1'b0;
    end else if(N1228) begin
      btb_q[1537] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1536] <= 1'b0;
    end else if(N1228) begin
      btb_q[1536] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1535] <= 1'b0;
    end else if(N1228) begin
      btb_q[1535] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1534] <= 1'b0;
    end else if(N1228) begin
      btb_q[1534] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1533] <= 1'b0;
    end else if(N1228) begin
      btb_q[1533] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1532] <= 1'b0;
    end else if(N1228) begin
      btb_q[1532] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1531] <= 1'b0;
    end else if(N1228) begin
      btb_q[1531] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1530] <= 1'b0;
    end else if(N1228) begin
      btb_q[1530] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1529] <= 1'b0;
    end else if(N1228) begin
      btb_q[1529] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1528] <= 1'b0;
    end else if(N1228) begin
      btb_q[1528] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1527] <= 1'b0;
    end else if(N1228) begin
      btb_q[1527] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1526] <= 1'b0;
    end else if(N1228) begin
      btb_q[1526] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1525] <= 1'b0;
    end else if(N1228) begin
      btb_q[1525] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1524] <= 1'b0;
    end else if(N1228) begin
      btb_q[1524] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1523] <= 1'b0;
    end else if(N1228) begin
      btb_q[1523] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1522] <= 1'b0;
    end else if(N1228) begin
      btb_q[1522] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1521] <= 1'b0;
    end else if(N1228) begin
      btb_q[1521] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1520] <= 1'b0;
    end else if(N1228) begin
      btb_q[1520] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1519] <= 1'b0;
    end else if(N1228) begin
      btb_q[1519] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1518] <= 1'b0;
    end else if(N1228) begin
      btb_q[1518] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1517] <= 1'b0;
    end else if(N1228) begin
      btb_q[1517] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1516] <= 1'b0;
    end else if(N1228) begin
      btb_q[1516] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1515] <= 1'b0;
    end else if(N1228) begin
      btb_q[1515] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1514] <= 1'b0;
    end else if(N1228) begin
      btb_q[1514] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1513] <= 1'b0;
    end else if(N1228) begin
      btb_q[1513] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1512] <= 1'b0;
    end else if(N1228) begin
      btb_q[1512] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1511] <= 1'b0;
    end else if(N1228) begin
      btb_q[1511] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1510] <= 1'b0;
    end else if(N1228) begin
      btb_q[1510] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1509] <= 1'b0;
    end else if(N1228) begin
      btb_q[1509] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1508] <= 1'b0;
    end else if(N1228) begin
      btb_q[1508] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1507] <= 1'b0;
    end else if(N1232) begin
      btb_q[1507] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1506] <= 1'b0;
    end else if(N1232) begin
      btb_q[1506] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1505] <= 1'b0;
    end else if(N1232) begin
      btb_q[1505] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1504] <= 1'b0;
    end else if(N1232) begin
      btb_q[1504] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1503] <= 1'b0;
    end else if(N1232) begin
      btb_q[1503] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1502] <= 1'b0;
    end else if(N1232) begin
      btb_q[1502] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1501] <= 1'b0;
    end else if(N1232) begin
      btb_q[1501] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1500] <= 1'b0;
    end else if(N1232) begin
      btb_q[1500] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1499] <= 1'b0;
    end else if(N1232) begin
      btb_q[1499] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1498] <= 1'b0;
    end else if(N1232) begin
      btb_q[1498] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1497] <= 1'b0;
    end else if(N1232) begin
      btb_q[1497] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1496] <= 1'b0;
    end else if(N1232) begin
      btb_q[1496] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1495] <= 1'b0;
    end else if(N1232) begin
      btb_q[1495] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1494] <= 1'b0;
    end else if(N1223) begin
      btb_q[1494] <= N552;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1493] <= 1'b0;
    end else if(N1236) begin
      btb_q[1493] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1492] <= 1'b0;
    end else if(N1236) begin
      btb_q[1492] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1491] <= 1'b0;
    end else if(N1236) begin
      btb_q[1491] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1490] <= 1'b0;
    end else if(N1236) begin
      btb_q[1490] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1489] <= 1'b0;
    end else if(N1236) begin
      btb_q[1489] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1488] <= 1'b0;
    end else if(N1236) begin
      btb_q[1488] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1487] <= 1'b0;
    end else if(N1236) begin
      btb_q[1487] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1486] <= 1'b0;
    end else if(N1236) begin
      btb_q[1486] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1485] <= 1'b0;
    end else if(N1236) begin
      btb_q[1485] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1484] <= 1'b0;
    end else if(N1239) begin
      btb_q[1484] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1483] <= 1'b0;
    end else if(N1239) begin
      btb_q[1483] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1482] <= 1'b0;
    end else if(N1239) begin
      btb_q[1482] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1481] <= 1'b0;
    end else if(N1239) begin
      btb_q[1481] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1480] <= 1'b0;
    end else if(N1239) begin
      btb_q[1480] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1479] <= 1'b0;
    end else if(N1239) begin
      btb_q[1479] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1478] <= 1'b0;
    end else if(N1239) begin
      btb_q[1478] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1477] <= 1'b0;
    end else if(N1239) begin
      btb_q[1477] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1476] <= 1'b0;
    end else if(N1239) begin
      btb_q[1476] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1475] <= 1'b0;
    end else if(N1239) begin
      btb_q[1475] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1474] <= 1'b0;
    end else if(N1239) begin
      btb_q[1474] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1473] <= 1'b0;
    end else if(N1239) begin
      btb_q[1473] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1472] <= 1'b0;
    end else if(N1239) begin
      btb_q[1472] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1471] <= 1'b0;
    end else if(N1239) begin
      btb_q[1471] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1470] <= 1'b0;
    end else if(N1239) begin
      btb_q[1470] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1469] <= 1'b0;
    end else if(N1239) begin
      btb_q[1469] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1468] <= 1'b0;
    end else if(N1239) begin
      btb_q[1468] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1467] <= 1'b0;
    end else if(N1239) begin
      btb_q[1467] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1466] <= 1'b0;
    end else if(N1239) begin
      btb_q[1466] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1465] <= 1'b0;
    end else if(N1239) begin
      btb_q[1465] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1464] <= 1'b0;
    end else if(N1239) begin
      btb_q[1464] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1463] <= 1'b0;
    end else if(N1239) begin
      btb_q[1463] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1462] <= 1'b0;
    end else if(N1239) begin
      btb_q[1462] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1461] <= 1'b0;
    end else if(N1239) begin
      btb_q[1461] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1460] <= 1'b0;
    end else if(N1239) begin
      btb_q[1460] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1459] <= 1'b0;
    end else if(N1239) begin
      btb_q[1459] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1458] <= 1'b0;
    end else if(N1239) begin
      btb_q[1458] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1457] <= 1'b0;
    end else if(N1239) begin
      btb_q[1457] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1456] <= 1'b0;
    end else if(N1239) begin
      btb_q[1456] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1455] <= 1'b0;
    end else if(N1239) begin
      btb_q[1455] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1454] <= 1'b0;
    end else if(N1239) begin
      btb_q[1454] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1453] <= 1'b0;
    end else if(N1239) begin
      btb_q[1453] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1452] <= 1'b0;
    end else if(N1239) begin
      btb_q[1452] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1451] <= 1'b0;
    end else if(N1239) begin
      btb_q[1451] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1450] <= 1'b0;
    end else if(N1239) begin
      btb_q[1450] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1449] <= 1'b0;
    end else if(N1239) begin
      btb_q[1449] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1448] <= 1'b0;
    end else if(N1239) begin
      btb_q[1448] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1447] <= 1'b0;
    end else if(N1239) begin
      btb_q[1447] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1446] <= 1'b0;
    end else if(N1239) begin
      btb_q[1446] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1445] <= 1'b0;
    end else if(N1239) begin
      btb_q[1445] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1444] <= 1'b0;
    end else if(N1240) begin
      btb_q[1444] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1443] <= 1'b0;
    end else if(N1240) begin
      btb_q[1443] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1442] <= 1'b0;
    end else if(N1240) begin
      btb_q[1442] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1441] <= 1'b0;
    end else if(N1240) begin
      btb_q[1441] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1440] <= 1'b0;
    end else if(N1240) begin
      btb_q[1440] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1439] <= 1'b0;
    end else if(N1240) begin
      btb_q[1439] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1438] <= 1'b0;
    end else if(N1240) begin
      btb_q[1438] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1437] <= 1'b0;
    end else if(N1240) begin
      btb_q[1437] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1436] <= 1'b0;
    end else if(N1240) begin
      btb_q[1436] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1435] <= 1'b0;
    end else if(N1240) begin
      btb_q[1435] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1434] <= 1'b0;
    end else if(N1240) begin
      btb_q[1434] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1433] <= 1'b0;
    end else if(N1240) begin
      btb_q[1433] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1432] <= 1'b0;
    end else if(N1240) begin
      btb_q[1432] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1431] <= 1'b0;
    end else if(N1240) begin
      btb_q[1431] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1430] <= 1'b0;
    end else if(N1240) begin
      btb_q[1430] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1429] <= 1'b0;
    end else if(N1241) begin
      btb_q[1429] <= N551;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1428] <= 1'b0;
    end else if(N1245) begin
      btb_q[1428] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1427] <= 1'b0;
    end else if(N1245) begin
      btb_q[1427] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1426] <= 1'b0;
    end else if(N1245) begin
      btb_q[1426] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1425] <= 1'b0;
    end else if(N1245) begin
      btb_q[1425] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1424] <= 1'b0;
    end else if(N1245) begin
      btb_q[1424] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1423] <= 1'b0;
    end else if(N1245) begin
      btb_q[1423] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1422] <= 1'b0;
    end else if(N1245) begin
      btb_q[1422] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1421] <= 1'b0;
    end else if(N1245) begin
      btb_q[1421] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1420] <= 1'b0;
    end else if(N1245) begin
      btb_q[1420] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1419] <= 1'b0;
    end else if(N1245) begin
      btb_q[1419] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1418] <= 1'b0;
    end else if(N1245) begin
      btb_q[1418] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1417] <= 1'b0;
    end else if(N1245) begin
      btb_q[1417] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1416] <= 1'b0;
    end else if(N1245) begin
      btb_q[1416] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1415] <= 1'b0;
    end else if(N1245) begin
      btb_q[1415] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1414] <= 1'b0;
    end else if(N1245) begin
      btb_q[1414] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1413] <= 1'b0;
    end else if(N1245) begin
      btb_q[1413] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1412] <= 1'b0;
    end else if(N1245) begin
      btb_q[1412] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1411] <= 1'b0;
    end else if(N1245) begin
      btb_q[1411] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1410] <= 1'b0;
    end else if(N1245) begin
      btb_q[1410] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1409] <= 1'b0;
    end else if(N1245) begin
      btb_q[1409] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1408] <= 1'b0;
    end else if(N1245) begin
      btb_q[1408] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1407] <= 1'b0;
    end else if(N1245) begin
      btb_q[1407] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1406] <= 1'b0;
    end else if(N1249) begin
      btb_q[1406] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1405] <= 1'b0;
    end else if(N1249) begin
      btb_q[1405] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1404] <= 1'b0;
    end else if(N1249) begin
      btb_q[1404] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1403] <= 1'b0;
    end else if(N1249) begin
      btb_q[1403] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1402] <= 1'b0;
    end else if(N1249) begin
      btb_q[1402] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1401] <= 1'b0;
    end else if(N1249) begin
      btb_q[1401] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1400] <= 1'b0;
    end else if(N1249) begin
      btb_q[1400] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1399] <= 1'b0;
    end else if(N1249) begin
      btb_q[1399] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1398] <= 1'b0;
    end else if(N1249) begin
      btb_q[1398] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1397] <= 1'b0;
    end else if(N1249) begin
      btb_q[1397] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1396] <= 1'b0;
    end else if(N1249) begin
      btb_q[1396] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1395] <= 1'b0;
    end else if(N1249) begin
      btb_q[1395] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1394] <= 1'b0;
    end else if(N1249) begin
      btb_q[1394] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1393] <= 1'b0;
    end else if(N1249) begin
      btb_q[1393] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1392] <= 1'b0;
    end else if(N1249) begin
      btb_q[1392] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1391] <= 1'b0;
    end else if(N1249) begin
      btb_q[1391] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1390] <= 1'b0;
    end else if(N1249) begin
      btb_q[1390] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1389] <= 1'b0;
    end else if(N1249) begin
      btb_q[1389] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1388] <= 1'b0;
    end else if(N1249) begin
      btb_q[1388] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1387] <= 1'b0;
    end else if(N1249) begin
      btb_q[1387] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1386] <= 1'b0;
    end else if(N1249) begin
      btb_q[1386] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1385] <= 1'b0;
    end else if(N1252) begin
      btb_q[1385] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1384] <= 1'b0;
    end else if(N1252) begin
      btb_q[1384] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1383] <= 1'b0;
    end else if(N1252) begin
      btb_q[1383] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1382] <= 1'b0;
    end else if(N1252) begin
      btb_q[1382] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1381] <= 1'b0;
    end else if(N1252) begin
      btb_q[1381] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1380] <= 1'b0;
    end else if(N1252) begin
      btb_q[1380] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1379] <= 1'b0;
    end else if(N1252) begin
      btb_q[1379] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1378] <= 1'b0;
    end else if(N1252) begin
      btb_q[1378] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1377] <= 1'b0;
    end else if(N1252) begin
      btb_q[1377] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1376] <= 1'b0;
    end else if(N1252) begin
      btb_q[1376] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1375] <= 1'b0;
    end else if(N1252) begin
      btb_q[1375] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1374] <= 1'b0;
    end else if(N1252) begin
      btb_q[1374] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1373] <= 1'b0;
    end else if(N1252) begin
      btb_q[1373] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1372] <= 1'b0;
    end else if(N1252) begin
      btb_q[1372] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1371] <= 1'b0;
    end else if(N1252) begin
      btb_q[1371] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1370] <= 1'b0;
    end else if(N1252) begin
      btb_q[1370] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1369] <= 1'b0;
    end else if(N1252) begin
      btb_q[1369] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1368] <= 1'b0;
    end else if(N1252) begin
      btb_q[1368] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1367] <= 1'b0;
    end else if(N1252) begin
      btb_q[1367] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1366] <= 1'b0;
    end else if(N1252) begin
      btb_q[1366] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1365] <= 1'b0;
    end else if(N1252) begin
      btb_q[1365] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1364] <= 1'b0;
    end else if(N1253) begin
      btb_q[1364] <= N550;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1363] <= 1'b0;
    end else if(N1257) begin
      btb_q[1363] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1362] <= 1'b0;
    end else if(N1257) begin
      btb_q[1362] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1361] <= 1'b0;
    end else if(N1257) begin
      btb_q[1361] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1360] <= 1'b0;
    end else if(N1257) begin
      btb_q[1360] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1359] <= 1'b0;
    end else if(N1257) begin
      btb_q[1359] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1358] <= 1'b0;
    end else if(N1257) begin
      btb_q[1358] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1357] <= 1'b0;
    end else if(N1257) begin
      btb_q[1357] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1356] <= 1'b0;
    end else if(N1257) begin
      btb_q[1356] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1355] <= 1'b0;
    end else if(N1257) begin
      btb_q[1355] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1354] <= 1'b0;
    end else if(N1257) begin
      btb_q[1354] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1353] <= 1'b0;
    end else if(N1257) begin
      btb_q[1353] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1352] <= 1'b0;
    end else if(N1257) begin
      btb_q[1352] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1351] <= 1'b0;
    end else if(N1257) begin
      btb_q[1351] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1350] <= 1'b0;
    end else if(N1257) begin
      btb_q[1350] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1349] <= 1'b0;
    end else if(N1257) begin
      btb_q[1349] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1348] <= 1'b0;
    end else if(N1257) begin
      btb_q[1348] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1347] <= 1'b0;
    end else if(N1257) begin
      btb_q[1347] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1346] <= 1'b0;
    end else if(N1257) begin
      btb_q[1346] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1345] <= 1'b0;
    end else if(N1257) begin
      btb_q[1345] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1344] <= 1'b0;
    end else if(N1257) begin
      btb_q[1344] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1343] <= 1'b0;
    end else if(N1258) begin
      btb_q[1343] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1342] <= 1'b0;
    end else if(N1258) begin
      btb_q[1342] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1341] <= 1'b0;
    end else if(N1258) begin
      btb_q[1341] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1340] <= 1'b0;
    end else if(N1258) begin
      btb_q[1340] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1339] <= 1'b0;
    end else if(N1258) begin
      btb_q[1339] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1338] <= 1'b0;
    end else if(N1258) begin
      btb_q[1338] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1337] <= 1'b0;
    end else if(N1258) begin
      btb_q[1337] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1336] <= 1'b0;
    end else if(N1258) begin
      btb_q[1336] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1335] <= 1'b0;
    end else if(N1258) begin
      btb_q[1335] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1334] <= 1'b0;
    end else if(N1258) begin
      btb_q[1334] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1333] <= 1'b0;
    end else if(N1258) begin
      btb_q[1333] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1332] <= 1'b0;
    end else if(N1258) begin
      btb_q[1332] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1331] <= 1'b0;
    end else if(N1258) begin
      btb_q[1331] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1330] <= 1'b0;
    end else if(N1258) begin
      btb_q[1330] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1329] <= 1'b0;
    end else if(N1258) begin
      btb_q[1329] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1328] <= 1'b0;
    end else if(N1258) begin
      btb_q[1328] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1327] <= 1'b0;
    end else if(N1258) begin
      btb_q[1327] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1326] <= 1'b0;
    end else if(N1258) begin
      btb_q[1326] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1325] <= 1'b0;
    end else if(N1258) begin
      btb_q[1325] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1324] <= 1'b0;
    end else if(N1258) begin
      btb_q[1324] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1323] <= 1'b0;
    end else if(N1258) begin
      btb_q[1323] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1322] <= 1'b0;
    end else if(N1258) begin
      btb_q[1322] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1321] <= 1'b0;
    end else if(N1258) begin
      btb_q[1321] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1320] <= 1'b0;
    end else if(N1258) begin
      btb_q[1320] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1319] <= 1'b0;
    end else if(N1258) begin
      btb_q[1319] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1318] <= 1'b0;
    end else if(N1258) begin
      btb_q[1318] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1317] <= 1'b0;
    end else if(N1258) begin
      btb_q[1317] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1316] <= 1'b0;
    end else if(N1258) begin
      btb_q[1316] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1315] <= 1'b0;
    end else if(N1258) begin
      btb_q[1315] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1314] <= 1'b0;
    end else if(N1258) begin
      btb_q[1314] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1313] <= 1'b0;
    end else if(N1258) begin
      btb_q[1313] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1312] <= 1'b0;
    end else if(N1258) begin
      btb_q[1312] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1311] <= 1'b0;
    end else if(N1258) begin
      btb_q[1311] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1310] <= 1'b0;
    end else if(N1258) begin
      btb_q[1310] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1309] <= 1'b0;
    end else if(N1258) begin
      btb_q[1309] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1308] <= 1'b0;
    end else if(N1258) begin
      btb_q[1308] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1307] <= 1'b0;
    end else if(N1258) begin
      btb_q[1307] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1306] <= 1'b0;
    end else if(N1262) begin
      btb_q[1306] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1305] <= 1'b0;
    end else if(N1262) begin
      btb_q[1305] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1304] <= 1'b0;
    end else if(N1262) begin
      btb_q[1304] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1303] <= 1'b0;
    end else if(N1262) begin
      btb_q[1303] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1302] <= 1'b0;
    end else if(N1262) begin
      btb_q[1302] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1301] <= 1'b0;
    end else if(N1262) begin
      btb_q[1301] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1300] <= 1'b0;
    end else if(N1262) begin
      btb_q[1300] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1299] <= 1'b0;
    end else if(N1253) begin
      btb_q[1299] <= N549;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1298] <= 1'b0;
    end else if(N1266) begin
      btb_q[1298] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1297] <= 1'b0;
    end else if(N1266) begin
      btb_q[1297] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1296] <= 1'b0;
    end else if(N1266) begin
      btb_q[1296] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1295] <= 1'b0;
    end else if(N1266) begin
      btb_q[1295] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1294] <= 1'b0;
    end else if(N1266) begin
      btb_q[1294] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1293] <= 1'b0;
    end else if(N1266) begin
      btb_q[1293] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1292] <= 1'b0;
    end else if(N1266) begin
      btb_q[1292] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1291] <= 1'b0;
    end else if(N1266) begin
      btb_q[1291] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1290] <= 1'b0;
    end else if(N1266) begin
      btb_q[1290] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1289] <= 1'b0;
    end else if(N1266) begin
      btb_q[1289] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1288] <= 1'b0;
    end else if(N1266) begin
      btb_q[1288] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1287] <= 1'b0;
    end else if(N1266) begin
      btb_q[1287] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1286] <= 1'b0;
    end else if(N1269) begin
      btb_q[1286] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1285] <= 1'b0;
    end else if(N1269) begin
      btb_q[1285] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1284] <= 1'b0;
    end else if(N1269) begin
      btb_q[1284] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1283] <= 1'b0;
    end else if(N1269) begin
      btb_q[1283] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1282] <= 1'b0;
    end else if(N1269) begin
      btb_q[1282] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1281] <= 1'b0;
    end else if(N1269) begin
      btb_q[1281] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1280] <= 1'b0;
    end else if(N1269) begin
      btb_q[1280] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1279] <= 1'b0;
    end else if(N1269) begin
      btb_q[1279] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1278] <= 1'b0;
    end else if(N1269) begin
      btb_q[1278] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1277] <= 1'b0;
    end else if(N1269) begin
      btb_q[1277] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1276] <= 1'b0;
    end else if(N1269) begin
      btb_q[1276] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1275] <= 1'b0;
    end else if(N1269) begin
      btb_q[1275] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1274] <= 1'b0;
    end else if(N1269) begin
      btb_q[1274] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1273] <= 1'b0;
    end else if(N1269) begin
      btb_q[1273] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1272] <= 1'b0;
    end else if(N1269) begin
      btb_q[1272] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1271] <= 1'b0;
    end else if(N1269) begin
      btb_q[1271] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1270] <= 1'b0;
    end else if(N1269) begin
      btb_q[1270] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1269] <= 1'b0;
    end else if(N1269) begin
      btb_q[1269] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1268] <= 1'b0;
    end else if(N1269) begin
      btb_q[1268] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1267] <= 1'b0;
    end else if(N1269) begin
      btb_q[1267] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1266] <= 1'b0;
    end else if(N1269) begin
      btb_q[1266] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1265] <= 1'b0;
    end else if(N1269) begin
      btb_q[1265] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1264] <= 1'b0;
    end else if(N1269) begin
      btb_q[1264] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1263] <= 1'b0;
    end else if(N1269) begin
      btb_q[1263] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1262] <= 1'b0;
    end else if(N1269) begin
      btb_q[1262] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1261] <= 1'b0;
    end else if(N1269) begin
      btb_q[1261] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1260] <= 1'b0;
    end else if(N1269) begin
      btb_q[1260] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1259] <= 1'b0;
    end else if(N1269) begin
      btb_q[1259] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1258] <= 1'b0;
    end else if(N1269) begin
      btb_q[1258] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1257] <= 1'b0;
    end else if(N1269) begin
      btb_q[1257] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1256] <= 1'b0;
    end else if(N1269) begin
      btb_q[1256] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1255] <= 1'b0;
    end else if(N1269) begin
      btb_q[1255] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1254] <= 1'b0;
    end else if(N1269) begin
      btb_q[1254] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1253] <= 1'b0;
    end else if(N1269) begin
      btb_q[1253] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1252] <= 1'b0;
    end else if(N1269) begin
      btb_q[1252] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1251] <= 1'b0;
    end else if(N1269) begin
      btb_q[1251] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1250] <= 1'b0;
    end else if(N1269) begin
      btb_q[1250] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1249] <= 1'b0;
    end else if(N1269) begin
      btb_q[1249] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1248] <= 1'b0;
    end else if(N1269) begin
      btb_q[1248] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1247] <= 1'b0;
    end else if(N1269) begin
      btb_q[1247] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1246] <= 1'b0;
    end else if(N1269) begin
      btb_q[1246] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1245] <= 1'b0;
    end else if(N1269) begin
      btb_q[1245] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1244] <= 1'b0;
    end else if(N1269) begin
      btb_q[1244] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1243] <= 1'b0;
    end else if(N1270) begin
      btb_q[1243] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1242] <= 1'b0;
    end else if(N1270) begin
      btb_q[1242] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1241] <= 1'b0;
    end else if(N1270) begin
      btb_q[1241] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1240] <= 1'b0;
    end else if(N1270) begin
      btb_q[1240] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1239] <= 1'b0;
    end else if(N1270) begin
      btb_q[1239] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1238] <= 1'b0;
    end else if(N1270) begin
      btb_q[1238] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1237] <= 1'b0;
    end else if(N1270) begin
      btb_q[1237] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1236] <= 1'b0;
    end else if(N1270) begin
      btb_q[1236] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1235] <= 1'b0;
    end else if(N1270) begin
      btb_q[1235] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1234] <= 1'b0;
    end else if(N1271) begin
      btb_q[1234] <= N548;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1233] <= 1'b0;
    end else if(N1275) begin
      btb_q[1233] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1232] <= 1'b0;
    end else if(N1275) begin
      btb_q[1232] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1231] <= 1'b0;
    end else if(N1275) begin
      btb_q[1231] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1230] <= 1'b0;
    end else if(N1275) begin
      btb_q[1230] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1229] <= 1'b0;
    end else if(N1275) begin
      btb_q[1229] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1228] <= 1'b0;
    end else if(N1275) begin
      btb_q[1228] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1227] <= 1'b0;
    end else if(N1275) begin
      btb_q[1227] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1226] <= 1'b0;
    end else if(N1275) begin
      btb_q[1226] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1225] <= 1'b0;
    end else if(N1275) begin
      btb_q[1225] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1224] <= 1'b0;
    end else if(N1275) begin
      btb_q[1224] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1223] <= 1'b0;
    end else if(N1275) begin
      btb_q[1223] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1222] <= 1'b0;
    end else if(N1275) begin
      btb_q[1222] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1221] <= 1'b0;
    end else if(N1275) begin
      btb_q[1221] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1220] <= 1'b0;
    end else if(N1275) begin
      btb_q[1220] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1219] <= 1'b0;
    end else if(N1275) begin
      btb_q[1219] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1218] <= 1'b0;
    end else if(N1275) begin
      btb_q[1218] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1217] <= 1'b0;
    end else if(N1275) begin
      btb_q[1217] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1216] <= 1'b0;
    end else if(N1275) begin
      btb_q[1216] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1215] <= 1'b0;
    end else if(N1275) begin
      btb_q[1215] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1214] <= 1'b0;
    end else if(N1275) begin
      btb_q[1214] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1213] <= 1'b0;
    end else if(N1275) begin
      btb_q[1213] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1212] <= 1'b0;
    end else if(N1275) begin
      btb_q[1212] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1211] <= 1'b0;
    end else if(N1275) begin
      btb_q[1211] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1210] <= 1'b0;
    end else if(N1275) begin
      btb_q[1210] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1209] <= 1'b0;
    end else if(N1275) begin
      btb_q[1209] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1208] <= 1'b0;
    end else if(N1275) begin
      btb_q[1208] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1207] <= 1'b0;
    end else if(N1275) begin
      btb_q[1207] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1206] <= 1'b0;
    end else if(N1275) begin
      btb_q[1206] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1205] <= 1'b0;
    end else if(N1279) begin
      btb_q[1205] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1204] <= 1'b0;
    end else if(N1279) begin
      btb_q[1204] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1203] <= 1'b0;
    end else if(N1279) begin
      btb_q[1203] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1202] <= 1'b0;
    end else if(N1279) begin
      btb_q[1202] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1201] <= 1'b0;
    end else if(N1279) begin
      btb_q[1201] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1200] <= 1'b0;
    end else if(N1279) begin
      btb_q[1200] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1199] <= 1'b0;
    end else if(N1279) begin
      btb_q[1199] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1198] <= 1'b0;
    end else if(N1279) begin
      btb_q[1198] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1197] <= 1'b0;
    end else if(N1279) begin
      btb_q[1197] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1196] <= 1'b0;
    end else if(N1279) begin
      btb_q[1196] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1195] <= 1'b0;
    end else if(N1279) begin
      btb_q[1195] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1194] <= 1'b0;
    end else if(N1279) begin
      btb_q[1194] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1193] <= 1'b0;
    end else if(N1279) begin
      btb_q[1193] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1192] <= 1'b0;
    end else if(N1279) begin
      btb_q[1192] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1191] <= 1'b0;
    end else if(N1279) begin
      btb_q[1191] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1190] <= 1'b0;
    end else if(N1279) begin
      btb_q[1190] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1189] <= 1'b0;
    end else if(N1279) begin
      btb_q[1189] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1188] <= 1'b0;
    end else if(N1279) begin
      btb_q[1188] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1187] <= 1'b0;
    end else if(N1282) begin
      btb_q[1187] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1186] <= 1'b0;
    end else if(N1282) begin
      btb_q[1186] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1185] <= 1'b0;
    end else if(N1282) begin
      btb_q[1185] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1184] <= 1'b0;
    end else if(N1282) begin
      btb_q[1184] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1183] <= 1'b0;
    end else if(N1282) begin
      btb_q[1183] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1182] <= 1'b0;
    end else if(N1282) begin
      btb_q[1182] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1181] <= 1'b0;
    end else if(N1282) begin
      btb_q[1181] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1180] <= 1'b0;
    end else if(N1282) begin
      btb_q[1180] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1179] <= 1'b0;
    end else if(N1282) begin
      btb_q[1179] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1178] <= 1'b0;
    end else if(N1282) begin
      btb_q[1178] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1177] <= 1'b0;
    end else if(N1282) begin
      btb_q[1177] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1176] <= 1'b0;
    end else if(N1282) begin
      btb_q[1176] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1175] <= 1'b0;
    end else if(N1282) begin
      btb_q[1175] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1174] <= 1'b0;
    end else if(N1282) begin
      btb_q[1174] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1173] <= 1'b0;
    end else if(N1282) begin
      btb_q[1173] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1172] <= 1'b0;
    end else if(N1282) begin
      btb_q[1172] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1171] <= 1'b0;
    end else if(N1282) begin
      btb_q[1171] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1170] <= 1'b0;
    end else if(N1282) begin
      btb_q[1170] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1169] <= 1'b0;
    end else if(N1283) begin
      btb_q[1169] <= N547;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1168] <= 1'b0;
    end else if(N1287) begin
      btb_q[1168] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1167] <= 1'b0;
    end else if(N1287) begin
      btb_q[1167] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1166] <= 1'b0;
    end else if(N1287) begin
      btb_q[1166] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1165] <= 1'b0;
    end else if(N1287) begin
      btb_q[1165] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1164] <= 1'b0;
    end else if(N1287) begin
      btb_q[1164] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1163] <= 1'b0;
    end else if(N1287) begin
      btb_q[1163] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1162] <= 1'b0;
    end else if(N1287) begin
      btb_q[1162] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1161] <= 1'b0;
    end else if(N1287) begin
      btb_q[1161] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1160] <= 1'b0;
    end else if(N1287) begin
      btb_q[1160] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1159] <= 1'b0;
    end else if(N1287) begin
      btb_q[1159] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1158] <= 1'b0;
    end else if(N1287) begin
      btb_q[1158] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1157] <= 1'b0;
    end else if(N1287) begin
      btb_q[1157] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1156] <= 1'b0;
    end else if(N1287) begin
      btb_q[1156] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1155] <= 1'b0;
    end else if(N1287) begin
      btb_q[1155] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1154] <= 1'b0;
    end else if(N1287) begin
      btb_q[1154] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1153] <= 1'b0;
    end else if(N1287) begin
      btb_q[1153] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1152] <= 1'b0;
    end else if(N1287) begin
      btb_q[1152] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1151] <= 1'b0;
    end else if(N1287) begin
      btb_q[1151] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1150] <= 1'b0;
    end else if(N1287) begin
      btb_q[1150] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1149] <= 1'b0;
    end else if(N1287) begin
      btb_q[1149] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1148] <= 1'b0;
    end else if(N1287) begin
      btb_q[1148] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1147] <= 1'b0;
    end else if(N1287) begin
      btb_q[1147] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1146] <= 1'b0;
    end else if(N1287) begin
      btb_q[1146] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1145] <= 1'b0;
    end else if(N1287) begin
      btb_q[1145] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1144] <= 1'b0;
    end else if(N1287) begin
      btb_q[1144] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1143] <= 1'b0;
    end else if(N1287) begin
      btb_q[1143] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1142] <= 1'b0;
    end else if(N1288) begin
      btb_q[1142] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1141] <= 1'b0;
    end else if(N1288) begin
      btb_q[1141] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1140] <= 1'b0;
    end else if(N1288) begin
      btb_q[1140] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1139] <= 1'b0;
    end else if(N1288) begin
      btb_q[1139] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1138] <= 1'b0;
    end else if(N1288) begin
      btb_q[1138] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1137] <= 1'b0;
    end else if(N1288) begin
      btb_q[1137] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1136] <= 1'b0;
    end else if(N1288) begin
      btb_q[1136] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1135] <= 1'b0;
    end else if(N1288) begin
      btb_q[1135] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1134] <= 1'b0;
    end else if(N1288) begin
      btb_q[1134] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1133] <= 1'b0;
    end else if(N1288) begin
      btb_q[1133] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1132] <= 1'b0;
    end else if(N1288) begin
      btb_q[1132] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1131] <= 1'b0;
    end else if(N1288) begin
      btb_q[1131] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1130] <= 1'b0;
    end else if(N1288) begin
      btb_q[1130] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1129] <= 1'b0;
    end else if(N1288) begin
      btb_q[1129] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1128] <= 1'b0;
    end else if(N1288) begin
      btb_q[1128] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1127] <= 1'b0;
    end else if(N1288) begin
      btb_q[1127] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1126] <= 1'b0;
    end else if(N1288) begin
      btb_q[1126] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1125] <= 1'b0;
    end else if(N1288) begin
      btb_q[1125] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1124] <= 1'b0;
    end else if(N1288) begin
      btb_q[1124] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1123] <= 1'b0;
    end else if(N1288) begin
      btb_q[1123] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1122] <= 1'b0;
    end else if(N1288) begin
      btb_q[1122] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1121] <= 1'b0;
    end else if(N1288) begin
      btb_q[1121] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1120] <= 1'b0;
    end else if(N1288) begin
      btb_q[1120] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1119] <= 1'b0;
    end else if(N1288) begin
      btb_q[1119] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1118] <= 1'b0;
    end else if(N1288) begin
      btb_q[1118] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1117] <= 1'b0;
    end else if(N1288) begin
      btb_q[1117] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1116] <= 1'b0;
    end else if(N1288) begin
      btb_q[1116] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1115] <= 1'b0;
    end else if(N1288) begin
      btb_q[1115] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1114] <= 1'b0;
    end else if(N1288) begin
      btb_q[1114] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1113] <= 1'b0;
    end else if(N1288) begin
      btb_q[1113] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1112] <= 1'b0;
    end else if(N1288) begin
      btb_q[1112] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1111] <= 1'b0;
    end else if(N1288) begin
      btb_q[1111] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1110] <= 1'b0;
    end else if(N1288) begin
      btb_q[1110] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1109] <= 1'b0;
    end else if(N1288) begin
      btb_q[1109] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1108] <= 1'b0;
    end else if(N1288) begin
      btb_q[1108] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1107] <= 1'b0;
    end else if(N1288) begin
      btb_q[1107] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1106] <= 1'b0;
    end else if(N1288) begin
      btb_q[1106] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1105] <= 1'b0;
    end else if(N1292) begin
      btb_q[1105] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1104] <= 1'b0;
    end else if(N1283) begin
      btb_q[1104] <= N546;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1103] <= 1'b0;
    end else if(N1296) begin
      btb_q[1103] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1102] <= 1'b0;
    end else if(N1296) begin
      btb_q[1102] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1101] <= 1'b0;
    end else if(N1296) begin
      btb_q[1101] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1100] <= 1'b0;
    end else if(N1296) begin
      btb_q[1100] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1099] <= 1'b0;
    end else if(N1296) begin
      btb_q[1099] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1098] <= 1'b0;
    end else if(N1296) begin
      btb_q[1098] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1097] <= 1'b0;
    end else if(N1296) begin
      btb_q[1097] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1096] <= 1'b0;
    end else if(N1296) begin
      btb_q[1096] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1095] <= 1'b0;
    end else if(N1296) begin
      btb_q[1095] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1094] <= 1'b0;
    end else if(N1296) begin
      btb_q[1094] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1093] <= 1'b0;
    end else if(N1296) begin
      btb_q[1093] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1092] <= 1'b0;
    end else if(N1296) begin
      btb_q[1092] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1091] <= 1'b0;
    end else if(N1296) begin
      btb_q[1091] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1090] <= 1'b0;
    end else if(N1296) begin
      btb_q[1090] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1089] <= 1'b0;
    end else if(N1296) begin
      btb_q[1089] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1088] <= 1'b0;
    end else if(N1299) begin
      btb_q[1088] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1087] <= 1'b0;
    end else if(N1299) begin
      btb_q[1087] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1086] <= 1'b0;
    end else if(N1299) begin
      btb_q[1086] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1085] <= 1'b0;
    end else if(N1299) begin
      btb_q[1085] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1084] <= 1'b0;
    end else if(N1299) begin
      btb_q[1084] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1083] <= 1'b0;
    end else if(N1299) begin
      btb_q[1083] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1082] <= 1'b0;
    end else if(N1299) begin
      btb_q[1082] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1081] <= 1'b0;
    end else if(N1299) begin
      btb_q[1081] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1080] <= 1'b0;
    end else if(N1299) begin
      btb_q[1080] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1079] <= 1'b0;
    end else if(N1299) begin
      btb_q[1079] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1078] <= 1'b0;
    end else if(N1299) begin
      btb_q[1078] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1077] <= 1'b0;
    end else if(N1299) begin
      btb_q[1077] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1076] <= 1'b0;
    end else if(N1299) begin
      btb_q[1076] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1075] <= 1'b0;
    end else if(N1299) begin
      btb_q[1075] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1074] <= 1'b0;
    end else if(N1299) begin
      btb_q[1074] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1073] <= 1'b0;
    end else if(N1299) begin
      btb_q[1073] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1072] <= 1'b0;
    end else if(N1299) begin
      btb_q[1072] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1071] <= 1'b0;
    end else if(N1299) begin
      btb_q[1071] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1070] <= 1'b0;
    end else if(N1299) begin
      btb_q[1070] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1069] <= 1'b0;
    end else if(N1299) begin
      btb_q[1069] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1068] <= 1'b0;
    end else if(N1299) begin
      btb_q[1068] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1067] <= 1'b0;
    end else if(N1299) begin
      btb_q[1067] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1066] <= 1'b0;
    end else if(N1299) begin
      btb_q[1066] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1065] <= 1'b0;
    end else if(N1299) begin
      btb_q[1065] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1064] <= 1'b0;
    end else if(N1299) begin
      btb_q[1064] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1063] <= 1'b0;
    end else if(N1299) begin
      btb_q[1063] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1062] <= 1'b0;
    end else if(N1299) begin
      btb_q[1062] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1061] <= 1'b0;
    end else if(N1299) begin
      btb_q[1061] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1060] <= 1'b0;
    end else if(N1299) begin
      btb_q[1060] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1059] <= 1'b0;
    end else if(N1299) begin
      btb_q[1059] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1058] <= 1'b0;
    end else if(N1299) begin
      btb_q[1058] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1057] <= 1'b0;
    end else if(N1299) begin
      btb_q[1057] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1056] <= 1'b0;
    end else if(N1299) begin
      btb_q[1056] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1055] <= 1'b0;
    end else if(N1299) begin
      btb_q[1055] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1054] <= 1'b0;
    end else if(N1299) begin
      btb_q[1054] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1053] <= 1'b0;
    end else if(N1299) begin
      btb_q[1053] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1052] <= 1'b0;
    end else if(N1299) begin
      btb_q[1052] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1051] <= 1'b0;
    end else if(N1299) begin
      btb_q[1051] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1050] <= 1'b0;
    end else if(N1299) begin
      btb_q[1050] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1049] <= 1'b0;
    end else if(N1299) begin
      btb_q[1049] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1048] <= 1'b0;
    end else if(N1299) begin
      btb_q[1048] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1047] <= 1'b0;
    end else if(N1299) begin
      btb_q[1047] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1046] <= 1'b0;
    end else if(N1299) begin
      btb_q[1046] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1045] <= 1'b0;
    end else if(N1299) begin
      btb_q[1045] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1044] <= 1'b0;
    end else if(N1299) begin
      btb_q[1044] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1043] <= 1'b0;
    end else if(N1299) begin
      btb_q[1043] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1042] <= 1'b0;
    end else if(N1300) begin
      btb_q[1042] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1041] <= 1'b0;
    end else if(N1300) begin
      btb_q[1041] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1040] <= 1'b0;
    end else if(N1300) begin
      btb_q[1040] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1039] <= 1'b0;
    end else if(N1301) begin
      btb_q[1039] <= N545;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1038] <= 1'b0;
    end else if(N1305) begin
      btb_q[1038] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1037] <= 1'b0;
    end else if(N1305) begin
      btb_q[1037] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1036] <= 1'b0;
    end else if(N1305) begin
      btb_q[1036] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1035] <= 1'b0;
    end else if(N1305) begin
      btb_q[1035] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1034] <= 1'b0;
    end else if(N1305) begin
      btb_q[1034] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1033] <= 1'b0;
    end else if(N1305) begin
      btb_q[1033] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1032] <= 1'b0;
    end else if(N1305) begin
      btb_q[1032] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1031] <= 1'b0;
    end else if(N1305) begin
      btb_q[1031] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1030] <= 1'b0;
    end else if(N1305) begin
      btb_q[1030] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1029] <= 1'b0;
    end else if(N1305) begin
      btb_q[1029] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1028] <= 1'b0;
    end else if(N1305) begin
      btb_q[1028] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1027] <= 1'b0;
    end else if(N1305) begin
      btb_q[1027] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1026] <= 1'b0;
    end else if(N1305) begin
      btb_q[1026] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1025] <= 1'b0;
    end else if(N1305) begin
      btb_q[1025] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1024] <= 1'b0;
    end else if(N1305) begin
      btb_q[1024] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1023] <= 1'b0;
    end else if(N1305) begin
      btb_q[1023] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1022] <= 1'b0;
    end else if(N1305) begin
      btb_q[1022] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1021] <= 1'b0;
    end else if(N1305) begin
      btb_q[1021] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1020] <= 1'b0;
    end else if(N1305) begin
      btb_q[1020] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1019] <= 1'b0;
    end else if(N1305) begin
      btb_q[1019] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1018] <= 1'b0;
    end else if(N1305) begin
      btb_q[1018] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1017] <= 1'b0;
    end else if(N1305) begin
      btb_q[1017] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1016] <= 1'b0;
    end else if(N1305) begin
      btb_q[1016] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1015] <= 1'b0;
    end else if(N1305) begin
      btb_q[1015] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1014] <= 1'b0;
    end else if(N1305) begin
      btb_q[1014] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1013] <= 1'b0;
    end else if(N1305) begin
      btb_q[1013] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1012] <= 1'b0;
    end else if(N1305) begin
      btb_q[1012] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1011] <= 1'b0;
    end else if(N1305) begin
      btb_q[1011] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1010] <= 1'b0;
    end else if(N1305) begin
      btb_q[1010] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1009] <= 1'b0;
    end else if(N1305) begin
      btb_q[1009] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1008] <= 1'b0;
    end else if(N1305) begin
      btb_q[1008] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1007] <= 1'b0;
    end else if(N1305) begin
      btb_q[1007] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1006] <= 1'b0;
    end else if(N1305) begin
      btb_q[1006] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1005] <= 1'b0;
    end else if(N1305) begin
      btb_q[1005] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1004] <= 1'b0;
    end else if(N1309) begin
      btb_q[1004] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1003] <= 1'b0;
    end else if(N1309) begin
      btb_q[1003] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1002] <= 1'b0;
    end else if(N1309) begin
      btb_q[1002] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1001] <= 1'b0;
    end else if(N1309) begin
      btb_q[1001] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1000] <= 1'b0;
    end else if(N1309) begin
      btb_q[1000] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[999] <= 1'b0;
    end else if(N1309) begin
      btb_q[999] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[998] <= 1'b0;
    end else if(N1309) begin
      btb_q[998] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[997] <= 1'b0;
    end else if(N1309) begin
      btb_q[997] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[996] <= 1'b0;
    end else if(N1309) begin
      btb_q[996] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[995] <= 1'b0;
    end else if(N1309) begin
      btb_q[995] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[994] <= 1'b0;
    end else if(N1309) begin
      btb_q[994] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[993] <= 1'b0;
    end else if(N1309) begin
      btb_q[993] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[992] <= 1'b0;
    end else if(N1309) begin
      btb_q[992] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[991] <= 1'b0;
    end else if(N1309) begin
      btb_q[991] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[990] <= 1'b0;
    end else if(N1309) begin
      btb_q[990] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[989] <= 1'b0;
    end else if(N1312) begin
      btb_q[989] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[988] <= 1'b0;
    end else if(N1312) begin
      btb_q[988] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[987] <= 1'b0;
    end else if(N1312) begin
      btb_q[987] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[986] <= 1'b0;
    end else if(N1312) begin
      btb_q[986] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[985] <= 1'b0;
    end else if(N1312) begin
      btb_q[985] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[984] <= 1'b0;
    end else if(N1312) begin
      btb_q[984] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[983] <= 1'b0;
    end else if(N1312) begin
      btb_q[983] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[982] <= 1'b0;
    end else if(N1312) begin
      btb_q[982] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[981] <= 1'b0;
    end else if(N1312) begin
      btb_q[981] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[980] <= 1'b0;
    end else if(N1312) begin
      btb_q[980] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[979] <= 1'b0;
    end else if(N1312) begin
      btb_q[979] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[978] <= 1'b0;
    end else if(N1312) begin
      btb_q[978] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[977] <= 1'b0;
    end else if(N1312) begin
      btb_q[977] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[976] <= 1'b0;
    end else if(N1312) begin
      btb_q[976] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[975] <= 1'b0;
    end else if(N1312) begin
      btb_q[975] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[974] <= 1'b0;
    end else if(N1313) begin
      btb_q[974] <= N544;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[973] <= 1'b0;
    end else if(N1317) begin
      btb_q[973] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[972] <= 1'b0;
    end else if(N1317) begin
      btb_q[972] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[971] <= 1'b0;
    end else if(N1317) begin
      btb_q[971] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[970] <= 1'b0;
    end else if(N1317) begin
      btb_q[970] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[969] <= 1'b0;
    end else if(N1317) begin
      btb_q[969] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[968] <= 1'b0;
    end else if(N1317) begin
      btb_q[968] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[967] <= 1'b0;
    end else if(N1317) begin
      btb_q[967] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[966] <= 1'b0;
    end else if(N1317) begin
      btb_q[966] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[965] <= 1'b0;
    end else if(N1317) begin
      btb_q[965] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[964] <= 1'b0;
    end else if(N1317) begin
      btb_q[964] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[963] <= 1'b0;
    end else if(N1317) begin
      btb_q[963] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[962] <= 1'b0;
    end else if(N1317) begin
      btb_q[962] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[961] <= 1'b0;
    end else if(N1317) begin
      btb_q[961] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[960] <= 1'b0;
    end else if(N1317) begin
      btb_q[960] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[959] <= 1'b0;
    end else if(N1317) begin
      btb_q[959] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[958] <= 1'b0;
    end else if(N1317) begin
      btb_q[958] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[957] <= 1'b0;
    end else if(N1317) begin
      btb_q[957] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[956] <= 1'b0;
    end else if(N1317) begin
      btb_q[956] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[955] <= 1'b0;
    end else if(N1317) begin
      btb_q[955] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[954] <= 1'b0;
    end else if(N1317) begin
      btb_q[954] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[953] <= 1'b0;
    end else if(N1317) begin
      btb_q[953] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[952] <= 1'b0;
    end else if(N1317) begin
      btb_q[952] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[951] <= 1'b0;
    end else if(N1317) begin
      btb_q[951] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[950] <= 1'b0;
    end else if(N1317) begin
      btb_q[950] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[949] <= 1'b0;
    end else if(N1317) begin
      btb_q[949] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[948] <= 1'b0;
    end else if(N1317) begin
      btb_q[948] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[947] <= 1'b0;
    end else if(N1317) begin
      btb_q[947] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[946] <= 1'b0;
    end else if(N1317) begin
      btb_q[946] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[945] <= 1'b0;
    end else if(N1317) begin
      btb_q[945] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[944] <= 1'b0;
    end else if(N1317) begin
      btb_q[944] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[943] <= 1'b0;
    end else if(N1317) begin
      btb_q[943] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[942] <= 1'b0;
    end else if(N1317) begin
      btb_q[942] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[941] <= 1'b0;
    end else if(N1318) begin
      btb_q[941] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[940] <= 1'b0;
    end else if(N1318) begin
      btb_q[940] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[939] <= 1'b0;
    end else if(N1318) begin
      btb_q[939] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[938] <= 1'b0;
    end else if(N1318) begin
      btb_q[938] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[937] <= 1'b0;
    end else if(N1318) begin
      btb_q[937] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[936] <= 1'b0;
    end else if(N1318) begin
      btb_q[936] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[935] <= 1'b0;
    end else if(N1318) begin
      btb_q[935] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[934] <= 1'b0;
    end else if(N1318) begin
      btb_q[934] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[933] <= 1'b0;
    end else if(N1318) begin
      btb_q[933] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[932] <= 1'b0;
    end else if(N1318) begin
      btb_q[932] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[931] <= 1'b0;
    end else if(N1318) begin
      btb_q[931] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[930] <= 1'b0;
    end else if(N1318) begin
      btb_q[930] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[929] <= 1'b0;
    end else if(N1318) begin
      btb_q[929] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[928] <= 1'b0;
    end else if(N1318) begin
      btb_q[928] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[927] <= 1'b0;
    end else if(N1318) begin
      btb_q[927] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[926] <= 1'b0;
    end else if(N1318) begin
      btb_q[926] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[925] <= 1'b0;
    end else if(N1318) begin
      btb_q[925] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[924] <= 1'b0;
    end else if(N1318) begin
      btb_q[924] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[923] <= 1'b0;
    end else if(N1318) begin
      btb_q[923] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[922] <= 1'b0;
    end else if(N1318) begin
      btb_q[922] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[921] <= 1'b0;
    end else if(N1318) begin
      btb_q[921] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[920] <= 1'b0;
    end else if(N1318) begin
      btb_q[920] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[919] <= 1'b0;
    end else if(N1318) begin
      btb_q[919] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[918] <= 1'b0;
    end else if(N1318) begin
      btb_q[918] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[917] <= 1'b0;
    end else if(N1318) begin
      btb_q[917] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[916] <= 1'b0;
    end else if(N1318) begin
      btb_q[916] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[915] <= 1'b0;
    end else if(N1318) begin
      btb_q[915] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[914] <= 1'b0;
    end else if(N1318) begin
      btb_q[914] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[913] <= 1'b0;
    end else if(N1318) begin
      btb_q[913] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[912] <= 1'b0;
    end else if(N1318) begin
      btb_q[912] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[911] <= 1'b0;
    end else if(N1318) begin
      btb_q[911] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[910] <= 1'b0;
    end else if(N1318) begin
      btb_q[910] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[909] <= 1'b0;
    end else if(N1313) begin
      btb_q[909] <= N543;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[908] <= 1'b0;
    end else if(N1322) begin
      btb_q[908] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[907] <= 1'b0;
    end else if(N1322) begin
      btb_q[907] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[906] <= 1'b0;
    end else if(N1322) begin
      btb_q[906] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[905] <= 1'b0;
    end else if(N1322) begin
      btb_q[905] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[904] <= 1'b0;
    end else if(N1322) begin
      btb_q[904] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[903] <= 1'b0;
    end else if(N1326) begin
      btb_q[903] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[902] <= 1'b0;
    end else if(N1326) begin
      btb_q[902] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[901] <= 1'b0;
    end else if(N1326) begin
      btb_q[901] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[900] <= 1'b0;
    end else if(N1326) begin
      btb_q[900] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[899] <= 1'b0;
    end else if(N1326) begin
      btb_q[899] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[898] <= 1'b0;
    end else if(N1326) begin
      btb_q[898] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[897] <= 1'b0;
    end else if(N1326) begin
      btb_q[897] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[896] <= 1'b0;
    end else if(N1326) begin
      btb_q[896] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[895] <= 1'b0;
    end else if(N1326) begin
      btb_q[895] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[894] <= 1'b0;
    end else if(N1326) begin
      btb_q[894] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[893] <= 1'b0;
    end else if(N1326) begin
      btb_q[893] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[892] <= 1'b0;
    end else if(N1326) begin
      btb_q[892] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[891] <= 1'b0;
    end else if(N1326) begin
      btb_q[891] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[890] <= 1'b0;
    end else if(N1329) begin
      btb_q[890] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[889] <= 1'b0;
    end else if(N1329) begin
      btb_q[889] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[888] <= 1'b0;
    end else if(N1329) begin
      btb_q[888] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[887] <= 1'b0;
    end else if(N1329) begin
      btb_q[887] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[886] <= 1'b0;
    end else if(N1329) begin
      btb_q[886] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[885] <= 1'b0;
    end else if(N1329) begin
      btb_q[885] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[884] <= 1'b0;
    end else if(N1329) begin
      btb_q[884] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[883] <= 1'b0;
    end else if(N1329) begin
      btb_q[883] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[882] <= 1'b0;
    end else if(N1329) begin
      btb_q[882] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[881] <= 1'b0;
    end else if(N1329) begin
      btb_q[881] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[880] <= 1'b0;
    end else if(N1329) begin
      btb_q[880] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[879] <= 1'b0;
    end else if(N1329) begin
      btb_q[879] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[878] <= 1'b0;
    end else if(N1329) begin
      btb_q[878] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[877] <= 1'b0;
    end else if(N1329) begin
      btb_q[877] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[876] <= 1'b0;
    end else if(N1329) begin
      btb_q[876] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[875] <= 1'b0;
    end else if(N1329) begin
      btb_q[875] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[874] <= 1'b0;
    end else if(N1329) begin
      btb_q[874] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[873] <= 1'b0;
    end else if(N1329) begin
      btb_q[873] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[872] <= 1'b0;
    end else if(N1329) begin
      btb_q[872] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[871] <= 1'b0;
    end else if(N1329) begin
      btb_q[871] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[870] <= 1'b0;
    end else if(N1329) begin
      btb_q[870] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[869] <= 1'b0;
    end else if(N1329) begin
      btb_q[869] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[868] <= 1'b0;
    end else if(N1329) begin
      btb_q[868] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[867] <= 1'b0;
    end else if(N1329) begin
      btb_q[867] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[866] <= 1'b0;
    end else if(N1329) begin
      btb_q[866] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[865] <= 1'b0;
    end else if(N1329) begin
      btb_q[865] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[864] <= 1'b0;
    end else if(N1329) begin
      btb_q[864] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[863] <= 1'b0;
    end else if(N1329) begin
      btb_q[863] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[862] <= 1'b0;
    end else if(N1329) begin
      btb_q[862] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[861] <= 1'b0;
    end else if(N1329) begin
      btb_q[861] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[860] <= 1'b0;
    end else if(N1329) begin
      btb_q[860] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[859] <= 1'b0;
    end else if(N1329) begin
      btb_q[859] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[858] <= 1'b0;
    end else if(N1329) begin
      btb_q[858] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[857] <= 1'b0;
    end else if(N1329) begin
      btb_q[857] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[856] <= 1'b0;
    end else if(N1329) begin
      btb_q[856] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[855] <= 1'b0;
    end else if(N1329) begin
      btb_q[855] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[854] <= 1'b0;
    end else if(N1329) begin
      btb_q[854] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[853] <= 1'b0;
    end else if(N1329) begin
      btb_q[853] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[852] <= 1'b0;
    end else if(N1329) begin
      btb_q[852] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[851] <= 1'b0;
    end else if(N1329) begin
      btb_q[851] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[850] <= 1'b0;
    end else if(N1329) begin
      btb_q[850] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[849] <= 1'b0;
    end else if(N1329) begin
      btb_q[849] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[848] <= 1'b0;
    end else if(N1329) begin
      btb_q[848] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[847] <= 1'b0;
    end else if(N1329) begin
      btb_q[847] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[846] <= 1'b0;
    end else if(N1329) begin
      btb_q[846] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[845] <= 1'b0;
    end else if(N1329) begin
      btb_q[845] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[844] <= 1'b0;
    end else if(N1330) begin
      btb_q[844] <= N542;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[843] <= 1'b0;
    end else if(N1334) begin
      btb_q[843] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[842] <= 1'b0;
    end else if(N1334) begin
      btb_q[842] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[841] <= 1'b0;
    end else if(N1334) begin
      btb_q[841] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[840] <= 1'b0;
    end else if(N1335) begin
      btb_q[840] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[839] <= 1'b0;
    end else if(N1335) begin
      btb_q[839] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[838] <= 1'b0;
    end else if(N1335) begin
      btb_q[838] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[837] <= 1'b0;
    end else if(N1335) begin
      btb_q[837] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[836] <= 1'b0;
    end else if(N1335) begin
      btb_q[836] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[835] <= 1'b0;
    end else if(N1335) begin
      btb_q[835] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[834] <= 1'b0;
    end else if(N1335) begin
      btb_q[834] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[833] <= 1'b0;
    end else if(N1335) begin
      btb_q[833] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[832] <= 1'b0;
    end else if(N1335) begin
      btb_q[832] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[831] <= 1'b0;
    end else if(N1335) begin
      btb_q[831] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[830] <= 1'b0;
    end else if(N1335) begin
      btb_q[830] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[829] <= 1'b0;
    end else if(N1335) begin
      btb_q[829] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[828] <= 1'b0;
    end else if(N1335) begin
      btb_q[828] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[827] <= 1'b0;
    end else if(N1335) begin
      btb_q[827] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[826] <= 1'b0;
    end else if(N1335) begin
      btb_q[826] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[825] <= 1'b0;
    end else if(N1335) begin
      btb_q[825] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[824] <= 1'b0;
    end else if(N1335) begin
      btb_q[824] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[823] <= 1'b0;
    end else if(N1335) begin
      btb_q[823] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[822] <= 1'b0;
    end else if(N1335) begin
      btb_q[822] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[821] <= 1'b0;
    end else if(N1335) begin
      btb_q[821] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[820] <= 1'b0;
    end else if(N1335) begin
      btb_q[820] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[819] <= 1'b0;
    end else if(N1335) begin
      btb_q[819] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[818] <= 1'b0;
    end else if(N1335) begin
      btb_q[818] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[817] <= 1'b0;
    end else if(N1335) begin
      btb_q[817] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[816] <= 1'b0;
    end else if(N1335) begin
      btb_q[816] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[815] <= 1'b0;
    end else if(N1335) begin
      btb_q[815] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[814] <= 1'b0;
    end else if(N1335) begin
      btb_q[814] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[813] <= 1'b0;
    end else if(N1335) begin
      btb_q[813] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[812] <= 1'b0;
    end else if(N1335) begin
      btb_q[812] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[811] <= 1'b0;
    end else if(N1335) begin
      btb_q[811] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[810] <= 1'b0;
    end else if(N1335) begin
      btb_q[810] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[809] <= 1'b0;
    end else if(N1335) begin
      btb_q[809] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[808] <= 1'b0;
    end else if(N1335) begin
      btb_q[808] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[807] <= 1'b0;
    end else if(N1335) begin
      btb_q[807] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[806] <= 1'b0;
    end else if(N1335) begin
      btb_q[806] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[805] <= 1'b0;
    end else if(N1335) begin
      btb_q[805] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[804] <= 1'b0;
    end else if(N1335) begin
      btb_q[804] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[803] <= 1'b0;
    end else if(N1339) begin
      btb_q[803] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[802] <= 1'b0;
    end else if(N1339) begin
      btb_q[802] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[801] <= 1'b0;
    end else if(N1339) begin
      btb_q[801] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[800] <= 1'b0;
    end else if(N1339) begin
      btb_q[800] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[799] <= 1'b0;
    end else if(N1339) begin
      btb_q[799] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[798] <= 1'b0;
    end else if(N1339) begin
      btb_q[798] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[797] <= 1'b0;
    end else if(N1339) begin
      btb_q[797] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[796] <= 1'b0;
    end else if(N1339) begin
      btb_q[796] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[795] <= 1'b0;
    end else if(N1339) begin
      btb_q[795] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[794] <= 1'b0;
    end else if(N1339) begin
      btb_q[794] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[793] <= 1'b0;
    end else if(N1339) begin
      btb_q[793] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[792] <= 1'b0;
    end else if(N1339) begin
      btb_q[792] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[791] <= 1'b0;
    end else if(N1342) begin
      btb_q[791] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[790] <= 1'b0;
    end else if(N1342) begin
      btb_q[790] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[789] <= 1'b0;
    end else if(N1342) begin
      btb_q[789] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[788] <= 1'b0;
    end else if(N1342) begin
      btb_q[788] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[787] <= 1'b0;
    end else if(N1342) begin
      btb_q[787] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[786] <= 1'b0;
    end else if(N1342) begin
      btb_q[786] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[785] <= 1'b0;
    end else if(N1342) begin
      btb_q[785] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[784] <= 1'b0;
    end else if(N1342) begin
      btb_q[784] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[783] <= 1'b0;
    end else if(N1342) begin
      btb_q[783] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[782] <= 1'b0;
    end else if(N1342) begin
      btb_q[782] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[781] <= 1'b0;
    end else if(N1342) begin
      btb_q[781] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[780] <= 1'b0;
    end else if(N1342) begin
      btb_q[780] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[779] <= 1'b0;
    end else if(N1343) begin
      btb_q[779] <= N541;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[778] <= 1'b0;
    end else if(N1347) begin
      btb_q[778] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[777] <= 1'b0;
    end else if(N1347) begin
      btb_q[777] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[776] <= 1'b0;
    end else if(N1347) begin
      btb_q[776] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[775] <= 1'b0;
    end else if(N1347) begin
      btb_q[775] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[774] <= 1'b0;
    end else if(N1347) begin
      btb_q[774] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[773] <= 1'b0;
    end else if(N1347) begin
      btb_q[773] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[772] <= 1'b0;
    end else if(N1347) begin
      btb_q[772] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[771] <= 1'b0;
    end else if(N1347) begin
      btb_q[771] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[770] <= 1'b0;
    end else if(N1347) begin
      btb_q[770] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[769] <= 1'b0;
    end else if(N1347) begin
      btb_q[769] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[768] <= 1'b0;
    end else if(N1347) begin
      btb_q[768] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[767] <= 1'b0;
    end else if(N1347) begin
      btb_q[767] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[766] <= 1'b0;
    end else if(N1347) begin
      btb_q[766] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[765] <= 1'b0;
    end else if(N1347) begin
      btb_q[765] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[764] <= 1'b0;
    end else if(N1347) begin
      btb_q[764] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[763] <= 1'b0;
    end else if(N1347) begin
      btb_q[763] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[762] <= 1'b0;
    end else if(N1347) begin
      btb_q[762] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[761] <= 1'b0;
    end else if(N1347) begin
      btb_q[761] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[760] <= 1'b0;
    end else if(N1347) begin
      btb_q[760] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[759] <= 1'b0;
    end else if(N1347) begin
      btb_q[759] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[758] <= 1'b0;
    end else if(N1347) begin
      btb_q[758] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[757] <= 1'b0;
    end else if(N1347) begin
      btb_q[757] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[756] <= 1'b0;
    end else if(N1347) begin
      btb_q[756] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[755] <= 1'b0;
    end else if(N1347) begin
      btb_q[755] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[754] <= 1'b0;
    end else if(N1347) begin
      btb_q[754] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[753] <= 1'b0;
    end else if(N1347) begin
      btb_q[753] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[752] <= 1'b0;
    end else if(N1347) begin
      btb_q[752] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[751] <= 1'b0;
    end else if(N1347) begin
      btb_q[751] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[750] <= 1'b0;
    end else if(N1347) begin
      btb_q[750] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[749] <= 1'b0;
    end else if(N1347) begin
      btb_q[749] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[748] <= 1'b0;
    end else if(N1347) begin
      btb_q[748] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[747] <= 1'b0;
    end else if(N1347) begin
      btb_q[747] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[746] <= 1'b0;
    end else if(N1347) begin
      btb_q[746] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[745] <= 1'b0;
    end else if(N1347) begin
      btb_q[745] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[744] <= 1'b0;
    end else if(N1347) begin
      btb_q[744] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[743] <= 1'b0;
    end else if(N1347) begin
      btb_q[743] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[742] <= 1'b0;
    end else if(N1347) begin
      btb_q[742] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[741] <= 1'b0;
    end else if(N1347) begin
      btb_q[741] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[740] <= 1'b0;
    end else if(N1348) begin
      btb_q[740] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[739] <= 1'b0;
    end else if(N1348) begin
      btb_q[739] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[738] <= 1'b0;
    end else if(N1348) begin
      btb_q[738] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[737] <= 1'b0;
    end else if(N1348) begin
      btb_q[737] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[736] <= 1'b0;
    end else if(N1348) begin
      btb_q[736] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[735] <= 1'b0;
    end else if(N1348) begin
      btb_q[735] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[734] <= 1'b0;
    end else if(N1348) begin
      btb_q[734] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[733] <= 1'b0;
    end else if(N1348) begin
      btb_q[733] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[732] <= 1'b0;
    end else if(N1348) begin
      btb_q[732] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[731] <= 1'b0;
    end else if(N1348) begin
      btb_q[731] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[730] <= 1'b0;
    end else if(N1348) begin
      btb_q[730] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[729] <= 1'b0;
    end else if(N1348) begin
      btb_q[729] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[728] <= 1'b0;
    end else if(N1348) begin
      btb_q[728] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[727] <= 1'b0;
    end else if(N1348) begin
      btb_q[727] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[726] <= 1'b0;
    end else if(N1348) begin
      btb_q[726] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[725] <= 1'b0;
    end else if(N1348) begin
      btb_q[725] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[724] <= 1'b0;
    end else if(N1348) begin
      btb_q[724] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[723] <= 1'b0;
    end else if(N1348) begin
      btb_q[723] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[722] <= 1'b0;
    end else if(N1348) begin
      btb_q[722] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[721] <= 1'b0;
    end else if(N1348) begin
      btb_q[721] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[720] <= 1'b0;
    end else if(N1348) begin
      btb_q[720] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[719] <= 1'b0;
    end else if(N1348) begin
      btb_q[719] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[718] <= 1'b0;
    end else if(N1348) begin
      btb_q[718] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[717] <= 1'b0;
    end else if(N1348) begin
      btb_q[717] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[716] <= 1'b0;
    end else if(N1348) begin
      btb_q[716] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[715] <= 1'b0;
    end else if(N1348) begin
      btb_q[715] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[714] <= 1'b0;
    end else if(N1343) begin
      btb_q[714] <= N540;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[713] <= 1'b0;
    end else if(N1352) begin
      btb_q[713] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[712] <= 1'b0;
    end else if(N1352) begin
      btb_q[712] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[711] <= 1'b0;
    end else if(N1352) begin
      btb_q[711] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[710] <= 1'b0;
    end else if(N1352) begin
      btb_q[710] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[709] <= 1'b0;
    end else if(N1352) begin
      btb_q[709] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[708] <= 1'b0;
    end else if(N1352) begin
      btb_q[708] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[707] <= 1'b0;
    end else if(N1352) begin
      btb_q[707] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[706] <= 1'b0;
    end else if(N1352) begin
      btb_q[706] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[705] <= 1'b0;
    end else if(N1352) begin
      btb_q[705] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[704] <= 1'b0;
    end else if(N1352) begin
      btb_q[704] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[703] <= 1'b0;
    end else if(N1352) begin
      btb_q[703] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[702] <= 1'b0;
    end else if(N1356) begin
      btb_q[702] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[701] <= 1'b0;
    end else if(N1356) begin
      btb_q[701] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[700] <= 1'b0;
    end else if(N1356) begin
      btb_q[700] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[699] <= 1'b0;
    end else if(N1356) begin
      btb_q[699] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[698] <= 1'b0;
    end else if(N1356) begin
      btb_q[698] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[697] <= 1'b0;
    end else if(N1356) begin
      btb_q[697] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[696] <= 1'b0;
    end else if(N1356) begin
      btb_q[696] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[695] <= 1'b0;
    end else if(N1356) begin
      btb_q[695] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[694] <= 1'b0;
    end else if(N1356) begin
      btb_q[694] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[693] <= 1'b0;
    end else if(N1356) begin
      btb_q[693] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[692] <= 1'b0;
    end else if(N1359) begin
      btb_q[692] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[691] <= 1'b0;
    end else if(N1359) begin
      btb_q[691] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[690] <= 1'b0;
    end else if(N1359) begin
      btb_q[690] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[689] <= 1'b0;
    end else if(N1359) begin
      btb_q[689] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[688] <= 1'b0;
    end else if(N1359) begin
      btb_q[688] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[687] <= 1'b0;
    end else if(N1359) begin
      btb_q[687] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[686] <= 1'b0;
    end else if(N1359) begin
      btb_q[686] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[685] <= 1'b0;
    end else if(N1359) begin
      btb_q[685] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[684] <= 1'b0;
    end else if(N1359) begin
      btb_q[684] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[683] <= 1'b0;
    end else if(N1359) begin
      btb_q[683] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[682] <= 1'b0;
    end else if(N1359) begin
      btb_q[682] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[681] <= 1'b0;
    end else if(N1359) begin
      btb_q[681] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[680] <= 1'b0;
    end else if(N1359) begin
      btb_q[680] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[679] <= 1'b0;
    end else if(N1359) begin
      btb_q[679] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[678] <= 1'b0;
    end else if(N1359) begin
      btb_q[678] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[677] <= 1'b0;
    end else if(N1359) begin
      btb_q[677] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[676] <= 1'b0;
    end else if(N1359) begin
      btb_q[676] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[675] <= 1'b0;
    end else if(N1359) begin
      btb_q[675] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[674] <= 1'b0;
    end else if(N1359) begin
      btb_q[674] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[673] <= 1'b0;
    end else if(N1359) begin
      btb_q[673] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[672] <= 1'b0;
    end else if(N1359) begin
      btb_q[672] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[671] <= 1'b0;
    end else if(N1359) begin
      btb_q[671] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[670] <= 1'b0;
    end else if(N1359) begin
      btb_q[670] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[669] <= 1'b0;
    end else if(N1359) begin
      btb_q[669] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[668] <= 1'b0;
    end else if(N1359) begin
      btb_q[668] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[667] <= 1'b0;
    end else if(N1359) begin
      btb_q[667] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[666] <= 1'b0;
    end else if(N1359) begin
      btb_q[666] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[665] <= 1'b0;
    end else if(N1359) begin
      btb_q[665] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[664] <= 1'b0;
    end else if(N1359) begin
      btb_q[664] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[663] <= 1'b0;
    end else if(N1359) begin
      btb_q[663] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[662] <= 1'b0;
    end else if(N1359) begin
      btb_q[662] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[661] <= 1'b0;
    end else if(N1359) begin
      btb_q[661] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[660] <= 1'b0;
    end else if(N1359) begin
      btb_q[660] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[659] <= 1'b0;
    end else if(N1359) begin
      btb_q[659] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[658] <= 1'b0;
    end else if(N1359) begin
      btb_q[658] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[657] <= 1'b0;
    end else if(N1359) begin
      btb_q[657] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[656] <= 1'b0;
    end else if(N1359) begin
      btb_q[656] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[655] <= 1'b0;
    end else if(N1359) begin
      btb_q[655] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[654] <= 1'b0;
    end else if(N1359) begin
      btb_q[654] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[653] <= 1'b0;
    end else if(N1359) begin
      btb_q[653] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[652] <= 1'b0;
    end else if(N1359) begin
      btb_q[652] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[651] <= 1'b0;
    end else if(N1359) begin
      btb_q[651] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[650] <= 1'b0;
    end else if(N1359) begin
      btb_q[650] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[649] <= 1'b0;
    end else if(N1360) begin
      btb_q[649] <= N539;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[648] <= 1'b0;
    end else if(N1364) begin
      btb_q[648] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[647] <= 1'b0;
    end else if(N1364) begin
      btb_q[647] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[646] <= 1'b0;
    end else if(N1364) begin
      btb_q[646] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[645] <= 1'b0;
    end else if(N1364) begin
      btb_q[645] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[644] <= 1'b0;
    end else if(N1364) begin
      btb_q[644] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[643] <= 1'b0;
    end else if(N1364) begin
      btb_q[643] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[642] <= 1'b0;
    end else if(N1364) begin
      btb_q[642] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[641] <= 1'b0;
    end else if(N1364) begin
      btb_q[641] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[640] <= 1'b0;
    end else if(N1364) begin
      btb_q[640] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[639] <= 1'b0;
    end else if(N1365) begin
      btb_q[639] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[638] <= 1'b0;
    end else if(N1365) begin
      btb_q[638] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[637] <= 1'b0;
    end else if(N1365) begin
      btb_q[637] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[636] <= 1'b0;
    end else if(N1365) begin
      btb_q[636] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[635] <= 1'b0;
    end else if(N1365) begin
      btb_q[635] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[634] <= 1'b0;
    end else if(N1365) begin
      btb_q[634] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[633] <= 1'b0;
    end else if(N1365) begin
      btb_q[633] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[632] <= 1'b0;
    end else if(N1365) begin
      btb_q[632] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[631] <= 1'b0;
    end else if(N1365) begin
      btb_q[631] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[630] <= 1'b0;
    end else if(N1365) begin
      btb_q[630] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[629] <= 1'b0;
    end else if(N1365) begin
      btb_q[629] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[628] <= 1'b0;
    end else if(N1365) begin
      btb_q[628] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[627] <= 1'b0;
    end else if(N1365) begin
      btb_q[627] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[626] <= 1'b0;
    end else if(N1365) begin
      btb_q[626] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[625] <= 1'b0;
    end else if(N1365) begin
      btb_q[625] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[624] <= 1'b0;
    end else if(N1365) begin
      btb_q[624] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[623] <= 1'b0;
    end else if(N1365) begin
      btb_q[623] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[622] <= 1'b0;
    end else if(N1365) begin
      btb_q[622] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[621] <= 1'b0;
    end else if(N1365) begin
      btb_q[621] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[620] <= 1'b0;
    end else if(N1365) begin
      btb_q[620] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[619] <= 1'b0;
    end else if(N1365) begin
      btb_q[619] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[618] <= 1'b0;
    end else if(N1365) begin
      btb_q[618] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[617] <= 1'b0;
    end else if(N1365) begin
      btb_q[617] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[616] <= 1'b0;
    end else if(N1365) begin
      btb_q[616] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[615] <= 1'b0;
    end else if(N1365) begin
      btb_q[615] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[614] <= 1'b0;
    end else if(N1365) begin
      btb_q[614] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[613] <= 1'b0;
    end else if(N1365) begin
      btb_q[613] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[612] <= 1'b0;
    end else if(N1365) begin
      btb_q[612] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[611] <= 1'b0;
    end else if(N1365) begin
      btb_q[611] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[610] <= 1'b0;
    end else if(N1365) begin
      btb_q[610] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[609] <= 1'b0;
    end else if(N1365) begin
      btb_q[609] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[608] <= 1'b0;
    end else if(N1365) begin
      btb_q[608] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[607] <= 1'b0;
    end else if(N1365) begin
      btb_q[607] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[606] <= 1'b0;
    end else if(N1365) begin
      btb_q[606] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[605] <= 1'b0;
    end else if(N1365) begin
      btb_q[605] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[604] <= 1'b0;
    end else if(N1365) begin
      btb_q[604] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[603] <= 1'b0;
    end else if(N1365) begin
      btb_q[603] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[602] <= 1'b0;
    end else if(N1369) begin
      btb_q[602] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[601] <= 1'b0;
    end else if(N1369) begin
      btb_q[601] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[600] <= 1'b0;
    end else if(N1369) begin
      btb_q[600] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[599] <= 1'b0;
    end else if(N1369) begin
      btb_q[599] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[598] <= 1'b0;
    end else if(N1369) begin
      btb_q[598] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[597] <= 1'b0;
    end else if(N1369) begin
      btb_q[597] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[596] <= 1'b0;
    end else if(N1369) begin
      btb_q[596] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[595] <= 1'b0;
    end else if(N1369) begin
      btb_q[595] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[594] <= 1'b0;
    end else if(N1369) begin
      btb_q[594] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[593] <= 1'b0;
    end else if(N1372) begin
      btb_q[593] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[592] <= 1'b0;
    end else if(N1372) begin
      btb_q[592] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[591] <= 1'b0;
    end else if(N1372) begin
      btb_q[591] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[590] <= 1'b0;
    end else if(N1372) begin
      btb_q[590] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[589] <= 1'b0;
    end else if(N1372) begin
      btb_q[589] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[588] <= 1'b0;
    end else if(N1372) begin
      btb_q[588] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[587] <= 1'b0;
    end else if(N1372) begin
      btb_q[587] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[586] <= 1'b0;
    end else if(N1372) begin
      btb_q[586] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[585] <= 1'b0;
    end else if(N1372) begin
      btb_q[585] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[584] <= 1'b0;
    end else if(N1373) begin
      btb_q[584] <= N538;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[583] <= 1'b0;
    end else if(N1377) begin
      btb_q[583] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[582] <= 1'b0;
    end else if(N1377) begin
      btb_q[582] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[581] <= 1'b0;
    end else if(N1377) begin
      btb_q[581] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[580] <= 1'b0;
    end else if(N1377) begin
      btb_q[580] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[579] <= 1'b0;
    end else if(N1377) begin
      btb_q[579] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[578] <= 1'b0;
    end else if(N1377) begin
      btb_q[578] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[577] <= 1'b0;
    end else if(N1377) begin
      btb_q[577] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[576] <= 1'b0;
    end else if(N1377) begin
      btb_q[576] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[575] <= 1'b0;
    end else if(N1377) begin
      btb_q[575] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[574] <= 1'b0;
    end else if(N1377) begin
      btb_q[574] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[573] <= 1'b0;
    end else if(N1377) begin
      btb_q[573] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[572] <= 1'b0;
    end else if(N1377) begin
      btb_q[572] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[571] <= 1'b0;
    end else if(N1377) begin
      btb_q[571] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[570] <= 1'b0;
    end else if(N1377) begin
      btb_q[570] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[569] <= 1'b0;
    end else if(N1377) begin
      btb_q[569] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[568] <= 1'b0;
    end else if(N1377) begin
      btb_q[568] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[567] <= 1'b0;
    end else if(N1377) begin
      btb_q[567] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[566] <= 1'b0;
    end else if(N1377) begin
      btb_q[566] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[565] <= 1'b0;
    end else if(N1377) begin
      btb_q[565] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[564] <= 1'b0;
    end else if(N1377) begin
      btb_q[564] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[563] <= 1'b0;
    end else if(N1377) begin
      btb_q[563] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[562] <= 1'b0;
    end else if(N1377) begin
      btb_q[562] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[561] <= 1'b0;
    end else if(N1377) begin
      btb_q[561] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[560] <= 1'b0;
    end else if(N1377) begin
      btb_q[560] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[559] <= 1'b0;
    end else if(N1377) begin
      btb_q[559] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[558] <= 1'b0;
    end else if(N1377) begin
      btb_q[558] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[557] <= 1'b0;
    end else if(N1377) begin
      btb_q[557] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[556] <= 1'b0;
    end else if(N1377) begin
      btb_q[556] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[555] <= 1'b0;
    end else if(N1377) begin
      btb_q[555] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[554] <= 1'b0;
    end else if(N1377) begin
      btb_q[554] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[553] <= 1'b0;
    end else if(N1377) begin
      btb_q[553] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[552] <= 1'b0;
    end else if(N1377) begin
      btb_q[552] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[551] <= 1'b0;
    end else if(N1377) begin
      btb_q[551] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[550] <= 1'b0;
    end else if(N1377) begin
      btb_q[550] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[549] <= 1'b0;
    end else if(N1377) begin
      btb_q[549] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[548] <= 1'b0;
    end else if(N1377) begin
      btb_q[548] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[547] <= 1'b0;
    end else if(N1377) begin
      btb_q[547] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[546] <= 1'b0;
    end else if(N1377) begin
      btb_q[546] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[545] <= 1'b0;
    end else if(N1377) begin
      btb_q[545] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[544] <= 1'b0;
    end else if(N1377) begin
      btb_q[544] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[543] <= 1'b0;
    end else if(N1377) begin
      btb_q[543] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[542] <= 1'b0;
    end else if(N1377) begin
      btb_q[542] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[541] <= 1'b0;
    end else if(N1377) begin
      btb_q[541] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[540] <= 1'b0;
    end else if(N1377) begin
      btb_q[540] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[539] <= 1'b0;
    end else if(N1378) begin
      btb_q[539] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[538] <= 1'b0;
    end else if(N1378) begin
      btb_q[538] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[537] <= 1'b0;
    end else if(N1378) begin
      btb_q[537] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[536] <= 1'b0;
    end else if(N1378) begin
      btb_q[536] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[535] <= 1'b0;
    end else if(N1378) begin
      btb_q[535] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[534] <= 1'b0;
    end else if(N1378) begin
      btb_q[534] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[533] <= 1'b0;
    end else if(N1378) begin
      btb_q[533] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[532] <= 1'b0;
    end else if(N1378) begin
      btb_q[532] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[531] <= 1'b0;
    end else if(N1378) begin
      btb_q[531] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[530] <= 1'b0;
    end else if(N1378) begin
      btb_q[530] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[529] <= 1'b0;
    end else if(N1378) begin
      btb_q[529] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[528] <= 1'b0;
    end else if(N1378) begin
      btb_q[528] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[527] <= 1'b0;
    end else if(N1378) begin
      btb_q[527] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[526] <= 1'b0;
    end else if(N1378) begin
      btb_q[526] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[525] <= 1'b0;
    end else if(N1378) begin
      btb_q[525] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[524] <= 1'b0;
    end else if(N1378) begin
      btb_q[524] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[523] <= 1'b0;
    end else if(N1378) begin
      btb_q[523] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[522] <= 1'b0;
    end else if(N1378) begin
      btb_q[522] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[521] <= 1'b0;
    end else if(N1378) begin
      btb_q[521] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[520] <= 1'b0;
    end else if(N1378) begin
      btb_q[520] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[519] <= 1'b0;
    end else if(N1373) begin
      btb_q[519] <= N537;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[518] <= 1'b0;
    end else if(N1382) begin
      btb_q[518] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[517] <= 1'b0;
    end else if(N1382) begin
      btb_q[517] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[516] <= 1'b0;
    end else if(N1382) begin
      btb_q[516] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[515] <= 1'b0;
    end else if(N1382) begin
      btb_q[515] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[514] <= 1'b0;
    end else if(N1382) begin
      btb_q[514] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[513] <= 1'b0;
    end else if(N1382) begin
      btb_q[513] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[512] <= 1'b0;
    end else if(N1382) begin
      btb_q[512] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[511] <= 1'b0;
    end else if(N1382) begin
      btb_q[511] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[510] <= 1'b0;
    end else if(N1382) begin
      btb_q[510] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[509] <= 1'b0;
    end else if(N1382) begin
      btb_q[509] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[508] <= 1'b0;
    end else if(N1382) begin
      btb_q[508] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[507] <= 1'b0;
    end else if(N1382) begin
      btb_q[507] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[506] <= 1'b0;
    end else if(N1382) begin
      btb_q[506] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[505] <= 1'b0;
    end else if(N1382) begin
      btb_q[505] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[504] <= 1'b0;
    end else if(N1382) begin
      btb_q[504] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[503] <= 1'b0;
    end else if(N1382) begin
      btb_q[503] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[502] <= 1'b0;
    end else if(N1382) begin
      btb_q[502] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[501] <= 1'b0;
    end else if(N1386) begin
      btb_q[501] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[500] <= 1'b0;
    end else if(N1386) begin
      btb_q[500] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[499] <= 1'b0;
    end else if(N1386) begin
      btb_q[499] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[498] <= 1'b0;
    end else if(N1386) begin
      btb_q[498] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[497] <= 1'b0;
    end else if(N1386) begin
      btb_q[497] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[496] <= 1'b0;
    end else if(N1386) begin
      btb_q[496] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[495] <= 1'b0;
    end else if(N1386) begin
      btb_q[495] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[494] <= 1'b0;
    end else if(N1389) begin
      btb_q[494] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[493] <= 1'b0;
    end else if(N1389) begin
      btb_q[493] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[492] <= 1'b0;
    end else if(N1389) begin
      btb_q[492] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[491] <= 1'b0;
    end else if(N1389) begin
      btb_q[491] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[490] <= 1'b0;
    end else if(N1389) begin
      btb_q[490] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[489] <= 1'b0;
    end else if(N1389) begin
      btb_q[489] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[488] <= 1'b0;
    end else if(N1389) begin
      btb_q[488] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[487] <= 1'b0;
    end else if(N1389) begin
      btb_q[487] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[486] <= 1'b0;
    end else if(N1389) begin
      btb_q[486] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[485] <= 1'b0;
    end else if(N1389) begin
      btb_q[485] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[484] <= 1'b0;
    end else if(N1389) begin
      btb_q[484] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[483] <= 1'b0;
    end else if(N1389) begin
      btb_q[483] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[482] <= 1'b0;
    end else if(N1389) begin
      btb_q[482] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[481] <= 1'b0;
    end else if(N1389) begin
      btb_q[481] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[480] <= 1'b0;
    end else if(N1389) begin
      btb_q[480] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[479] <= 1'b0;
    end else if(N1389) begin
      btb_q[479] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[478] <= 1'b0;
    end else if(N1389) begin
      btb_q[478] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[477] <= 1'b0;
    end else if(N1389) begin
      btb_q[477] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[476] <= 1'b0;
    end else if(N1389) begin
      btb_q[476] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[475] <= 1'b0;
    end else if(N1389) begin
      btb_q[475] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[474] <= 1'b0;
    end else if(N1389) begin
      btb_q[474] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[473] <= 1'b0;
    end else if(N1389) begin
      btb_q[473] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[472] <= 1'b0;
    end else if(N1389) begin
      btb_q[472] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[471] <= 1'b0;
    end else if(N1389) begin
      btb_q[471] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[470] <= 1'b0;
    end else if(N1389) begin
      btb_q[470] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[469] <= 1'b0;
    end else if(N1389) begin
      btb_q[469] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[468] <= 1'b0;
    end else if(N1389) begin
      btb_q[468] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[467] <= 1'b0;
    end else if(N1389) begin
      btb_q[467] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[466] <= 1'b0;
    end else if(N1389) begin
      btb_q[466] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[465] <= 1'b0;
    end else if(N1389) begin
      btb_q[465] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[464] <= 1'b0;
    end else if(N1389) begin
      btb_q[464] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[463] <= 1'b0;
    end else if(N1389) begin
      btb_q[463] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[462] <= 1'b0;
    end else if(N1389) begin
      btb_q[462] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[461] <= 1'b0;
    end else if(N1389) begin
      btb_q[461] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[460] <= 1'b0;
    end else if(N1389) begin
      btb_q[460] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[459] <= 1'b0;
    end else if(N1389) begin
      btb_q[459] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[458] <= 1'b0;
    end else if(N1389) begin
      btb_q[458] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[457] <= 1'b0;
    end else if(N1389) begin
      btb_q[457] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[456] <= 1'b0;
    end else if(N1389) begin
      btb_q[456] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[455] <= 1'b0;
    end else if(N1389) begin
      btb_q[455] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[454] <= 1'b0;
    end else if(N1390) begin
      btb_q[454] <= N536;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[453] <= 1'b0;
    end else if(N1394) begin
      btb_q[453] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[452] <= 1'b0;
    end else if(N1394) begin
      btb_q[452] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[451] <= 1'b0;
    end else if(N1394) begin
      btb_q[451] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[450] <= 1'b0;
    end else if(N1394) begin
      btb_q[450] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[449] <= 1'b0;
    end else if(N1394) begin
      btb_q[449] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[448] <= 1'b0;
    end else if(N1394) begin
      btb_q[448] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[447] <= 1'b0;
    end else if(N1394) begin
      btb_q[447] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[446] <= 1'b0;
    end else if(N1394) begin
      btb_q[446] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[445] <= 1'b0;
    end else if(N1394) begin
      btb_q[445] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[444] <= 1'b0;
    end else if(N1394) begin
      btb_q[444] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[443] <= 1'b0;
    end else if(N1394) begin
      btb_q[443] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[442] <= 1'b0;
    end else if(N1394) begin
      btb_q[442] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[441] <= 1'b0;
    end else if(N1394) begin
      btb_q[441] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[440] <= 1'b0;
    end else if(N1394) begin
      btb_q[440] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[439] <= 1'b0;
    end else if(N1394) begin
      btb_q[439] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[438] <= 1'b0;
    end else if(N1395) begin
      btb_q[438] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[437] <= 1'b0;
    end else if(N1395) begin
      btb_q[437] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[436] <= 1'b0;
    end else if(N1395) begin
      btb_q[436] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[435] <= 1'b0;
    end else if(N1395) begin
      btb_q[435] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[434] <= 1'b0;
    end else if(N1395) begin
      btb_q[434] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[433] <= 1'b0;
    end else if(N1395) begin
      btb_q[433] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[432] <= 1'b0;
    end else if(N1395) begin
      btb_q[432] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[431] <= 1'b0;
    end else if(N1395) begin
      btb_q[431] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[430] <= 1'b0;
    end else if(N1395) begin
      btb_q[430] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[429] <= 1'b0;
    end else if(N1395) begin
      btb_q[429] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[428] <= 1'b0;
    end else if(N1395) begin
      btb_q[428] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[427] <= 1'b0;
    end else if(N1395) begin
      btb_q[427] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[426] <= 1'b0;
    end else if(N1395) begin
      btb_q[426] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[425] <= 1'b0;
    end else if(N1395) begin
      btb_q[425] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[424] <= 1'b0;
    end else if(N1395) begin
      btb_q[424] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[423] <= 1'b0;
    end else if(N1395) begin
      btb_q[423] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[422] <= 1'b0;
    end else if(N1395) begin
      btb_q[422] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[421] <= 1'b0;
    end else if(N1395) begin
      btb_q[421] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[420] <= 1'b0;
    end else if(N1395) begin
      btb_q[420] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[419] <= 1'b0;
    end else if(N1395) begin
      btb_q[419] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[418] <= 1'b0;
    end else if(N1395) begin
      btb_q[418] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[417] <= 1'b0;
    end else if(N1395) begin
      btb_q[417] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[416] <= 1'b0;
    end else if(N1395) begin
      btb_q[416] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[415] <= 1'b0;
    end else if(N1395) begin
      btb_q[415] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[414] <= 1'b0;
    end else if(N1395) begin
      btb_q[414] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[413] <= 1'b0;
    end else if(N1395) begin
      btb_q[413] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[412] <= 1'b0;
    end else if(N1395) begin
      btb_q[412] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[411] <= 1'b0;
    end else if(N1395) begin
      btb_q[411] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[410] <= 1'b0;
    end else if(N1395) begin
      btb_q[410] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[409] <= 1'b0;
    end else if(N1395) begin
      btb_q[409] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[408] <= 1'b0;
    end else if(N1395) begin
      btb_q[408] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[407] <= 1'b0;
    end else if(N1395) begin
      btb_q[407] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[406] <= 1'b0;
    end else if(N1395) begin
      btb_q[406] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[405] <= 1'b0;
    end else if(N1395) begin
      btb_q[405] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[404] <= 1'b0;
    end else if(N1395) begin
      btb_q[404] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[403] <= 1'b0;
    end else if(N1395) begin
      btb_q[403] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[402] <= 1'b0;
    end else if(N1395) begin
      btb_q[402] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[401] <= 1'b0;
    end else if(N1399) begin
      btb_q[401] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[400] <= 1'b0;
    end else if(N1399) begin
      btb_q[400] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[399] <= 1'b0;
    end else if(N1399) begin
      btb_q[399] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[398] <= 1'b0;
    end else if(N1399) begin
      btb_q[398] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[397] <= 1'b0;
    end else if(N1399) begin
      btb_q[397] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[396] <= 1'b0;
    end else if(N1399) begin
      btb_q[396] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[395] <= 1'b0;
    end else if(N1402) begin
      btb_q[395] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[394] <= 1'b0;
    end else if(N1402) begin
      btb_q[394] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[393] <= 1'b0;
    end else if(N1402) begin
      btb_q[393] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[392] <= 1'b0;
    end else if(N1402) begin
      btb_q[392] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[391] <= 1'b0;
    end else if(N1402) begin
      btb_q[391] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[390] <= 1'b0;
    end else if(N1402) begin
      btb_q[390] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[389] <= 1'b0;
    end else if(N1403) begin
      btb_q[389] <= N535;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[388] <= 1'b0;
    end else if(N1407) begin
      btb_q[388] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[387] <= 1'b0;
    end else if(N1407) begin
      btb_q[387] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[386] <= 1'b0;
    end else if(N1407) begin
      btb_q[386] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[385] <= 1'b0;
    end else if(N1407) begin
      btb_q[385] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[384] <= 1'b0;
    end else if(N1407) begin
      btb_q[384] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[383] <= 1'b0;
    end else if(N1407) begin
      btb_q[383] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[382] <= 1'b0;
    end else if(N1407) begin
      btb_q[382] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[381] <= 1'b0;
    end else if(N1407) begin
      btb_q[381] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[380] <= 1'b0;
    end else if(N1407) begin
      btb_q[380] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[379] <= 1'b0;
    end else if(N1407) begin
      btb_q[379] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[378] <= 1'b0;
    end else if(N1407) begin
      btb_q[378] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[377] <= 1'b0;
    end else if(N1407) begin
      btb_q[377] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[376] <= 1'b0;
    end else if(N1407) begin
      btb_q[376] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[375] <= 1'b0;
    end else if(N1407) begin
      btb_q[375] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[374] <= 1'b0;
    end else if(N1407) begin
      btb_q[374] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[373] <= 1'b0;
    end else if(N1407) begin
      btb_q[373] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[372] <= 1'b0;
    end else if(N1407) begin
      btb_q[372] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[371] <= 1'b0;
    end else if(N1407) begin
      btb_q[371] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[370] <= 1'b0;
    end else if(N1407) begin
      btb_q[370] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[369] <= 1'b0;
    end else if(N1407) begin
      btb_q[369] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[368] <= 1'b0;
    end else if(N1407) begin
      btb_q[368] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[367] <= 1'b0;
    end else if(N1407) begin
      btb_q[367] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[366] <= 1'b0;
    end else if(N1407) begin
      btb_q[366] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[365] <= 1'b0;
    end else if(N1407) begin
      btb_q[365] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[364] <= 1'b0;
    end else if(N1407) begin
      btb_q[364] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[363] <= 1'b0;
    end else if(N1407) begin
      btb_q[363] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[362] <= 1'b0;
    end else if(N1407) begin
      btb_q[362] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[361] <= 1'b0;
    end else if(N1407) begin
      btb_q[361] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[360] <= 1'b0;
    end else if(N1407) begin
      btb_q[360] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[359] <= 1'b0;
    end else if(N1407) begin
      btb_q[359] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[358] <= 1'b0;
    end else if(N1407) begin
      btb_q[358] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[357] <= 1'b0;
    end else if(N1407) begin
      btb_q[357] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[356] <= 1'b0;
    end else if(N1407) begin
      btb_q[356] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[355] <= 1'b0;
    end else if(N1407) begin
      btb_q[355] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[354] <= 1'b0;
    end else if(N1407) begin
      btb_q[354] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[353] <= 1'b0;
    end else if(N1407) begin
      btb_q[353] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[352] <= 1'b0;
    end else if(N1407) begin
      btb_q[352] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[351] <= 1'b0;
    end else if(N1407) begin
      btb_q[351] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[350] <= 1'b0;
    end else if(N1407) begin
      btb_q[350] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[349] <= 1'b0;
    end else if(N1407) begin
      btb_q[349] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[348] <= 1'b0;
    end else if(N1407) begin
      btb_q[348] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[347] <= 1'b0;
    end else if(N1407) begin
      btb_q[347] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[346] <= 1'b0;
    end else if(N1407) begin
      btb_q[346] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[345] <= 1'b0;
    end else if(N1407) begin
      btb_q[345] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[344] <= 1'b0;
    end else if(N1407) begin
      btb_q[344] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[343] <= 1'b0;
    end else if(N1407) begin
      btb_q[343] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[342] <= 1'b0;
    end else if(N1407) begin
      btb_q[342] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[341] <= 1'b0;
    end else if(N1407) begin
      btb_q[341] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[340] <= 1'b0;
    end else if(N1407) begin
      btb_q[340] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[339] <= 1'b0;
    end else if(N1407) begin
      btb_q[339] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[338] <= 1'b0;
    end else if(N1408) begin
      btb_q[338] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[337] <= 1'b0;
    end else if(N1408) begin
      btb_q[337] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[336] <= 1'b0;
    end else if(N1408) begin
      btb_q[336] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[335] <= 1'b0;
    end else if(N1408) begin
      btb_q[335] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[334] <= 1'b0;
    end else if(N1408) begin
      btb_q[334] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[333] <= 1'b0;
    end else if(N1408) begin
      btb_q[333] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[332] <= 1'b0;
    end else if(N1408) begin
      btb_q[332] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[331] <= 1'b0;
    end else if(N1408) begin
      btb_q[331] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[330] <= 1'b0;
    end else if(N1408) begin
      btb_q[330] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[329] <= 1'b0;
    end else if(N1408) begin
      btb_q[329] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[328] <= 1'b0;
    end else if(N1408) begin
      btb_q[328] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[327] <= 1'b0;
    end else if(N1408) begin
      btb_q[327] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[326] <= 1'b0;
    end else if(N1408) begin
      btb_q[326] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[325] <= 1'b0;
    end else if(N1408) begin
      btb_q[325] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[324] <= 1'b0;
    end else if(N1403) begin
      btb_q[324] <= N534;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[323] <= 1'b0;
    end else if(N1412) begin
      btb_q[323] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[322] <= 1'b0;
    end else if(N1412) begin
      btb_q[322] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[321] <= 1'b0;
    end else if(N1412) begin
      btb_q[321] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[320] <= 1'b0;
    end else if(N1412) begin
      btb_q[320] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[319] <= 1'b0;
    end else if(N1412) begin
      btb_q[319] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[318] <= 1'b0;
    end else if(N1412) begin
      btb_q[318] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[317] <= 1'b0;
    end else if(N1412) begin
      btb_q[317] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[316] <= 1'b0;
    end else if(N1412) begin
      btb_q[316] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[315] <= 1'b0;
    end else if(N1412) begin
      btb_q[315] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[314] <= 1'b0;
    end else if(N1412) begin
      btb_q[314] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[313] <= 1'b0;
    end else if(N1412) begin
      btb_q[313] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[312] <= 1'b0;
    end else if(N1412) begin
      btb_q[312] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[311] <= 1'b0;
    end else if(N1412) begin
      btb_q[311] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[310] <= 1'b0;
    end else if(N1412) begin
      btb_q[310] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[309] <= 1'b0;
    end else if(N1412) begin
      btb_q[309] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[308] <= 1'b0;
    end else if(N1412) begin
      btb_q[308] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[307] <= 1'b0;
    end else if(N1412) begin
      btb_q[307] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[306] <= 1'b0;
    end else if(N1412) begin
      btb_q[306] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[305] <= 1'b0;
    end else if(N1412) begin
      btb_q[305] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[304] <= 1'b0;
    end else if(N1412) begin
      btb_q[304] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[303] <= 1'b0;
    end else if(N1412) begin
      btb_q[303] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[302] <= 1'b0;
    end else if(N1412) begin
      btb_q[302] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[301] <= 1'b0;
    end else if(N1412) begin
      btb_q[301] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[300] <= 1'b0;
    end else if(N1416) begin
      btb_q[300] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[299] <= 1'b0;
    end else if(N1416) begin
      btb_q[299] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[298] <= 1'b0;
    end else if(N1416) begin
      btb_q[298] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[297] <= 1'b0;
    end else if(N1416) begin
      btb_q[297] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[296] <= 1'b0;
    end else if(N1419) begin
      btb_q[296] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[295] <= 1'b0;
    end else if(N1419) begin
      btb_q[295] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[294] <= 1'b0;
    end else if(N1419) begin
      btb_q[294] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[293] <= 1'b0;
    end else if(N1419) begin
      btb_q[293] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[292] <= 1'b0;
    end else if(N1419) begin
      btb_q[292] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[291] <= 1'b0;
    end else if(N1419) begin
      btb_q[291] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[290] <= 1'b0;
    end else if(N1419) begin
      btb_q[290] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[289] <= 1'b0;
    end else if(N1419) begin
      btb_q[289] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[288] <= 1'b0;
    end else if(N1419) begin
      btb_q[288] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[287] <= 1'b0;
    end else if(N1419) begin
      btb_q[287] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[286] <= 1'b0;
    end else if(N1419) begin
      btb_q[286] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[285] <= 1'b0;
    end else if(N1419) begin
      btb_q[285] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[284] <= 1'b0;
    end else if(N1419) begin
      btb_q[284] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[283] <= 1'b0;
    end else if(N1419) begin
      btb_q[283] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[282] <= 1'b0;
    end else if(N1419) begin
      btb_q[282] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[281] <= 1'b0;
    end else if(N1419) begin
      btb_q[281] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[280] <= 1'b0;
    end else if(N1419) begin
      btb_q[280] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[279] <= 1'b0;
    end else if(N1419) begin
      btb_q[279] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[278] <= 1'b0;
    end else if(N1419) begin
      btb_q[278] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[277] <= 1'b0;
    end else if(N1419) begin
      btb_q[277] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[276] <= 1'b0;
    end else if(N1419) begin
      btb_q[276] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[275] <= 1'b0;
    end else if(N1419) begin
      btb_q[275] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[274] <= 1'b0;
    end else if(N1419) begin
      btb_q[274] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[273] <= 1'b0;
    end else if(N1419) begin
      btb_q[273] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[272] <= 1'b0;
    end else if(N1419) begin
      btb_q[272] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[271] <= 1'b0;
    end else if(N1419) begin
      btb_q[271] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[270] <= 1'b0;
    end else if(N1419) begin
      btb_q[270] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[269] <= 1'b0;
    end else if(N1419) begin
      btb_q[269] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[268] <= 1'b0;
    end else if(N1419) begin
      btb_q[268] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[267] <= 1'b0;
    end else if(N1419) begin
      btb_q[267] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[266] <= 1'b0;
    end else if(N1419) begin
      btb_q[266] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[265] <= 1'b0;
    end else if(N1419) begin
      btb_q[265] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[264] <= 1'b0;
    end else if(N1419) begin
      btb_q[264] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[263] <= 1'b0;
    end else if(N1419) begin
      btb_q[263] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[262] <= 1'b0;
    end else if(N1419) begin
      btb_q[262] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[261] <= 1'b0;
    end else if(N1419) begin
      btb_q[261] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[260] <= 1'b0;
    end else if(N1419) begin
      btb_q[260] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[259] <= 1'b0;
    end else if(N1420) begin
      btb_q[259] <= N533;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[258] <= 1'b0;
    end else if(N1424) begin
      btb_q[258] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[257] <= 1'b0;
    end else if(N1424) begin
      btb_q[257] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[256] <= 1'b0;
    end else if(N1424) begin
      btb_q[256] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[255] <= 1'b0;
    end else if(N1424) begin
      btb_q[255] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[254] <= 1'b0;
    end else if(N1424) begin
      btb_q[254] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[253] <= 1'b0;
    end else if(N1424) begin
      btb_q[253] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[252] <= 1'b0;
    end else if(N1424) begin
      btb_q[252] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[251] <= 1'b0;
    end else if(N1424) begin
      btb_q[251] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[250] <= 1'b0;
    end else if(N1424) begin
      btb_q[250] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[249] <= 1'b0;
    end else if(N1424) begin
      btb_q[249] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[248] <= 1'b0;
    end else if(N1424) begin
      btb_q[248] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[247] <= 1'b0;
    end else if(N1424) begin
      btb_q[247] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[246] <= 1'b0;
    end else if(N1424) begin
      btb_q[246] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[245] <= 1'b0;
    end else if(N1424) begin
      btb_q[245] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[244] <= 1'b0;
    end else if(N1424) begin
      btb_q[244] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[243] <= 1'b0;
    end else if(N1424) begin
      btb_q[243] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[242] <= 1'b0;
    end else if(N1424) begin
      btb_q[242] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[241] <= 1'b0;
    end else if(N1424) begin
      btb_q[241] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[240] <= 1'b0;
    end else if(N1424) begin
      btb_q[240] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[239] <= 1'b0;
    end else if(N1424) begin
      btb_q[239] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[238] <= 1'b0;
    end else if(N1424) begin
      btb_q[238] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[237] <= 1'b0;
    end else if(N1425) begin
      btb_q[237] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[236] <= 1'b0;
    end else if(N1425) begin
      btb_q[236] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[235] <= 1'b0;
    end else if(N1425) begin
      btb_q[235] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[234] <= 1'b0;
    end else if(N1425) begin
      btb_q[234] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[233] <= 1'b0;
    end else if(N1425) begin
      btb_q[233] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[232] <= 1'b0;
    end else if(N1425) begin
      btb_q[232] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[231] <= 1'b0;
    end else if(N1425) begin
      btb_q[231] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[230] <= 1'b0;
    end else if(N1425) begin
      btb_q[230] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[229] <= 1'b0;
    end else if(N1425) begin
      btb_q[229] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[228] <= 1'b0;
    end else if(N1425) begin
      btb_q[228] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[227] <= 1'b0;
    end else if(N1425) begin
      btb_q[227] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[226] <= 1'b0;
    end else if(N1425) begin
      btb_q[226] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[225] <= 1'b0;
    end else if(N1425) begin
      btb_q[225] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[224] <= 1'b0;
    end else if(N1425) begin
      btb_q[224] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[223] <= 1'b0;
    end else if(N1425) begin
      btb_q[223] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[222] <= 1'b0;
    end else if(N1425) begin
      btb_q[222] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[221] <= 1'b0;
    end else if(N1425) begin
      btb_q[221] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[220] <= 1'b0;
    end else if(N1425) begin
      btb_q[220] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[219] <= 1'b0;
    end else if(N1425) begin
      btb_q[219] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[218] <= 1'b0;
    end else if(N1425) begin
      btb_q[218] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[217] <= 1'b0;
    end else if(N1425) begin
      btb_q[217] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[216] <= 1'b0;
    end else if(N1425) begin
      btb_q[216] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[215] <= 1'b0;
    end else if(N1425) begin
      btb_q[215] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[214] <= 1'b0;
    end else if(N1425) begin
      btb_q[214] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[213] <= 1'b0;
    end else if(N1425) begin
      btb_q[213] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[212] <= 1'b0;
    end else if(N1425) begin
      btb_q[212] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[211] <= 1'b0;
    end else if(N1425) begin
      btb_q[211] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[210] <= 1'b0;
    end else if(N1425) begin
      btb_q[210] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[209] <= 1'b0;
    end else if(N1425) begin
      btb_q[209] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[208] <= 1'b0;
    end else if(N1425) begin
      btb_q[208] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[207] <= 1'b0;
    end else if(N1425) begin
      btb_q[207] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[206] <= 1'b0;
    end else if(N1425) begin
      btb_q[206] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[205] <= 1'b0;
    end else if(N1425) begin
      btb_q[205] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[204] <= 1'b0;
    end else if(N1425) begin
      btb_q[204] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[203] <= 1'b0;
    end else if(N1425) begin
      btb_q[203] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[202] <= 1'b0;
    end else if(N1425) begin
      btb_q[202] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[201] <= 1'b0;
    end else if(N1425) begin
      btb_q[201] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[200] <= 1'b0;
    end else if(N1429) begin
      btb_q[200] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[199] <= 1'b0;
    end else if(N1429) begin
      btb_q[199] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[198] <= 1'b0;
    end else if(N1429) begin
      btb_q[198] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[197] <= 1'b0;
    end else if(N1432) begin
      btb_q[197] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[196] <= 1'b0;
    end else if(N1432) begin
      btb_q[196] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[195] <= 1'b0;
    end else if(N1432) begin
      btb_q[195] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[194] <= 1'b0;
    end else if(N1433) begin
      btb_q[194] <= N532;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[193] <= 1'b0;
    end else if(N1437) begin
      btb_q[193] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[192] <= 1'b0;
    end else if(N1437) begin
      btb_q[192] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[191] <= 1'b0;
    end else if(N1437) begin
      btb_q[191] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[190] <= 1'b0;
    end else if(N1437) begin
      btb_q[190] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[189] <= 1'b0;
    end else if(N1437) begin
      btb_q[189] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[188] <= 1'b0;
    end else if(N1437) begin
      btb_q[188] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[187] <= 1'b0;
    end else if(N1437) begin
      btb_q[187] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[186] <= 1'b0;
    end else if(N1437) begin
      btb_q[186] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[185] <= 1'b0;
    end else if(N1437) begin
      btb_q[185] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[184] <= 1'b0;
    end else if(N1437) begin
      btb_q[184] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[183] <= 1'b0;
    end else if(N1437) begin
      btb_q[183] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[182] <= 1'b0;
    end else if(N1437) begin
      btb_q[182] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[181] <= 1'b0;
    end else if(N1437) begin
      btb_q[181] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[180] <= 1'b0;
    end else if(N1437) begin
      btb_q[180] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[179] <= 1'b0;
    end else if(N1437) begin
      btb_q[179] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[178] <= 1'b0;
    end else if(N1437) begin
      btb_q[178] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[177] <= 1'b0;
    end else if(N1437) begin
      btb_q[177] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[176] <= 1'b0;
    end else if(N1437) begin
      btb_q[176] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[175] <= 1'b0;
    end else if(N1437) begin
      btb_q[175] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[174] <= 1'b0;
    end else if(N1437) begin
      btb_q[174] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[173] <= 1'b0;
    end else if(N1437) begin
      btb_q[173] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[172] <= 1'b0;
    end else if(N1437) begin
      btb_q[172] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[171] <= 1'b0;
    end else if(N1437) begin
      btb_q[171] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[170] <= 1'b0;
    end else if(N1437) begin
      btb_q[170] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[169] <= 1'b0;
    end else if(N1437) begin
      btb_q[169] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[168] <= 1'b0;
    end else if(N1437) begin
      btb_q[168] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[167] <= 1'b0;
    end else if(N1437) begin
      btb_q[167] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[166] <= 1'b0;
    end else if(N1437) begin
      btb_q[166] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[165] <= 1'b0;
    end else if(N1437) begin
      btb_q[165] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[164] <= 1'b0;
    end else if(N1437) begin
      btb_q[164] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[163] <= 1'b0;
    end else if(N1437) begin
      btb_q[163] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[162] <= 1'b0;
    end else if(N1437) begin
      btb_q[162] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[161] <= 1'b0;
    end else if(N1437) begin
      btb_q[161] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[160] <= 1'b0;
    end else if(N1437) begin
      btb_q[160] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[159] <= 1'b0;
    end else if(N1437) begin
      btb_q[159] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[158] <= 1'b0;
    end else if(N1437) begin
      btb_q[158] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[157] <= 1'b0;
    end else if(N1437) begin
      btb_q[157] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[156] <= 1'b0;
    end else if(N1437) begin
      btb_q[156] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[155] <= 1'b0;
    end else if(N1437) begin
      btb_q[155] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[154] <= 1'b0;
    end else if(N1437) begin
      btb_q[154] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[153] <= 1'b0;
    end else if(N1437) begin
      btb_q[153] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[152] <= 1'b0;
    end else if(N1437) begin
      btb_q[152] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[151] <= 1'b0;
    end else if(N1437) begin
      btb_q[151] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[150] <= 1'b0;
    end else if(N1437) begin
      btb_q[150] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[149] <= 1'b0;
    end else if(N1437) begin
      btb_q[149] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[148] <= 1'b0;
    end else if(N1437) begin
      btb_q[148] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[147] <= 1'b0;
    end else if(N1437) begin
      btb_q[147] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[146] <= 1'b0;
    end else if(N1437) begin
      btb_q[146] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[145] <= 1'b0;
    end else if(N1437) begin
      btb_q[145] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[144] <= 1'b0;
    end else if(N1437) begin
      btb_q[144] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[143] <= 1'b0;
    end else if(N1437) begin
      btb_q[143] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[142] <= 1'b0;
    end else if(N1437) begin
      btb_q[142] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[141] <= 1'b0;
    end else if(N1437) begin
      btb_q[141] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[140] <= 1'b0;
    end else if(N1437) begin
      btb_q[140] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[139] <= 1'b0;
    end else if(N1437) begin
      btb_q[139] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[138] <= 1'b0;
    end else if(N1437) begin
      btb_q[138] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[137] <= 1'b0;
    end else if(N1438) begin
      btb_q[137] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[136] <= 1'b0;
    end else if(N1438) begin
      btb_q[136] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[135] <= 1'b0;
    end else if(N1438) begin
      btb_q[135] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[134] <= 1'b0;
    end else if(N1438) begin
      btb_q[134] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[133] <= 1'b0;
    end else if(N1438) begin
      btb_q[133] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[132] <= 1'b0;
    end else if(N1438) begin
      btb_q[132] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[131] <= 1'b0;
    end else if(N1438) begin
      btb_q[131] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[130] <= 1'b0;
    end else if(N1438) begin
      btb_q[130] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[129] <= 1'b0;
    end else if(N1433) begin
      btb_q[129] <= N531;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[128] <= 1'b0;
    end else if(N1442) begin
      btb_q[128] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[127] <= 1'b0;
    end else if(N1442) begin
      btb_q[127] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[126] <= 1'b0;
    end else if(N1442) begin
      btb_q[126] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[125] <= 1'b0;
    end else if(N1442) begin
      btb_q[125] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[124] <= 1'b0;
    end else if(N1442) begin
      btb_q[124] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[123] <= 1'b0;
    end else if(N1442) begin
      btb_q[123] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[122] <= 1'b0;
    end else if(N1442) begin
      btb_q[122] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[121] <= 1'b0;
    end else if(N1442) begin
      btb_q[121] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[120] <= 1'b0;
    end else if(N1442) begin
      btb_q[120] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[119] <= 1'b0;
    end else if(N1442) begin
      btb_q[119] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[118] <= 1'b0;
    end else if(N1442) begin
      btb_q[118] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[117] <= 1'b0;
    end else if(N1442) begin
      btb_q[117] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[116] <= 1'b0;
    end else if(N1442) begin
      btb_q[116] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[115] <= 1'b0;
    end else if(N1442) begin
      btb_q[115] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[114] <= 1'b0;
    end else if(N1442) begin
      btb_q[114] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[113] <= 1'b0;
    end else if(N1442) begin
      btb_q[113] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[112] <= 1'b0;
    end else if(N1442) begin
      btb_q[112] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[111] <= 1'b0;
    end else if(N1442) begin
      btb_q[111] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[110] <= 1'b0;
    end else if(N1442) begin
      btb_q[110] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[109] <= 1'b0;
    end else if(N1442) begin
      btb_q[109] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[108] <= 1'b0;
    end else if(N1442) begin
      btb_q[108] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[107] <= 1'b0;
    end else if(N1442) begin
      btb_q[107] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[106] <= 1'b0;
    end else if(N1442) begin
      btb_q[106] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[105] <= 1'b0;
    end else if(N1442) begin
      btb_q[105] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[104] <= 1'b0;
    end else if(N1442) begin
      btb_q[104] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[103] <= 1'b0;
    end else if(N1442) begin
      btb_q[103] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[102] <= 1'b0;
    end else if(N1442) begin
      btb_q[102] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[101] <= 1'b0;
    end else if(N1442) begin
      btb_q[101] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[100] <= 1'b0;
    end else if(N1442) begin
      btb_q[100] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[99] <= 1'b0;
    end else if(N1446) begin
      btb_q[99] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[98] <= 1'b0;
    end else if(N1449) begin
      btb_q[98] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[97] <= 1'b0;
    end else if(N1449) begin
      btb_q[97] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[96] <= 1'b0;
    end else if(N1449) begin
      btb_q[96] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[95] <= 1'b0;
    end else if(N1449) begin
      btb_q[95] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[94] <= 1'b0;
    end else if(N1449) begin
      btb_q[94] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[93] <= 1'b0;
    end else if(N1449) begin
      btb_q[93] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[92] <= 1'b0;
    end else if(N1449) begin
      btb_q[92] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[91] <= 1'b0;
    end else if(N1449) begin
      btb_q[91] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[90] <= 1'b0;
    end else if(N1449) begin
      btb_q[90] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[89] <= 1'b0;
    end else if(N1449) begin
      btb_q[89] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[88] <= 1'b0;
    end else if(N1449) begin
      btb_q[88] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[87] <= 1'b0;
    end else if(N1449) begin
      btb_q[87] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[86] <= 1'b0;
    end else if(N1449) begin
      btb_q[86] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[85] <= 1'b0;
    end else if(N1449) begin
      btb_q[85] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[84] <= 1'b0;
    end else if(N1449) begin
      btb_q[84] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[83] <= 1'b0;
    end else if(N1449) begin
      btb_q[83] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[82] <= 1'b0;
    end else if(N1449) begin
      btb_q[82] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[81] <= 1'b0;
    end else if(N1449) begin
      btb_q[81] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[80] <= 1'b0;
    end else if(N1449) begin
      btb_q[80] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[79] <= 1'b0;
    end else if(N1449) begin
      btb_q[79] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[78] <= 1'b0;
    end else if(N1449) begin
      btb_q[78] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[77] <= 1'b0;
    end else if(N1449) begin
      btb_q[77] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[76] <= 1'b0;
    end else if(N1449) begin
      btb_q[76] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[75] <= 1'b0;
    end else if(N1449) begin
      btb_q[75] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[74] <= 1'b0;
    end else if(N1449) begin
      btb_q[74] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[73] <= 1'b0;
    end else if(N1449) begin
      btb_q[73] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[72] <= 1'b0;
    end else if(N1449) begin
      btb_q[72] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[71] <= 1'b0;
    end else if(N1449) begin
      btb_q[71] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[70] <= 1'b0;
    end else if(N1449) begin
      btb_q[70] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[69] <= 1'b0;
    end else if(N1449) begin
      btb_q[69] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[68] <= 1'b0;
    end else if(N1449) begin
      btb_q[68] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[67] <= 1'b0;
    end else if(N1449) begin
      btb_q[67] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[66] <= 1'b0;
    end else if(N1449) begin
      btb_q[66] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[65] <= 1'b0;
    end else if(N1449) begin
      btb_q[65] <= btb_update_i[1];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[64] <= 1'b0;
    end else if(N595) begin
      btb_q[64] <= N530;
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[63] <= 1'b0;
    end else if(N1453) begin
      btb_q[63] <= btb_update_i[64];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[62] <= 1'b0;
    end else if(N1453) begin
      btb_q[62] <= btb_update_i[63];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[61] <= 1'b0;
    end else if(N1453) begin
      btb_q[61] <= btb_update_i[62];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[60] <= 1'b0;
    end else if(N1453) begin
      btb_q[60] <= btb_update_i[61];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[59] <= 1'b0;
    end else if(N1453) begin
      btb_q[59] <= btb_update_i[60];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[58] <= 1'b0;
    end else if(N1453) begin
      btb_q[58] <= btb_update_i[59];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[57] <= 1'b0;
    end else if(N1453) begin
      btb_q[57] <= btb_update_i[58];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[56] <= 1'b0;
    end else if(N1453) begin
      btb_q[56] <= btb_update_i[57];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[55] <= 1'b0;
    end else if(N1453) begin
      btb_q[55] <= btb_update_i[56];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[54] <= 1'b0;
    end else if(N1453) begin
      btb_q[54] <= btb_update_i[55];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[53] <= 1'b0;
    end else if(N1453) begin
      btb_q[53] <= btb_update_i[54];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[52] <= 1'b0;
    end else if(N1453) begin
      btb_q[52] <= btb_update_i[53];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[51] <= 1'b0;
    end else if(N1453) begin
      btb_q[51] <= btb_update_i[52];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[50] <= 1'b0;
    end else if(N1453) begin
      btb_q[50] <= btb_update_i[51];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[49] <= 1'b0;
    end else if(N1453) begin
      btb_q[49] <= btb_update_i[50];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[48] <= 1'b0;
    end else if(N1453) begin
      btb_q[48] <= btb_update_i[49];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[47] <= 1'b0;
    end else if(N1453) begin
      btb_q[47] <= btb_update_i[48];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[46] <= 1'b0;
    end else if(N1453) begin
      btb_q[46] <= btb_update_i[47];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[45] <= 1'b0;
    end else if(N1453) begin
      btb_q[45] <= btb_update_i[46];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[44] <= 1'b0;
    end else if(N1453) begin
      btb_q[44] <= btb_update_i[45];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[43] <= 1'b0;
    end else if(N1453) begin
      btb_q[43] <= btb_update_i[44];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[42] <= 1'b0;
    end else if(N1453) begin
      btb_q[42] <= btb_update_i[43];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[41] <= 1'b0;
    end else if(N1453) begin
      btb_q[41] <= btb_update_i[42];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[40] <= 1'b0;
    end else if(N1453) begin
      btb_q[40] <= btb_update_i[41];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[39] <= 1'b0;
    end else if(N1454) begin
      btb_q[39] <= btb_update_i[40];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[38] <= 1'b0;
    end else if(N1455) begin
      btb_q[38] <= btb_update_i[39];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[37] <= 1'b0;
    end else if(N1456) begin
      btb_q[37] <= btb_update_i[38];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[36] <= 1'b0;
    end else if(N1457) begin
      btb_q[36] <= btb_update_i[37];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[35] <= 1'b0;
    end else if(N1458) begin
      btb_q[35] <= btb_update_i[36];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[34] <= 1'b0;
    end else if(N1459) begin
      btb_q[34] <= btb_update_i[35];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[33] <= 1'b0;
    end else if(N1460) begin
      btb_q[33] <= btb_update_i[34];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[32] <= 1'b0;
    end else if(N1461) begin
      btb_q[32] <= btb_update_i[33];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[31] <= 1'b0;
    end else if(N1462) begin
      btb_q[31] <= btb_update_i[32];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[30] <= 1'b0;
    end else if(N1463) begin
      btb_q[30] <= btb_update_i[31];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[29] <= 1'b0;
    end else if(N1464) begin
      btb_q[29] <= btb_update_i[30];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[28] <= 1'b0;
    end else if(N1465) begin
      btb_q[28] <= btb_update_i[29];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[27] <= 1'b0;
    end else if(N1466) begin
      btb_q[27] <= btb_update_i[28];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[26] <= 1'b0;
    end else if(N1467) begin
      btb_q[26] <= btb_update_i[27];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[25] <= 1'b0;
    end else if(N1468) begin
      btb_q[25] <= btb_update_i[26];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[24] <= 1'b0;
    end else if(N1469) begin
      btb_q[24] <= btb_update_i[25];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[23] <= 1'b0;
    end else if(N1470) begin
      btb_q[23] <= btb_update_i[24];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[22] <= 1'b0;
    end else if(N1471) begin
      btb_q[22] <= btb_update_i[23];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[21] <= 1'b0;
    end else if(N1472) begin
      btb_q[21] <= btb_update_i[22];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[20] <= 1'b0;
    end else if(N1473) begin
      btb_q[20] <= btb_update_i[21];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[19] <= 1'b0;
    end else if(N1474) begin
      btb_q[19] <= btb_update_i[20];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[18] <= 1'b0;
    end else if(N1475) begin
      btb_q[18] <= btb_update_i[19];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[17] <= 1'b0;
    end else if(N1476) begin
      btb_q[17] <= btb_update_i[18];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[16] <= 1'b0;
    end else if(N1477) begin
      btb_q[16] <= btb_update_i[17];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[15] <= 1'b0;
    end else if(N1478) begin
      btb_q[15] <= btb_update_i[16];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[14] <= 1'b0;
    end else if(N1479) begin
      btb_q[14] <= btb_update_i[15];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[13] <= 1'b0;
    end else if(N1480) begin
      btb_q[13] <= btb_update_i[14];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[12] <= 1'b0;
    end else if(N1481) begin
      btb_q[12] <= btb_update_i[13];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[11] <= 1'b0;
    end else if(N1482) begin
      btb_q[11] <= btb_update_i[12];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[10] <= 1'b0;
    end else if(N1483) begin
      btb_q[10] <= btb_update_i[11];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[9] <= 1'b0;
    end else if(N1484) begin
      btb_q[9] <= btb_update_i[10];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[8] <= 1'b0;
    end else if(N1485) begin
      btb_q[8] <= btb_update_i[9];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[7] <= 1'b0;
    end else if(N1486) begin
      btb_q[7] <= btb_update_i[8];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[6] <= 1'b0;
    end else if(N1487) begin
      btb_q[6] <= btb_update_i[7];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[5] <= 1'b0;
    end else if(N1488) begin
      btb_q[5] <= btb_update_i[6];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[4] <= 1'b0;
    end else if(N1489) begin
      btb_q[4] <= btb_update_i[5];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[3] <= 1'b0;
    end else if(N1490) begin
      btb_q[3] <= btb_update_i[4];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[2] <= 1'b0;
    end else if(N1491) begin
      btb_q[2] <= btb_update_i[3];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[1] <= 1'b0;
    end else if(N1492) begin
      btb_q[1] <= btb_update_i[2];
    end 
  end


  always @(posedge clk_i or posedge N528) begin
    if(N528) begin
      btb_q[0] <= 1'b0;
    end else if(N1493) begin
      btb_q[0] <= btb_update_i[1];
    end 
  end

  assign N1494 = ~btb_update_i[71];
  assign N1495 = btb_update_i[69] & btb_update_i[70];
  assign N1496 = N0 & btb_update_i[70];
  assign N0 = ~btb_update_i[69];
  assign N1497 = btb_update_i[69] & N1;
  assign N1 = ~btb_update_i[70];
  assign N1498 = N2 & N3;
  assign N2 = ~btb_update_i[69];
  assign N3 = ~btb_update_i[70];
  assign N1499 = btb_update_i[71] & N1495;
  assign N1500 = btb_update_i[71] & N1496;
  assign N1501 = btb_update_i[71] & N1497;
  assign N1502 = btb_update_i[71] & N1498;
  assign N1503 = N1494 & N1495;
  assign N1504 = N1494 & N1496;
  assign N1505 = N1494 & N1497;
  assign N1506 = N1494 & N1498;
  assign N1507 = ~btb_update_i[68];
  assign N1508 = btb_update_i[66] & btb_update_i[67];
  assign N1509 = N4 & btb_update_i[67];
  assign N4 = ~btb_update_i[66];
  assign N1510 = btb_update_i[66] & N5;
  assign N5 = ~btb_update_i[67];
  assign N1511 = N6 & N7;
  assign N6 = ~btb_update_i[66];
  assign N7 = ~btb_update_i[67];
  assign N1512 = btb_update_i[68] & N1508;
  assign N1513 = btb_update_i[68] & N1509;
  assign N1514 = btb_update_i[68] & N1510;
  assign N1515 = btb_update_i[68] & N1511;
  assign N1516 = N1507 & N1508;
  assign N1517 = N1507 & N1509;
  assign N1518 = N1507 & N1510;
  assign N1519 = N1507 & N1511;
  assign N335 = N1499 & N1512;
  assign N334 = N1499 & N1513;
  assign N333 = N1499 & N1514;
  assign N332 = N1499 & N1515;
  assign N331 = N1499 & N1516;
  assign N330 = N1499 & N1517;
  assign N329 = N1499 & N1518;
  assign N328 = N1499 & N1519;
  assign N327 = N1500 & N1512;
  assign N326 = N1500 & N1513;
  assign N325 = N1500 & N1514;
  assign N324 = N1500 & N1515;
  assign N323 = N1500 & N1516;
  assign N322 = N1500 & N1517;
  assign N321 = N1500 & N1518;
  assign N320 = N1500 & N1519;
  assign N319 = N1501 & N1512;
  assign N318 = N1501 & N1513;
  assign N317 = N1501 & N1514;
  assign N316 = N1501 & N1515;
  assign N315 = N1501 & N1516;
  assign N314 = N1501 & N1517;
  assign N313 = N1501 & N1518;
  assign N312 = N1501 & N1519;
  assign N311 = N1502 & N1512;
  assign N310 = N1502 & N1513;
  assign N309 = N1502 & N1514;
  assign N308 = N1502 & N1515;
  assign N307 = N1502 & N1516;
  assign N306 = N1502 & N1517;
  assign N305 = N1502 & N1518;
  assign N304 = N1502 & N1519;
  assign N303 = N1503 & N1512;
  assign N302 = N1503 & N1513;
  assign N301 = N1503 & N1514;
  assign N300 = N1503 & N1515;
  assign N299 = N1503 & N1516;
  assign N298 = N1503 & N1517;
  assign N297 = N1503 & N1518;
  assign N296 = N1503 & N1519;
  assign N295 = N1504 & N1512;
  assign N294 = N1504 & N1513;
  assign N293 = N1504 & N1514;
  assign N292 = N1504 & N1515;
  assign N291 = N1504 & N1516;
  assign N290 = N1504 & N1517;
  assign N289 = N1504 & N1518;
  assign N288 = N1504 & N1519;
  assign N287 = N1505 & N1512;
  assign N286 = N1505 & N1513;
  assign N285 = N1505 & N1514;
  assign N284 = N1505 & N1515;
  assign N283 = N1505 & N1516;
  assign N282 = N1505 & N1517;
  assign N281 = N1505 & N1518;
  assign N280 = N1505 & N1519;
  assign N279 = N1506 & N1512;
  assign N278 = N1506 & N1513;
  assign N277 = N1506 & N1514;
  assign N276 = N1506 & N1515;
  assign N275 = N1506 & N1516;
  assign N274 = N1506 & N1517;
  assign N273 = N1506 & N1518;
  assign N272 = N1506 & N1519;
  assign N207 = (N8)? 1'b1 : 
                (N336)? btb_q[64] : 1'b0;
  assign N8 = N272;
  assign N208 = (N9)? 1'b1 : 
                (N338)? btb_q[129] : 1'b0;
  assign N9 = N273;
  assign N209 = (N10)? 1'b1 : 
                (N340)? btb_q[194] : 1'b0;
  assign N10 = N274;
  assign N210 = (N11)? 1'b1 : 
                (N342)? btb_q[259] : 1'b0;
  assign N11 = N275;
  assign N211 = (N12)? 1'b1 : 
                (N344)? btb_q[324] : 1'b0;
  assign N12 = N276;
  assign N212 = (N13)? 1'b1 : 
                (N346)? btb_q[389] : 1'b0;
  assign N13 = N277;
  assign N213 = (N14)? 1'b1 : 
                (N348)? btb_q[454] : 1'b0;
  assign N14 = N278;
  assign N214 = (N15)? 1'b1 : 
                (N350)? btb_q[519] : 1'b0;
  assign N15 = N279;
  assign N215 = (N16)? 1'b1 : 
                (N352)? btb_q[584] : 1'b0;
  assign N16 = N280;
  assign N216 = (N17)? 1'b1 : 
                (N354)? btb_q[649] : 1'b0;
  assign N17 = N281;
  assign N217 = (N18)? 1'b1 : 
                (N356)? btb_q[714] : 1'b0;
  assign N18 = N282;
  assign N218 = (N19)? 1'b1 : 
                (N358)? btb_q[779] : 1'b0;
  assign N19 = N283;
  assign N219 = (N20)? 1'b1 : 
                (N360)? btb_q[844] : 1'b0;
  assign N20 = N284;
  assign N220 = (N21)? 1'b1 : 
                (N362)? btb_q[909] : 1'b0;
  assign N21 = N285;
  assign N221 = (N22)? 1'b1 : 
                (N364)? btb_q[974] : 1'b0;
  assign N22 = N286;
  assign N222 = (N23)? 1'b1 : 
                (N366)? btb_q[1039] : 1'b0;
  assign N23 = N287;
  assign N223 = (N24)? 1'b1 : 
                (N368)? btb_q[1104] : 1'b0;
  assign N24 = N288;
  assign N224 = (N25)? 1'b1 : 
                (N370)? btb_q[1169] : 1'b0;
  assign N25 = N289;
  assign N225 = (N26)? 1'b1 : 
                (N372)? btb_q[1234] : 1'b0;
  assign N26 = N290;
  assign N226 = (N27)? 1'b1 : 
                (N374)? btb_q[1299] : 1'b0;
  assign N27 = N291;
  assign N227 = (N28)? 1'b1 : 
                (N376)? btb_q[1364] : 1'b0;
  assign N28 = N292;
  assign N228 = (N29)? 1'b1 : 
                (N378)? btb_q[1429] : 1'b0;
  assign N29 = N293;
  assign N229 = (N30)? 1'b1 : 
                (N380)? btb_q[1494] : 1'b0;
  assign N30 = N294;
  assign N230 = (N31)? 1'b1 : 
                (N382)? btb_q[1559] : 1'b0;
  assign N31 = N295;
  assign N231 = (N32)? 1'b1 : 
                (N384)? btb_q[1624] : 1'b0;
  assign N32 = N296;
  assign N232 = (N33)? 1'b1 : 
                (N386)? btb_q[1689] : 1'b0;
  assign N33 = N297;
  assign N233 = (N34)? 1'b1 : 
                (N388)? btb_q[1754] : 1'b0;
  assign N34 = N298;
  assign N234 = (N35)? 1'b1 : 
                (N390)? btb_q[1819] : 1'b0;
  assign N35 = N299;
  assign N235 = (N36)? 1'b1 : 
                (N392)? btb_q[1884] : 1'b0;
  assign N36 = N300;
  assign N236 = (N37)? 1'b1 : 
                (N394)? btb_q[1949] : 1'b0;
  assign N37 = N301;
  assign N237 = (N38)? 1'b1 : 
                (N396)? btb_q[2014] : 1'b0;
  assign N38 = N302;
  assign N238 = (N39)? 1'b1 : 
                (N398)? btb_q[2079] : 1'b0;
  assign N39 = N303;
  assign N239 = (N40)? 1'b1 : 
                (N400)? btb_q[2144] : 1'b0;
  assign N40 = N304;
  assign N240 = (N41)? 1'b1 : 
                (N402)? btb_q[2209] : 1'b0;
  assign N41 = N305;
  assign N241 = (N42)? 1'b1 : 
                (N404)? btb_q[2274] : 1'b0;
  assign N42 = N306;
  assign N242 = (N43)? 1'b1 : 
                (N406)? btb_q[2339] : 1'b0;
  assign N43 = N307;
  assign N243 = (N44)? 1'b1 : 
                (N408)? btb_q[2404] : 1'b0;
  assign N44 = N308;
  assign N244 = (N45)? 1'b1 : 
                (N410)? btb_q[2469] : 1'b0;
  assign N45 = N309;
  assign N245 = (N46)? 1'b1 : 
                (N412)? btb_q[2534] : 1'b0;
  assign N46 = N310;
  assign N246 = (N47)? 1'b1 : 
                (N414)? btb_q[2599] : 1'b0;
  assign N47 = N311;
  assign N247 = (N48)? 1'b1 : 
                (N416)? btb_q[2664] : 1'b0;
  assign N48 = N312;
  assign N248 = (N49)? 1'b1 : 
                (N418)? btb_q[2729] : 1'b0;
  assign N49 = N313;
  assign N249 = (N50)? 1'b1 : 
                (N420)? btb_q[2794] : 1'b0;
  assign N50 = N314;
  assign N250 = (N51)? 1'b1 : 
                (N422)? btb_q[2859] : 1'b0;
  assign N51 = N315;
  assign N251 = (N52)? 1'b1 : 
                (N424)? btb_q[2924] : 1'b0;
  assign N52 = N316;
  assign N252 = (N53)? 1'b1 : 
                (N426)? btb_q[2989] : 1'b0;
  assign N53 = N317;
  assign N253 = (N54)? 1'b1 : 
                (N428)? btb_q[3054] : 1'b0;
  assign N54 = N318;
  assign N254 = (N55)? 1'b1 : 
                (N430)? btb_q[3119] : 1'b0;
  assign N55 = N319;
  assign N255 = (N56)? 1'b1 : 
                (N432)? btb_q[3184] : 1'b0;
  assign N56 = N320;
  assign N256 = (N57)? 1'b1 : 
                (N434)? btb_q[3249] : 1'b0;
  assign N57 = N321;
  assign N257 = (N58)? 1'b1 : 
                (N436)? btb_q[3314] : 1'b0;
  assign N58 = N322;
  assign N258 = (N59)? 1'b1 : 
                (N438)? btb_q[3379] : 1'b0;
  assign N59 = N323;
  assign N259 = (N60)? 1'b1 : 
                (N440)? btb_q[3444] : 1'b0;
  assign N60 = N324;
  assign N260 = (N61)? 1'b1 : 
                (N442)? btb_q[3509] : 1'b0;
  assign N61 = N325;
  assign N261 = (N62)? 1'b1 : 
                (N444)? btb_q[3574] : 1'b0;
  assign N62 = N326;
  assign N262 = (N63)? 1'b1 : 
                (N446)? btb_q[3639] : 1'b0;
  assign N63 = N327;
  assign N263 = (N64)? 1'b1 : 
                (N448)? btb_q[3704] : 1'b0;
  assign N64 = N328;
  assign N264 = (N65)? 1'b1 : 
                (N450)? btb_q[3769] : 1'b0;
  assign N65 = N329;
  assign N265 = (N66)? 1'b1 : 
                (N452)? btb_q[3834] : 1'b0;
  assign N66 = N330;
  assign N266 = (N67)? 1'b1 : 
                (N454)? btb_q[3899] : 1'b0;
  assign N67 = N331;
  assign N267 = (N68)? 1'b1 : 
                (N456)? btb_q[3964] : 1'b0;
  assign N68 = N332;
  assign N268 = (N69)? 1'b1 : 
                (N458)? btb_q[4029] : 1'b0;
  assign N69 = N333;
  assign N269 = (N70)? 1'b1 : 
                (N460)? btb_q[4094] : 1'b0;
  assign N70 = N334;
  assign N270 = (N71)? 1'b1 : 
                (N462)? btb_q[4159] : 1'b0;
  assign N71 = N335;
  assign N337 = (N8)? 1'b0 : 
                (N336)? N207 : 1'b0;
  assign N339 = (N9)? 1'b0 : 
                (N338)? N208 : 1'b0;
  assign N341 = (N10)? 1'b0 : 
                (N340)? N209 : 1'b0;
  assign N343 = (N11)? 1'b0 : 
                (N342)? N210 : 1'b0;
  assign N345 = (N12)? 1'b0 : 
                (N344)? N211 : 1'b0;
  assign N347 = (N13)? 1'b0 : 
                (N346)? N212 : 1'b0;
  assign N349 = (N14)? 1'b0 : 
                (N348)? N213 : 1'b0;
  assign N351 = (N15)? 1'b0 : 
                (N350)? N214 : 1'b0;
  assign N353 = (N16)? 1'b0 : 
                (N352)? N215 : 1'b0;
  assign N355 = (N17)? 1'b0 : 
                (N354)? N216 : 1'b0;
  assign N357 = (N18)? 1'b0 : 
                (N356)? N217 : 1'b0;
  assign N359 = (N19)? 1'b0 : 
                (N358)? N218 : 1'b0;
  assign N361 = (N20)? 1'b0 : 
                (N360)? N219 : 1'b0;
  assign N363 = (N21)? 1'b0 : 
                (N362)? N220 : 1'b0;
  assign N365 = (N22)? 1'b0 : 
                (N364)? N221 : 1'b0;
  assign N367 = (N23)? 1'b0 : 
                (N366)? N222 : 1'b0;
  assign N369 = (N24)? 1'b0 : 
                (N368)? N223 : 1'b0;
  assign N371 = (N25)? 1'b0 : 
                (N370)? N224 : 1'b0;
  assign N373 = (N26)? 1'b0 : 
                (N372)? N225 : 1'b0;
  assign N375 = (N27)? 1'b0 : 
                (N374)? N226 : 1'b0;
  assign N377 = (N28)? 1'b0 : 
                (N376)? N227 : 1'b0;
  assign N379 = (N29)? 1'b0 : 
                (N378)? N228 : 1'b0;
  assign N381 = (N30)? 1'b0 : 
                (N380)? N229 : 1'b0;
  assign N383 = (N31)? 1'b0 : 
                (N382)? N230 : 1'b0;
  assign N385 = (N32)? 1'b0 : 
                (N384)? N231 : 1'b0;
  assign N387 = (N33)? 1'b0 : 
                (N386)? N232 : 1'b0;
  assign N389 = (N34)? 1'b0 : 
                (N388)? N233 : 1'b0;
  assign N391 = (N35)? 1'b0 : 
                (N390)? N234 : 1'b0;
  assign N393 = (N36)? 1'b0 : 
                (N392)? N235 : 1'b0;
  assign N395 = (N37)? 1'b0 : 
                (N394)? N236 : 1'b0;
  assign N397 = (N38)? 1'b0 : 
                (N396)? N237 : 1'b0;
  assign N399 = (N39)? 1'b0 : 
                (N398)? N238 : 1'b0;
  assign N401 = (N40)? 1'b0 : 
                (N400)? N239 : 1'b0;
  assign N403 = (N41)? 1'b0 : 
                (N402)? N240 : 1'b0;
  assign N405 = (N42)? 1'b0 : 
                (N404)? N241 : 1'b0;
  assign N407 = (N43)? 1'b0 : 
                (N406)? N242 : 1'b0;
  assign N409 = (N44)? 1'b0 : 
                (N408)? N243 : 1'b0;
  assign N411 = (N45)? 1'b0 : 
                (N410)? N244 : 1'b0;
  assign N413 = (N46)? 1'b0 : 
                (N412)? N245 : 1'b0;
  assign N415 = (N47)? 1'b0 : 
                (N414)? N246 : 1'b0;
  assign N417 = (N48)? 1'b0 : 
                (N416)? N247 : 1'b0;
  assign N419 = (N49)? 1'b0 : 
                (N418)? N248 : 1'b0;
  assign N421 = (N50)? 1'b0 : 
                (N420)? N249 : 1'b0;
  assign N423 = (N51)? 1'b0 : 
                (N422)? N250 : 1'b0;
  assign N425 = (N52)? 1'b0 : 
                (N424)? N251 : 1'b0;
  assign N427 = (N53)? 1'b0 : 
                (N426)? N252 : 1'b0;
  assign N429 = (N54)? 1'b0 : 
                (N428)? N253 : 1'b0;
  assign N431 = (N55)? 1'b0 : 
                (N430)? N254 : 1'b0;
  assign N433 = (N56)? 1'b0 : 
                (N432)? N255 : 1'b0;
  assign N435 = (N57)? 1'b0 : 
                (N434)? N256 : 1'b0;
  assign N437 = (N58)? 1'b0 : 
                (N436)? N257 : 1'b0;
  assign N439 = (N59)? 1'b0 : 
                (N438)? N258 : 1'b0;
  assign N441 = (N60)? 1'b0 : 
                (N440)? N259 : 1'b0;
  assign N443 = (N61)? 1'b0 : 
                (N442)? N260 : 1'b0;
  assign N445 = (N62)? 1'b0 : 
                (N444)? N261 : 1'b0;
  assign N447 = (N63)? 1'b0 : 
                (N446)? N262 : 1'b0;
  assign N449 = (N64)? 1'b0 : 
                (N448)? N263 : 1'b0;
  assign N451 = (N65)? 1'b0 : 
                (N450)? N264 : 1'b0;
  assign N453 = (N66)? 1'b0 : 
                (N452)? N265 : 1'b0;
  assign N455 = (N67)? 1'b0 : 
                (N454)? N266 : 1'b0;
  assign N457 = (N68)? 1'b0 : 
                (N456)? N267 : 1'b0;
  assign N459 = (N69)? 1'b0 : 
                (N458)? N268 : 1'b0;
  assign N461 = (N70)? 1'b0 : 
                (N460)? N269 : 1'b0;
  assign N463 = (N71)? 1'b0 : 
                (N462)? N270 : 1'b0;
  assign { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } = (N72)? { N463, N461, N459, N457, N455, N453, N451, N449, N447, N445, N443, N441, N439, N437, N435, N433, N431, N429, N427, N425, N423, N421, N419, N417, N415, N413, N411, N409, N407, N405, N403, N401, N399, N397, N395, N393, N391, N389, N387, N385, N383, N381, N379, N377, N375, N373, N371, N369, N367, N365, N363, N361, N359, N357, N355, N353, N351, N349, N347, N345, N343, N341, N339, N337 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N271)? { N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207 } : 1'b0;
  assign N72 = btb_update_i[0];
  assign { N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530 } = (N73)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N74)? { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } : 1'b0;
  assign N73 = flush_i;
  assign N74 = N529;
  assign N75 = ~vpc_i[1];
  assign N76 = ~vpc_i[2];
  assign N77 = N75 & N76;
  assign N78 = N75 & vpc_i[2];
  assign N79 = vpc_i[1] & N76;
  assign N80 = vpc_i[1] & vpc_i[2];
  assign N81 = ~vpc_i[3];
  assign N82 = N77 & N81;
  assign N83 = N77 & vpc_i[3];
  assign N84 = N79 & N81;
  assign N85 = N79 & vpc_i[3];
  assign N86 = N78 & N81;
  assign N87 = N78 & vpc_i[3];
  assign N88 = N80 & N81;
  assign N89 = N80 & vpc_i[3];
  assign N90 = ~vpc_i[4];
  assign N91 = N82 & N90;
  assign N92 = N82 & vpc_i[4];
  assign N93 = N84 & N90;
  assign N94 = N84 & vpc_i[4];
  assign N95 = N86 & N90;
  assign N96 = N86 & vpc_i[4];
  assign N97 = N88 & N90;
  assign N98 = N88 & vpc_i[4];
  assign N99 = N83 & N90;
  assign N100 = N83 & vpc_i[4];
  assign N101 = N85 & N90;
  assign N102 = N85 & vpc_i[4];
  assign N103 = N87 & N90;
  assign N104 = N87 & vpc_i[4];
  assign N105 = N89 & N90;
  assign N106 = N89 & vpc_i[4];
  assign N107 = ~vpc_i[5];
  assign N108 = N91 & N107;
  assign N109 = N91 & vpc_i[5];
  assign N110 = N93 & N107;
  assign N111 = N93 & vpc_i[5];
  assign N112 = N95 & N107;
  assign N113 = N95 & vpc_i[5];
  assign N114 = N97 & N107;
  assign N115 = N97 & vpc_i[5];
  assign N116 = N99 & N107;
  assign N117 = N99 & vpc_i[5];
  assign N118 = N101 & N107;
  assign N119 = N101 & vpc_i[5];
  assign N120 = N103 & N107;
  assign N121 = N103 & vpc_i[5];
  assign N122 = N105 & N107;
  assign N123 = N105 & vpc_i[5];
  assign N124 = N92 & N107;
  assign N125 = N92 & vpc_i[5];
  assign N126 = N94 & N107;
  assign N127 = N94 & vpc_i[5];
  assign N128 = N96 & N107;
  assign N129 = N96 & vpc_i[5];
  assign N130 = N98 & N107;
  assign N131 = N98 & vpc_i[5];
  assign N132 = N100 & N107;
  assign N133 = N100 & vpc_i[5];
  assign N134 = N102 & N107;
  assign N135 = N102 & vpc_i[5];
  assign N136 = N104 & N107;
  assign N137 = N104 & vpc_i[5];
  assign N138 = N106 & N107;
  assign N139 = N106 & vpc_i[5];
  assign N140 = ~vpc_i[6];
  assign N141 = N108 & N140;
  assign N142 = N108 & vpc_i[6];
  assign N143 = N110 & N140;
  assign N144 = N110 & vpc_i[6];
  assign N145 = N112 & N140;
  assign N146 = N112 & vpc_i[6];
  assign N147 = N114 & N140;
  assign N148 = N114 & vpc_i[6];
  assign N149 = N116 & N140;
  assign N150 = N116 & vpc_i[6];
  assign N151 = N118 & N140;
  assign N152 = N118 & vpc_i[6];
  assign N153 = N120 & N140;
  assign N154 = N120 & vpc_i[6];
  assign N155 = N122 & N140;
  assign N156 = N122 & vpc_i[6];
  assign N157 = N124 & N140;
  assign N158 = N124 & vpc_i[6];
  assign N159 = N126 & N140;
  assign N160 = N126 & vpc_i[6];
  assign N161 = N128 & N140;
  assign N162 = N128 & vpc_i[6];
  assign N163 = N130 & N140;
  assign N164 = N130 & vpc_i[6];
  assign N165 = N132 & N140;
  assign N166 = N132 & vpc_i[6];
  assign N167 = N134 & N140;
  assign N168 = N134 & vpc_i[6];
  assign N169 = N136 & N140;
  assign N170 = N136 & vpc_i[6];
  assign N171 = N138 & N140;
  assign N172 = N138 & vpc_i[6];
  assign N173 = N109 & N140;
  assign N174 = N109 & vpc_i[6];
  assign N175 = N111 & N140;
  assign N176 = N111 & vpc_i[6];
  assign N177 = N113 & N140;
  assign N178 = N113 & vpc_i[6];
  assign N179 = N115 & N140;
  assign N180 = N115 & vpc_i[6];
  assign N181 = N117 & N140;
  assign N182 = N117 & vpc_i[6];
  assign N183 = N119 & N140;
  assign N184 = N119 & vpc_i[6];
  assign N185 = N121 & N140;
  assign N186 = N121 & vpc_i[6];
  assign N187 = N123 & N140;
  assign N188 = N123 & vpc_i[6];
  assign N189 = N125 & N140;
  assign N190 = N125 & vpc_i[6];
  assign N191 = N127 & N140;
  assign N192 = N127 & vpc_i[6];
  assign N193 = N129 & N140;
  assign N194 = N129 & vpc_i[6];
  assign N195 = N131 & N140;
  assign N196 = N131 & vpc_i[6];
  assign N197 = N133 & N140;
  assign N198 = N133 & vpc_i[6];
  assign N199 = N135 & N140;
  assign N200 = N135 & vpc_i[6];
  assign N201 = N137 & N140;
  assign N202 = N137 & vpc_i[6];
  assign N203 = N139 & N140;
  assign N204 = N139 & vpc_i[6];
  assign N205 = btb_update_i[129] & N1520;
  assign N1520 = ~debug_mode_i;
  assign N206 = ~N205;
  assign N271 = ~btb_update_i[0];
  assign N336 = ~N272;
  assign N338 = ~N273;
  assign N340 = ~N274;
  assign N342 = ~N275;
  assign N344 = ~N276;
  assign N346 = ~N277;
  assign N348 = ~N278;
  assign N350 = ~N279;
  assign N352 = ~N280;
  assign N354 = ~N281;
  assign N356 = ~N282;
  assign N358 = ~N283;
  assign N360 = ~N284;
  assign N362 = ~N285;
  assign N364 = ~N286;
  assign N366 = ~N287;
  assign N368 = ~N288;
  assign N370 = ~N289;
  assign N372 = ~N290;
  assign N374 = ~N291;
  assign N376 = ~N292;
  assign N378 = ~N293;
  assign N380 = ~N294;
  assign N382 = ~N295;
  assign N384 = ~N296;
  assign N386 = ~N297;
  assign N388 = ~N298;
  assign N390 = ~N299;
  assign N392 = ~N300;
  assign N394 = ~N301;
  assign N396 = ~N302;
  assign N398 = ~N303;
  assign N400 = ~N304;
  assign N402 = ~N305;
  assign N404 = ~N306;
  assign N406 = ~N307;
  assign N408 = ~N308;
  assign N410 = ~N309;
  assign N412 = ~N310;
  assign N414 = ~N311;
  assign N416 = ~N312;
  assign N418 = ~N313;
  assign N420 = ~N314;
  assign N422 = ~N315;
  assign N424 = ~N316;
  assign N426 = ~N317;
  assign N428 = ~N318;
  assign N430 = ~N319;
  assign N432 = ~N320;
  assign N434 = ~N321;
  assign N436 = ~N322;
  assign N438 = ~N323;
  assign N440 = ~N324;
  assign N442 = ~N325;
  assign N444 = ~N326;
  assign N446 = ~N327;
  assign N448 = ~N328;
  assign N450 = ~N329;
  assign N452 = ~N330;
  assign N454 = ~N331;
  assign N456 = ~N332;
  assign N458 = ~N333;
  assign N460 = ~N334;
  assign N462 = ~N335;
  assign N528 = ~rst_ni;
  assign N529 = ~flush_i;
  assign N594 = N206 & N529;
  assign N595 = ~N594;
  assign N596 = N205 & N529;
  assign N597 = N462 & N596;
  assign N598 = N206 & N529;
  assign N599 = N597 | N598;
  assign N600 = ~N599;
  assign N601 = N529 & N600;
  assign N602 = N205 & N529;
  assign N603 = N462 & N602;
  assign N604 = N206 & N529;
  assign N605 = N603 | N604;
  assign N606 = ~N605;
  assign N607 = N529 & N606;
  assign N608 = N205 & N529;
  assign N609 = N462 & N608;
  assign N610 = N206 & N529;
  assign N611 = N609 | N610;
  assign N612 = ~N611;
  assign N613 = N529 & N612;
  assign N614 = N205 & N529;
  assign N615 = N462 & N614;
  assign N616 = N206 & N529;
  assign N617 = N615 | N616;
  assign N618 = ~N617;
  assign N619 = N529 & N618;
  assign N620 = N205 & N529;
  assign N621 = N462 & N620;
  assign N622 = N206 & N529;
  assign N623 = N621 | N622;
  assign N624 = ~N623;
  assign N625 = N529 & N624;
  assign N626 = N205 & N529;
  assign N627 = N462 & N626;
  assign N628 = N206 & N529;
  assign N629 = N627 | N628;
  assign N630 = ~N629;
  assign N631 = N529 & N630;
  assign N632 = N205 & N529;
  assign N633 = N462 & N632;
  assign N634 = N206 & N529;
  assign N635 = N633 | N634;
  assign N636 = ~N635;
  assign N637 = N529 & N636;
  assign N638 = N205 & N529;
  assign N639 = N462 & N638;
  assign N640 = N206 & N529;
  assign N641 = N639 | N640;
  assign N642 = ~N641;
  assign N643 = N529 & N642;
  assign N644 = N205 & N529;
  assign N645 = N462 & N644;
  assign N646 = N206 & N529;
  assign N647 = N645 | N646;
  assign N648 = ~N647;
  assign N649 = N529 & N648;
  assign N650 = N205 & N529;
  assign N651 = N462 & N650;
  assign N652 = N206 & N529;
  assign N653 = N651 | N652;
  assign N654 = ~N653;
  assign N655 = N529 & N654;
  assign N656 = N205 & N529;
  assign N657 = N462 & N656;
  assign N658 = N206 & N529;
  assign N659 = N657 | N658;
  assign N660 = ~N659;
  assign N661 = N529 & N660;
  assign N662 = N205 & N529;
  assign N663 = N462 & N662;
  assign N664 = N206 & N529;
  assign N665 = N663 | N664;
  assign N666 = ~N665;
  assign N667 = N529 & N666;
  assign N668 = N205 & N529;
  assign N669 = N462 & N668;
  assign N670 = N206 & N529;
  assign N671 = N669 | N670;
  assign N672 = ~N671;
  assign N673 = N529 & N672;
  assign N674 = N205 & N529;
  assign N675 = N462 & N674;
  assign N676 = N206 & N529;
  assign N677 = N675 | N676;
  assign N678 = ~N677;
  assign N679 = N529 & N678;
  assign N680 = N205 & N529;
  assign N681 = N462 & N680;
  assign N682 = N206 & N529;
  assign N683 = N681 | N682;
  assign N684 = ~N683;
  assign N685 = N529 & N684;
  assign N686 = N205 & N529;
  assign N687 = N462 & N686;
  assign N688 = N206 & N529;
  assign N689 = N687 | N688;
  assign N690 = ~N689;
  assign N691 = N529 & N690;
  assign N692 = N205 & N529;
  assign N693 = N462 & N692;
  assign N694 = N206 & N529;
  assign N695 = N693 | N694;
  assign N696 = ~N695;
  assign N697 = N529 & N696;
  assign N698 = N205 & N529;
  assign N699 = N462 & N698;
  assign N700 = N206 & N529;
  assign N701 = N699 | N700;
  assign N702 = ~N701;
  assign N703 = N529 & N702;
  assign N704 = N205 & N529;
  assign N705 = N462 & N704;
  assign N706 = N206 & N529;
  assign N707 = N705 | N706;
  assign N708 = ~N707;
  assign N709 = N529 & N708;
  assign N710 = N205 & N529;
  assign N711 = N462 & N710;
  assign N712 = N206 & N529;
  assign N713 = N711 | N712;
  assign N714 = ~N713;
  assign N715 = N529 & N714;
  assign N716 = N205 & N529;
  assign N717 = N462 & N716;
  assign N718 = N206 & N529;
  assign N719 = N717 | N718;
  assign N720 = ~N719;
  assign N721 = N529 & N720;
  assign N722 = N205 & N529;
  assign N723 = N462 & N722;
  assign N724 = N206 & N529;
  assign N725 = N723 | N724;
  assign N726 = ~N725;
  assign N727 = N529 & N726;
  assign N728 = N205 & N529;
  assign N729 = N462 & N728;
  assign N730 = N206 & N529;
  assign N731 = N729 | N730;
  assign N732 = ~N731;
  assign N733 = N529 & N732;
  assign N734 = N205 & N529;
  assign N735 = N462 & N734;
  assign N736 = N206 & N529;
  assign N737 = N735 | N736;
  assign N738 = ~N737;
  assign N739 = N529 & N738;
  assign N740 = N205 & N529;
  assign N741 = N462 & N740;
  assign N742 = N206 & N529;
  assign N743 = N741 | N742;
  assign N744 = ~N743;
  assign N745 = N529 & N744;
  assign N746 = N205 & N529;
  assign N747 = N462 & N746;
  assign N748 = N206 & N529;
  assign N749 = N747 | N748;
  assign N750 = ~N749;
  assign N751 = N529 & N750;
  assign N752 = N205 & N529;
  assign N753 = N462 & N752;
  assign N754 = N206 & N529;
  assign N755 = N753 | N754;
  assign N756 = ~N755;
  assign N757 = N529 & N756;
  assign N758 = N205 & N529;
  assign N759 = N462 & N758;
  assign N760 = N206 & N529;
  assign N761 = N759 | N760;
  assign N762 = ~N761;
  assign N763 = N529 & N762;
  assign N764 = N205 & N529;
  assign N765 = N462 & N764;
  assign N766 = N206 & N529;
  assign N767 = N765 | N766;
  assign N768 = ~N767;
  assign N769 = N529 & N768;
  assign N770 = N205 & N529;
  assign N771 = N462 & N770;
  assign N772 = N206 & N529;
  assign N773 = N771 | N772;
  assign N774 = ~N773;
  assign N775 = N529 & N774;
  assign N776 = N205 & N529;
  assign N777 = N462 & N776;
  assign N778 = N206 & N529;
  assign N779 = N777 | N778;
  assign N780 = ~N779;
  assign N781 = N529 & N780;
  assign N782 = N205 & N529;
  assign N783 = N462 & N782;
  assign N784 = N206 & N529;
  assign N785 = N783 | N784;
  assign N786 = ~N785;
  assign N787 = N529 & N786;
  assign N788 = N205 & N529;
  assign N789 = N462 & N788;
  assign N790 = N206 & N529;
  assign N791 = N789 | N790;
  assign N792 = ~N791;
  assign N793 = N529 & N792;
  assign N794 = N205 & N529;
  assign N795 = N462 & N794;
  assign N796 = N206 & N529;
  assign N797 = N795 | N796;
  assign N798 = ~N797;
  assign N799 = N529 & N798;
  assign N800 = N205 & N529;
  assign N801 = N462 & N800;
  assign N802 = N206 & N529;
  assign N803 = N801 | N802;
  assign N804 = ~N803;
  assign N805 = N529 & N804;
  assign N806 = N205 & N529;
  assign N807 = N462 & N806;
  assign N808 = N206 & N529;
  assign N809 = N807 | N808;
  assign N810 = ~N809;
  assign N811 = N529 & N810;
  assign N812 = N205 & N529;
  assign N813 = N462 & N812;
  assign N814 = N206 & N529;
  assign N815 = N813 | N814;
  assign N816 = ~N815;
  assign N817 = N529 & N816;
  assign N818 = N205 & N529;
  assign N819 = N462 & N818;
  assign N820 = N206 & N529;
  assign N821 = N819 | N820;
  assign N822 = ~N821;
  assign N823 = N529 & N822;
  assign N824 = N205 & N529;
  assign N825 = N462 & N824;
  assign N826 = N206 & N529;
  assign N827 = N825 | N826;
  assign N828 = ~N827;
  assign N829 = N529 & N828;
  assign N830 = N205 & N529;
  assign N831 = N462 & N830;
  assign N832 = N206 & N529;
  assign N833 = N831 | N832;
  assign N834 = ~N833;
  assign N835 = N529 & N834;
  assign N836 = N205 & N529;
  assign N837 = N462 & N836;
  assign N838 = N206 & N529;
  assign N839 = N837 | N838;
  assign N840 = ~N839;
  assign N841 = N529 & N840;
  assign N842 = ~N838;
  assign N843 = N460 & N836;
  assign N844 = N843 | N838;
  assign N845 = ~N844;
  assign N846 = N529 & N845;
  assign N847 = N843 | N832;
  assign N848 = ~N847;
  assign N849 = N529 & N848;
  assign N850 = ~N832;
  assign N851 = N458 & N836;
  assign N852 = N851 | N832;
  assign N853 = ~N852;
  assign N854 = N529 & N853;
  assign N855 = N458 & N830;
  assign N856 = N855 | N832;
  assign N857 = ~N856;
  assign N858 = N529 & N857;
  assign N859 = N456 & N830;
  assign N860 = N859 | N832;
  assign N861 = ~N860;
  assign N862 = N529 & N861;
  assign N863 = N859 | N826;
  assign N864 = ~N863;
  assign N865 = N529 & N864;
  assign N866 = N529 & N864;
  assign N867 = N456 & N824;
  assign N868 = N867 | N826;
  assign N869 = ~N868;
  assign N870 = N529 & N869;
  assign N871 = ~N826;
  assign N872 = N454 & N824;
  assign N873 = N872 | N826;
  assign N874 = ~N873;
  assign N875 = N529 & N874;
  assign N876 = N872 | N820;
  assign N877 = ~N876;
  assign N878 = N529 & N877;
  assign N879 = N529 & N877;
  assign N880 = ~N820;
  assign N881 = N452 & N824;
  assign N882 = N881 | N820;
  assign N883 = ~N882;
  assign N884 = N529 & N883;
  assign N885 = N452 & N818;
  assign N886 = N885 | N820;
  assign N887 = ~N886;
  assign N888 = N529 & N887;
  assign N889 = N450 & N818;
  assign N890 = N889 | N820;
  assign N891 = ~N890;
  assign N892 = N529 & N891;
  assign N893 = N889 | N814;
  assign N894 = ~N893;
  assign N895 = N529 & N894;
  assign N896 = N529 & N894;
  assign N897 = N450 & N812;
  assign N898 = N897 | N814;
  assign N899 = ~N898;
  assign N900 = N529 & N899;
  assign N901 = ~N814;
  assign N902 = N448 & N812;
  assign N903 = N902 | N814;
  assign N904 = ~N903;
  assign N905 = N529 & N904;
  assign N906 = N902 | N808;
  assign N907 = ~N906;
  assign N908 = N529 & N907;
  assign N909 = N529 & N907;
  assign N910 = ~N808;
  assign N911 = N446 & N812;
  assign N912 = N911 | N808;
  assign N913 = ~N912;
  assign N914 = N529 & N913;
  assign N915 = N446 & N806;
  assign N916 = N915 | N808;
  assign N917 = ~N916;
  assign N918 = N529 & N917;
  assign N919 = N444 & N806;
  assign N920 = N919 | N808;
  assign N921 = ~N920;
  assign N922 = N529 & N921;
  assign N923 = N919 | N802;
  assign N924 = ~N923;
  assign N925 = N529 & N924;
  assign N926 = N529 & N924;
  assign N927 = N444 & N800;
  assign N928 = N927 | N802;
  assign N929 = ~N928;
  assign N930 = N529 & N929;
  assign N931 = ~N802;
  assign N932 = N442 & N800;
  assign N933 = N932 | N802;
  assign N934 = ~N933;
  assign N935 = N529 & N934;
  assign N936 = N932 | N796;
  assign N937 = ~N936;
  assign N938 = N529 & N937;
  assign N939 = N529 & N937;
  assign N940 = ~N796;
  assign N941 = N440 & N800;
  assign N942 = N941 | N796;
  assign N943 = ~N942;
  assign N944 = N529 & N943;
  assign N945 = N440 & N794;
  assign N946 = N945 | N796;
  assign N947 = ~N946;
  assign N948 = N529 & N947;
  assign N949 = N438 & N794;
  assign N950 = N949 | N796;
  assign N951 = ~N950;
  assign N952 = N529 & N951;
  assign N953 = N949 | N790;
  assign N954 = ~N953;
  assign N955 = N529 & N954;
  assign N956 = N529 & N954;
  assign N957 = N438 & N788;
  assign N958 = N957 | N790;
  assign N959 = ~N958;
  assign N960 = N529 & N959;
  assign N961 = ~N790;
  assign N962 = N436 & N788;
  assign N963 = N962 | N790;
  assign N964 = ~N963;
  assign N965 = N529 & N964;
  assign N966 = N962 | N784;
  assign N967 = ~N966;
  assign N968 = N529 & N967;
  assign N969 = N529 & N967;
  assign N970 = ~N784;
  assign N971 = N434 & N788;
  assign N972 = N971 | N784;
  assign N973 = ~N972;
  assign N974 = N529 & N973;
  assign N975 = N434 & N782;
  assign N976 = N975 | N784;
  assign N977 = ~N976;
  assign N978 = N529 & N977;
  assign N979 = N432 & N782;
  assign N980 = N979 | N784;
  assign N981 = ~N980;
  assign N982 = N529 & N981;
  assign N983 = N979 | N778;
  assign N984 = ~N983;
  assign N985 = N529 & N984;
  assign N986 = N529 & N984;
  assign N987 = ~N778;
  assign N988 = N430 & N782;
  assign N989 = N988 | N778;
  assign N990 = ~N989;
  assign N991 = N529 & N990;
  assign N992 = N430 & N776;
  assign N993 = N992 | N778;
  assign N994 = ~N993;
  assign N995 = N529 & N994;
  assign N996 = N992 | N772;
  assign N997 = ~N996;
  assign N998 = N529 & N997;
  assign N999 = ~N772;
  assign N1000 = N428 & N776;
  assign N1001 = N1000 | N772;
  assign N1002 = ~N1001;
  assign N1003 = N529 & N1002;
  assign N1004 = N529 & N1002;
  assign N1005 = N428 & N770;
  assign N1006 = N1005 | N772;
  assign N1007 = ~N1006;
  assign N1008 = N529 & N1007;
  assign N1009 = N426 & N770;
  assign N1010 = N1009 | N772;
  assign N1011 = ~N1010;
  assign N1012 = N529 & N1011;
  assign N1013 = N1009 | N766;
  assign N1014 = ~N1013;
  assign N1015 = N529 & N1014;
  assign N1016 = N529 & N1014;
  assign N1017 = ~N766;
  assign N1018 = N424 & N770;
  assign N1019 = N1018 | N766;
  assign N1020 = ~N1019;
  assign N1021 = N529 & N1020;
  assign N1022 = N424 & N764;
  assign N1023 = N1022 | N766;
  assign N1024 = ~N1023;
  assign N1025 = N529 & N1024;
  assign N1026 = N1022 | N760;
  assign N1027 = ~N1026;
  assign N1028 = N529 & N1027;
  assign N1029 = ~N760;
  assign N1030 = N422 & N764;
  assign N1031 = N1030 | N760;
  assign N1032 = ~N1031;
  assign N1033 = N529 & N1032;
  assign N1034 = N529 & N1032;
  assign N1035 = N422 & N758;
  assign N1036 = N1035 | N760;
  assign N1037 = ~N1036;
  assign N1038 = N529 & N1037;
  assign N1039 = N420 & N758;
  assign N1040 = N1039 | N760;
  assign N1041 = ~N1040;
  assign N1042 = N529 & N1041;
  assign N1043 = N1039 | N754;
  assign N1044 = ~N1043;
  assign N1045 = N529 & N1044;
  assign N1046 = N529 & N1044;
  assign N1047 = ~N754;
  assign N1048 = N418 & N758;
  assign N1049 = N1048 | N754;
  assign N1050 = ~N1049;
  assign N1051 = N529 & N1050;
  assign N1052 = N418 & N752;
  assign N1053 = N1052 | N754;
  assign N1054 = ~N1053;
  assign N1055 = N529 & N1054;
  assign N1056 = N1052 | N748;
  assign N1057 = ~N1056;
  assign N1058 = N529 & N1057;
  assign N1059 = ~N748;
  assign N1060 = N416 & N752;
  assign N1061 = N1060 | N748;
  assign N1062 = ~N1061;
  assign N1063 = N529 & N1062;
  assign N1064 = N529 & N1062;
  assign N1065 = N416 & N746;
  assign N1066 = N1065 | N748;
  assign N1067 = ~N1066;
  assign N1068 = N529 & N1067;
  assign N1069 = N414 & N746;
  assign N1070 = N1069 | N748;
  assign N1071 = ~N1070;
  assign N1072 = N529 & N1071;
  assign N1073 = N1069 | N742;
  assign N1074 = ~N1073;
  assign N1075 = N529 & N1074;
  assign N1076 = N529 & N1074;
  assign N1077 = ~N742;
  assign N1078 = N412 & N746;
  assign N1079 = N1078 | N742;
  assign N1080 = ~N1079;
  assign N1081 = N529 & N1080;
  assign N1082 = N412 & N740;
  assign N1083 = N1082 | N742;
  assign N1084 = ~N1083;
  assign N1085 = N529 & N1084;
  assign N1086 = N1082 | N736;
  assign N1087 = ~N1086;
  assign N1088 = N529 & N1087;
  assign N1089 = ~N736;
  assign N1090 = N410 & N740;
  assign N1091 = N1090 | N736;
  assign N1092 = ~N1091;
  assign N1093 = N529 & N1092;
  assign N1094 = N529 & N1092;
  assign N1095 = N410 & N734;
  assign N1096 = N1095 | N736;
  assign N1097 = ~N1096;
  assign N1098 = N529 & N1097;
  assign N1099 = N408 & N734;
  assign N1100 = N1099 | N736;
  assign N1101 = ~N1100;
  assign N1102 = N529 & N1101;
  assign N1103 = N1099 | N730;
  assign N1104 = ~N1103;
  assign N1105 = N529 & N1104;
  assign N1106 = N529 & N1104;
  assign N1107 = ~N730;
  assign N1108 = N406 & N734;
  assign N1109 = N1108 | N730;
  assign N1110 = ~N1109;
  assign N1111 = N529 & N1110;
  assign N1112 = N406 & N728;
  assign N1113 = N1112 | N730;
  assign N1114 = ~N1113;
  assign N1115 = N529 & N1114;
  assign N1116 = N1112 | N724;
  assign N1117 = ~N1116;
  assign N1118 = N529 & N1117;
  assign N1119 = ~N724;
  assign N1120 = N404 & N728;
  assign N1121 = N1120 | N724;
  assign N1122 = ~N1121;
  assign N1123 = N529 & N1122;
  assign N1124 = N529 & N1122;
  assign N1125 = N404 & N722;
  assign N1126 = N1125 | N724;
  assign N1127 = ~N1126;
  assign N1128 = N529 & N1127;
  assign N1129 = N402 & N722;
  assign N1130 = N1129 | N724;
  assign N1131 = ~N1130;
  assign N1132 = N529 & N1131;
  assign N1133 = N1129 | N718;
  assign N1134 = ~N1133;
  assign N1135 = N529 & N1134;
  assign N1136 = N529 & N1134;
  assign N1137 = ~N718;
  assign N1138 = N400 & N722;
  assign N1139 = N1138 | N718;
  assign N1140 = ~N1139;
  assign N1141 = N529 & N1140;
  assign N1142 = N400 & N716;
  assign N1143 = N1142 | N718;
  assign N1144 = ~N1143;
  assign N1145 = N529 & N1144;
  assign N1146 = N398 & N716;
  assign N1147 = N1146 | N712;
  assign N1148 = ~N1147;
  assign N1149 = N529 & N1148;
  assign N1150 = N529 & N1148;
  assign N1151 = ~N712;
  assign N1152 = N396 & N716;
  assign N1153 = N1152 | N712;
  assign N1154 = ~N1153;
  assign N1155 = N529 & N1154;
  assign N1156 = N396 & N710;
  assign N1157 = N1156 | N712;
  assign N1158 = ~N1157;
  assign N1159 = N529 & N1158;
  assign N1160 = N1156 | N706;
  assign N1161 = ~N1160;
  assign N1162 = N529 & N1161;
  assign N1163 = ~N706;
  assign N1164 = N394 & N710;
  assign N1165 = N1164 | N706;
  assign N1166 = ~N1165;
  assign N1167 = N529 & N1166;
  assign N1168 = N529 & N1166;
  assign N1169 = N394 & N704;
  assign N1170 = N1169 | N706;
  assign N1171 = ~N1170;
  assign N1172 = N529 & N1171;
  assign N1173 = N392 & N704;
  assign N1174 = N1173 | N706;
  assign N1175 = ~N1174;
  assign N1176 = N529 & N1175;
  assign N1177 = N1173 | N700;
  assign N1178 = ~N1177;
  assign N1179 = N529 & N1178;
  assign N1180 = N529 & N1178;
  assign N1181 = ~N700;
  assign N1182 = N390 & N704;
  assign N1183 = N1182 | N700;
  assign N1184 = ~N1183;
  assign N1185 = N529 & N1184;
  assign N1186 = N390 & N698;
  assign N1187 = N1186 | N700;
  assign N1188 = ~N1187;
  assign N1189 = N529 & N1188;
  assign N1190 = N1186 | N694;
  assign N1191 = ~N1190;
  assign N1192 = N529 & N1191;
  assign N1193 = ~N694;
  assign N1194 = N388 & N698;
  assign N1195 = N1194 | N694;
  assign N1196 = ~N1195;
  assign N1197 = N529 & N1196;
  assign N1198 = N529 & N1196;
  assign N1199 = N388 & N692;
  assign N1200 = N1199 | N694;
  assign N1201 = ~N1200;
  assign N1202 = N529 & N1201;
  assign N1203 = N386 & N692;
  assign N1204 = N1203 | N694;
  assign N1205 = ~N1204;
  assign N1206 = N529 & N1205;
  assign N1207 = N1203 | N688;
  assign N1208 = ~N1207;
  assign N1209 = N529 & N1208;
  assign N1210 = N529 & N1208;
  assign N1211 = ~N688;
  assign N1212 = N384 & N692;
  assign N1213 = N1212 | N688;
  assign N1214 = ~N1213;
  assign N1215 = N529 & N1214;
  assign N1216 = N384 & N686;
  assign N1217 = N1216 | N688;
  assign N1218 = ~N1217;
  assign N1219 = N529 & N1218;
  assign N1220 = N1216 | N682;
  assign N1221 = ~N1220;
  assign N1222 = N529 & N1221;
  assign N1223 = ~N682;
  assign N1224 = N382 & N686;
  assign N1225 = N1224 | N682;
  assign N1226 = ~N1225;
  assign N1227 = N529 & N1226;
  assign N1228 = N529 & N1226;
  assign N1229 = N382 & N680;
  assign N1230 = N1229 | N682;
  assign N1231 = ~N1230;
  assign N1232 = N529 & N1231;
  assign N1233 = N380 & N680;
  assign N1234 = N1233 | N682;
  assign N1235 = ~N1234;
  assign N1236 = N529 & N1235;
  assign N1237 = N1233 | N676;
  assign N1238 = ~N1237;
  assign N1239 = N529 & N1238;
  assign N1240 = N529 & N1238;
  assign N1241 = ~N676;
  assign N1242 = N378 & N680;
  assign N1243 = N1242 | N676;
  assign N1244 = ~N1243;
  assign N1245 = N529 & N1244;
  assign N1246 = N378 & N674;
  assign N1247 = N1246 | N676;
  assign N1248 = ~N1247;
  assign N1249 = N529 & N1248;
  assign N1250 = N1246 | N670;
  assign N1251 = ~N1250;
  assign N1252 = N529 & N1251;
  assign N1253 = ~N670;
  assign N1254 = N376 & N674;
  assign N1255 = N1254 | N670;
  assign N1256 = ~N1255;
  assign N1257 = N529 & N1256;
  assign N1258 = N529 & N1256;
  assign N1259 = N376 & N668;
  assign N1260 = N1259 | N670;
  assign N1261 = ~N1260;
  assign N1262 = N529 & N1261;
  assign N1263 = N374 & N668;
  assign N1264 = N1263 | N670;
  assign N1265 = ~N1264;
  assign N1266 = N529 & N1265;
  assign N1267 = N1263 | N664;
  assign N1268 = ~N1267;
  assign N1269 = N529 & N1268;
  assign N1270 = N529 & N1268;
  assign N1271 = ~N664;
  assign N1272 = N372 & N668;
  assign N1273 = N1272 | N664;
  assign N1274 = ~N1273;
  assign N1275 = N529 & N1274;
  assign N1276 = N372 & N662;
  assign N1277 = N1276 | N664;
  assign N1278 = ~N1277;
  assign N1279 = N529 & N1278;
  assign N1280 = N1276 | N658;
  assign N1281 = ~N1280;
  assign N1282 = N529 & N1281;
  assign N1283 = ~N658;
  assign N1284 = N370 & N662;
  assign N1285 = N1284 | N658;
  assign N1286 = ~N1285;
  assign N1287 = N529 & N1286;
  assign N1288 = N529 & N1286;
  assign N1289 = N370 & N656;
  assign N1290 = N1289 | N658;
  assign N1291 = ~N1290;
  assign N1292 = N529 & N1291;
  assign N1293 = N368 & N656;
  assign N1294 = N1293 | N658;
  assign N1295 = ~N1294;
  assign N1296 = N529 & N1295;
  assign N1297 = N1293 | N652;
  assign N1298 = ~N1297;
  assign N1299 = N529 & N1298;
  assign N1300 = N529 & N1298;
  assign N1301 = ~N652;
  assign N1302 = N366 & N656;
  assign N1303 = N1302 | N652;
  assign N1304 = ~N1303;
  assign N1305 = N529 & N1304;
  assign N1306 = N366 & N650;
  assign N1307 = N1306 | N652;
  assign N1308 = ~N1307;
  assign N1309 = N529 & N1308;
  assign N1310 = N1306 | N646;
  assign N1311 = ~N1310;
  assign N1312 = N529 & N1311;
  assign N1313 = ~N646;
  assign N1314 = N364 & N650;
  assign N1315 = N1314 | N646;
  assign N1316 = ~N1315;
  assign N1317 = N529 & N1316;
  assign N1318 = N529 & N1316;
  assign N1319 = N362 & N650;
  assign N1320 = N1319 | N646;
  assign N1321 = ~N1320;
  assign N1322 = N529 & N1321;
  assign N1323 = N362 & N644;
  assign N1324 = N1323 | N646;
  assign N1325 = ~N1324;
  assign N1326 = N529 & N1325;
  assign N1327 = N1323 | N640;
  assign N1328 = ~N1327;
  assign N1329 = N529 & N1328;
  assign N1330 = ~N640;
  assign N1331 = N360 & N644;
  assign N1332 = N1331 | N640;
  assign N1333 = ~N1332;
  assign N1334 = N529 & N1333;
  assign N1335 = N529 & N1333;
  assign N1336 = N360 & N638;
  assign N1337 = N1336 | N640;
  assign N1338 = ~N1337;
  assign N1339 = N529 & N1338;
  assign N1340 = N1336 | N634;
  assign N1341 = ~N1340;
  assign N1342 = N529 & N1341;
  assign N1343 = ~N634;
  assign N1344 = N358 & N638;
  assign N1345 = N1344 | N634;
  assign N1346 = ~N1345;
  assign N1347 = N529 & N1346;
  assign N1348 = N529 & N1346;
  assign N1349 = N356 & N638;
  assign N1350 = N1349 | N634;
  assign N1351 = ~N1350;
  assign N1352 = N529 & N1351;
  assign N1353 = N356 & N632;
  assign N1354 = N1353 | N634;
  assign N1355 = ~N1354;
  assign N1356 = N529 & N1355;
  assign N1357 = N1353 | N628;
  assign N1358 = ~N1357;
  assign N1359 = N529 & N1358;
  assign N1360 = ~N628;
  assign N1361 = N354 & N632;
  assign N1362 = N1361 | N628;
  assign N1363 = ~N1362;
  assign N1364 = N529 & N1363;
  assign N1365 = N529 & N1363;
  assign N1366 = N354 & N626;
  assign N1367 = N1366 | N628;
  assign N1368 = ~N1367;
  assign N1369 = N529 & N1368;
  assign N1370 = N1366 | N622;
  assign N1371 = ~N1370;
  assign N1372 = N529 & N1371;
  assign N1373 = ~N622;
  assign N1374 = N352 & N626;
  assign N1375 = N1374 | N622;
  assign N1376 = ~N1375;
  assign N1377 = N529 & N1376;
  assign N1378 = N529 & N1376;
  assign N1379 = N350 & N626;
  assign N1380 = N1379 | N622;
  assign N1381 = ~N1380;
  assign N1382 = N529 & N1381;
  assign N1383 = N350 & N620;
  assign N1384 = N1383 | N622;
  assign N1385 = ~N1384;
  assign N1386 = N529 & N1385;
  assign N1387 = N1383 | N616;
  assign N1388 = ~N1387;
  assign N1389 = N529 & N1388;
  assign N1390 = ~N616;
  assign N1391 = N348 & N620;
  assign N1392 = N1391 | N616;
  assign N1393 = ~N1392;
  assign N1394 = N529 & N1393;
  assign N1395 = N529 & N1393;
  assign N1396 = N348 & N614;
  assign N1397 = N1396 | N616;
  assign N1398 = ~N1397;
  assign N1399 = N529 & N1398;
  assign N1400 = N1396 | N610;
  assign N1401 = ~N1400;
  assign N1402 = N529 & N1401;
  assign N1403 = ~N610;
  assign N1404 = N346 & N614;
  assign N1405 = N1404 | N610;
  assign N1406 = ~N1405;
  assign N1407 = N529 & N1406;
  assign N1408 = N529 & N1406;
  assign N1409 = N344 & N614;
  assign N1410 = N1409 | N610;
  assign N1411 = ~N1410;
  assign N1412 = N529 & N1411;
  assign N1413 = N344 & N608;
  assign N1414 = N1413 | N610;
  assign N1415 = ~N1414;
  assign N1416 = N529 & N1415;
  assign N1417 = N1413 | N604;
  assign N1418 = ~N1417;
  assign N1419 = N529 & N1418;
  assign N1420 = ~N604;
  assign N1421 = N342 & N608;
  assign N1422 = N1421 | N604;
  assign N1423 = ~N1422;
  assign N1424 = N529 & N1423;
  assign N1425 = N529 & N1423;
  assign N1426 = N342 & N602;
  assign N1427 = N1426 | N604;
  assign N1428 = ~N1427;
  assign N1429 = N529 & N1428;
  assign N1430 = N1426 | N598;
  assign N1431 = ~N1430;
  assign N1432 = N529 & N1431;
  assign N1433 = ~N598;
  assign N1434 = N340 & N602;
  assign N1435 = N1434 | N598;
  assign N1436 = ~N1435;
  assign N1437 = N529 & N1436;
  assign N1438 = N529 & N1436;
  assign N1439 = N338 & N602;
  assign N1440 = N1439 | N598;
  assign N1441 = ~N1440;
  assign N1442 = N529 & N1441;
  assign N1443 = N338 & N596;
  assign N1444 = N1443 | N598;
  assign N1445 = ~N1444;
  assign N1446 = N529 & N1445;
  assign N1447 = N1443 | N594;
  assign N1448 = ~N1447;
  assign N1449 = N529 & N1448;
  assign N1450 = N336 & N596;
  assign N1451 = N1450 | N594;
  assign N1452 = ~N1451;
  assign N1453 = N529 & N1452;
  assign N1454 = N529 & N1452;
  assign N1455 = N529 & N1452;
  assign N1456 = N529 & N1452;
  assign N1457 = N529 & N1452;
  assign N1458 = N529 & N1452;
  assign N1459 = N529 & N1452;
  assign N1460 = N529 & N1452;
  assign N1461 = N529 & N1452;
  assign N1462 = N529 & N1452;
  assign N1463 = N529 & N1452;
  assign N1464 = N529 & N1452;
  assign N1465 = N529 & N1452;
  assign N1466 = N529 & N1452;
  assign N1467 = N529 & N1452;
  assign N1468 = N529 & N1452;
  assign N1469 = N529 & N1452;
  assign N1470 = N529 & N1452;
  assign N1471 = N529 & N1452;
  assign N1472 = N529 & N1452;
  assign N1473 = N529 & N1452;
  assign N1474 = N529 & N1452;
  assign N1475 = N529 & N1452;
  assign N1476 = N529 & N1452;
  assign N1477 = N529 & N1452;
  assign N1478 = N529 & N1452;
  assign N1479 = N529 & N1452;
  assign N1480 = N529 & N1452;
  assign N1481 = N529 & N1452;
  assign N1482 = N529 & N1452;
  assign N1483 = N529 & N1452;
  assign N1484 = N529 & N1452;
  assign N1485 = N529 & N1452;
  assign N1486 = N529 & N1452;
  assign N1487 = N529 & N1452;
  assign N1488 = N529 & N1452;
  assign N1489 = N529 & N1452;
  assign N1490 = N529 & N1452;
  assign N1491 = N529 & N1452;
  assign N1492 = N529 & N1452;
  assign N1493 = N529 & N1452;

endmodule