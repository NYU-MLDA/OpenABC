module bsg_dff_reset_en_width_p173
(
  clk_i,
  reset_i,
  en_i,
  data_i,
  data_o
);

  input [172:0] data_i;
  output [172:0] data_o;
  input clk_i;
  input reset_i;
  input en_i;
  wire [172:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179;
  reg data_o_172_sv2v_reg,data_o_171_sv2v_reg,data_o_170_sv2v_reg,data_o_169_sv2v_reg,
  data_o_168_sv2v_reg,data_o_167_sv2v_reg,data_o_166_sv2v_reg,data_o_165_sv2v_reg,
  data_o_164_sv2v_reg,data_o_163_sv2v_reg,data_o_162_sv2v_reg,data_o_161_sv2v_reg,
  data_o_160_sv2v_reg,data_o_159_sv2v_reg,data_o_158_sv2v_reg,data_o_157_sv2v_reg,
  data_o_156_sv2v_reg,data_o_155_sv2v_reg,data_o_154_sv2v_reg,data_o_153_sv2v_reg,
  data_o_152_sv2v_reg,data_o_151_sv2v_reg,data_o_150_sv2v_reg,data_o_149_sv2v_reg,
  data_o_148_sv2v_reg,data_o_147_sv2v_reg,data_o_146_sv2v_reg,data_o_145_sv2v_reg,
  data_o_144_sv2v_reg,data_o_143_sv2v_reg,data_o_142_sv2v_reg,data_o_141_sv2v_reg,
  data_o_140_sv2v_reg,data_o_139_sv2v_reg,data_o_138_sv2v_reg,data_o_137_sv2v_reg,
  data_o_136_sv2v_reg,data_o_135_sv2v_reg,data_o_134_sv2v_reg,data_o_133_sv2v_reg,
  data_o_132_sv2v_reg,data_o_131_sv2v_reg,data_o_130_sv2v_reg,data_o_129_sv2v_reg,
  data_o_128_sv2v_reg,data_o_127_sv2v_reg,data_o_126_sv2v_reg,data_o_125_sv2v_reg,
  data_o_124_sv2v_reg,data_o_123_sv2v_reg,data_o_122_sv2v_reg,data_o_121_sv2v_reg,
  data_o_120_sv2v_reg,data_o_119_sv2v_reg,data_o_118_sv2v_reg,data_o_117_sv2v_reg,
  data_o_116_sv2v_reg,data_o_115_sv2v_reg,data_o_114_sv2v_reg,data_o_113_sv2v_reg,
  data_o_112_sv2v_reg,data_o_111_sv2v_reg,data_o_110_sv2v_reg,data_o_109_sv2v_reg,
  data_o_108_sv2v_reg,data_o_107_sv2v_reg,data_o_106_sv2v_reg,data_o_105_sv2v_reg,
  data_o_104_sv2v_reg,data_o_103_sv2v_reg,data_o_102_sv2v_reg,data_o_101_sv2v_reg,
  data_o_100_sv2v_reg,data_o_99_sv2v_reg,data_o_98_sv2v_reg,data_o_97_sv2v_reg,
  data_o_96_sv2v_reg,data_o_95_sv2v_reg,data_o_94_sv2v_reg,data_o_93_sv2v_reg,
  data_o_92_sv2v_reg,data_o_91_sv2v_reg,data_o_90_sv2v_reg,data_o_89_sv2v_reg,
  data_o_88_sv2v_reg,data_o_87_sv2v_reg,data_o_86_sv2v_reg,data_o_85_sv2v_reg,
  data_o_84_sv2v_reg,data_o_83_sv2v_reg,data_o_82_sv2v_reg,data_o_81_sv2v_reg,data_o_80_sv2v_reg,
  data_o_79_sv2v_reg,data_o_78_sv2v_reg,data_o_77_sv2v_reg,data_o_76_sv2v_reg,
  data_o_75_sv2v_reg,data_o_74_sv2v_reg,data_o_73_sv2v_reg,data_o_72_sv2v_reg,
  data_o_71_sv2v_reg,data_o_70_sv2v_reg,data_o_69_sv2v_reg,data_o_68_sv2v_reg,
  data_o_67_sv2v_reg,data_o_66_sv2v_reg,data_o_65_sv2v_reg,data_o_64_sv2v_reg,
  data_o_63_sv2v_reg,data_o_62_sv2v_reg,data_o_61_sv2v_reg,data_o_60_sv2v_reg,data_o_59_sv2v_reg,
  data_o_58_sv2v_reg,data_o_57_sv2v_reg,data_o_56_sv2v_reg,data_o_55_sv2v_reg,
  data_o_54_sv2v_reg,data_o_53_sv2v_reg,data_o_52_sv2v_reg,data_o_51_sv2v_reg,
  data_o_50_sv2v_reg,data_o_49_sv2v_reg,data_o_48_sv2v_reg,data_o_47_sv2v_reg,
  data_o_46_sv2v_reg,data_o_45_sv2v_reg,data_o_44_sv2v_reg,data_o_43_sv2v_reg,
  data_o_42_sv2v_reg,data_o_41_sv2v_reg,data_o_40_sv2v_reg,data_o_39_sv2v_reg,data_o_38_sv2v_reg,
  data_o_37_sv2v_reg,data_o_36_sv2v_reg,data_o_35_sv2v_reg,data_o_34_sv2v_reg,
  data_o_33_sv2v_reg,data_o_32_sv2v_reg,data_o_31_sv2v_reg,data_o_30_sv2v_reg,
  data_o_29_sv2v_reg,data_o_28_sv2v_reg,data_o_27_sv2v_reg,data_o_26_sv2v_reg,
  data_o_25_sv2v_reg,data_o_24_sv2v_reg,data_o_23_sv2v_reg,data_o_22_sv2v_reg,
  data_o_21_sv2v_reg,data_o_20_sv2v_reg,data_o_19_sv2v_reg,data_o_18_sv2v_reg,data_o_17_sv2v_reg,
  data_o_16_sv2v_reg,data_o_15_sv2v_reg,data_o_14_sv2v_reg,data_o_13_sv2v_reg,
  data_o_12_sv2v_reg,data_o_11_sv2v_reg,data_o_10_sv2v_reg,data_o_9_sv2v_reg,
  data_o_8_sv2v_reg,data_o_7_sv2v_reg,data_o_6_sv2v_reg,data_o_5_sv2v_reg,data_o_4_sv2v_reg,
  data_o_3_sv2v_reg,data_o_2_sv2v_reg,data_o_1_sv2v_reg,data_o_0_sv2v_reg;
  assign data_o[172] = data_o_172_sv2v_reg;
  assign data_o[171] = data_o_171_sv2v_reg;
  assign data_o[170] = data_o_170_sv2v_reg;
  assign data_o[169] = data_o_169_sv2v_reg;
  assign data_o[168] = data_o_168_sv2v_reg;
  assign data_o[167] = data_o_167_sv2v_reg;
  assign data_o[166] = data_o_166_sv2v_reg;
  assign data_o[165] = data_o_165_sv2v_reg;
  assign data_o[164] = data_o_164_sv2v_reg;
  assign data_o[163] = data_o_163_sv2v_reg;
  assign data_o[162] = data_o_162_sv2v_reg;
  assign data_o[161] = data_o_161_sv2v_reg;
  assign data_o[160] = data_o_160_sv2v_reg;
  assign data_o[159] = data_o_159_sv2v_reg;
  assign data_o[158] = data_o_158_sv2v_reg;
  assign data_o[157] = data_o_157_sv2v_reg;
  assign data_o[156] = data_o_156_sv2v_reg;
  assign data_o[155] = data_o_155_sv2v_reg;
  assign data_o[154] = data_o_154_sv2v_reg;
  assign data_o[153] = data_o_153_sv2v_reg;
  assign data_o[152] = data_o_152_sv2v_reg;
  assign data_o[151] = data_o_151_sv2v_reg;
  assign data_o[150] = data_o_150_sv2v_reg;
  assign data_o[149] = data_o_149_sv2v_reg;
  assign data_o[148] = data_o_148_sv2v_reg;
  assign data_o[147] = data_o_147_sv2v_reg;
  assign data_o[146] = data_o_146_sv2v_reg;
  assign data_o[145] = data_o_145_sv2v_reg;
  assign data_o[144] = data_o_144_sv2v_reg;
  assign data_o[143] = data_o_143_sv2v_reg;
  assign data_o[142] = data_o_142_sv2v_reg;
  assign data_o[141] = data_o_141_sv2v_reg;
  assign data_o[140] = data_o_140_sv2v_reg;
  assign data_o[139] = data_o_139_sv2v_reg;
  assign data_o[138] = data_o_138_sv2v_reg;
  assign data_o[137] = data_o_137_sv2v_reg;
  assign data_o[136] = data_o_136_sv2v_reg;
  assign data_o[135] = data_o_135_sv2v_reg;
  assign data_o[134] = data_o_134_sv2v_reg;
  assign data_o[133] = data_o_133_sv2v_reg;
  assign data_o[132] = data_o_132_sv2v_reg;
  assign data_o[131] = data_o_131_sv2v_reg;
  assign data_o[130] = data_o_130_sv2v_reg;
  assign data_o[129] = data_o_129_sv2v_reg;
  assign data_o[128] = data_o_128_sv2v_reg;
  assign data_o[127] = data_o_127_sv2v_reg;
  assign data_o[126] = data_o_126_sv2v_reg;
  assign data_o[125] = data_o_125_sv2v_reg;
  assign data_o[124] = data_o_124_sv2v_reg;
  assign data_o[123] = data_o_123_sv2v_reg;
  assign data_o[122] = data_o_122_sv2v_reg;
  assign data_o[121] = data_o_121_sv2v_reg;
  assign data_o[120] = data_o_120_sv2v_reg;
  assign data_o[119] = data_o_119_sv2v_reg;
  assign data_o[118] = data_o_118_sv2v_reg;
  assign data_o[117] = data_o_117_sv2v_reg;
  assign data_o[116] = data_o_116_sv2v_reg;
  assign data_o[115] = data_o_115_sv2v_reg;
  assign data_o[114] = data_o_114_sv2v_reg;
  assign data_o[113] = data_o_113_sv2v_reg;
  assign data_o[112] = data_o_112_sv2v_reg;
  assign data_o[111] = data_o_111_sv2v_reg;
  assign data_o[110] = data_o_110_sv2v_reg;
  assign data_o[109] = data_o_109_sv2v_reg;
  assign data_o[108] = data_o_108_sv2v_reg;
  assign data_o[107] = data_o_107_sv2v_reg;
  assign data_o[106] = data_o_106_sv2v_reg;
  assign data_o[105] = data_o_105_sv2v_reg;
  assign data_o[104] = data_o_104_sv2v_reg;
  assign data_o[103] = data_o_103_sv2v_reg;
  assign data_o[102] = data_o_102_sv2v_reg;
  assign data_o[101] = data_o_101_sv2v_reg;
  assign data_o[100] = data_o_100_sv2v_reg;
  assign data_o[99] = data_o_99_sv2v_reg;
  assign data_o[98] = data_o_98_sv2v_reg;
  assign data_o[97] = data_o_97_sv2v_reg;
  assign data_o[96] = data_o_96_sv2v_reg;
  assign data_o[95] = data_o_95_sv2v_reg;
  assign data_o[94] = data_o_94_sv2v_reg;
  assign data_o[93] = data_o_93_sv2v_reg;
  assign data_o[92] = data_o_92_sv2v_reg;
  assign data_o[91] = data_o_91_sv2v_reg;
  assign data_o[90] = data_o_90_sv2v_reg;
  assign data_o[89] = data_o_89_sv2v_reg;
  assign data_o[88] = data_o_88_sv2v_reg;
  assign data_o[87] = data_o_87_sv2v_reg;
  assign data_o[86] = data_o_86_sv2v_reg;
  assign data_o[85] = data_o_85_sv2v_reg;
  assign data_o[84] = data_o_84_sv2v_reg;
  assign data_o[83] = data_o_83_sv2v_reg;
  assign data_o[82] = data_o_82_sv2v_reg;
  assign data_o[81] = data_o_81_sv2v_reg;
  assign data_o[80] = data_o_80_sv2v_reg;
  assign data_o[79] = data_o_79_sv2v_reg;
  assign data_o[78] = data_o_78_sv2v_reg;
  assign data_o[77] = data_o_77_sv2v_reg;
  assign data_o[76] = data_o_76_sv2v_reg;
  assign data_o[75] = data_o_75_sv2v_reg;
  assign data_o[74] = data_o_74_sv2v_reg;
  assign data_o[73] = data_o_73_sv2v_reg;
  assign data_o[72] = data_o_72_sv2v_reg;
  assign data_o[71] = data_o_71_sv2v_reg;
  assign data_o[70] = data_o_70_sv2v_reg;
  assign data_o[69] = data_o_69_sv2v_reg;
  assign data_o[68] = data_o_68_sv2v_reg;
  assign data_o[67] = data_o_67_sv2v_reg;
  assign data_o[66] = data_o_66_sv2v_reg;
  assign data_o[65] = data_o_65_sv2v_reg;
  assign data_o[64] = data_o_64_sv2v_reg;
  assign data_o[63] = data_o_63_sv2v_reg;
  assign data_o[62] = data_o_62_sv2v_reg;
  assign data_o[61] = data_o_61_sv2v_reg;
  assign data_o[60] = data_o_60_sv2v_reg;
  assign data_o[59] = data_o_59_sv2v_reg;
  assign data_o[58] = data_o_58_sv2v_reg;
  assign data_o[57] = data_o_57_sv2v_reg;
  assign data_o[56] = data_o_56_sv2v_reg;
  assign data_o[55] = data_o_55_sv2v_reg;
  assign data_o[54] = data_o_54_sv2v_reg;
  assign data_o[53] = data_o_53_sv2v_reg;
  assign data_o[52] = data_o_52_sv2v_reg;
  assign data_o[51] = data_o_51_sv2v_reg;
  assign data_o[50] = data_o_50_sv2v_reg;
  assign data_o[49] = data_o_49_sv2v_reg;
  assign data_o[48] = data_o_48_sv2v_reg;
  assign data_o[47] = data_o_47_sv2v_reg;
  assign data_o[46] = data_o_46_sv2v_reg;
  assign data_o[45] = data_o_45_sv2v_reg;
  assign data_o[44] = data_o_44_sv2v_reg;
  assign data_o[43] = data_o_43_sv2v_reg;
  assign data_o[42] = data_o_42_sv2v_reg;
  assign data_o[41] = data_o_41_sv2v_reg;
  assign data_o[40] = data_o_40_sv2v_reg;
  assign data_o[39] = data_o_39_sv2v_reg;
  assign data_o[38] = data_o_38_sv2v_reg;
  assign data_o[37] = data_o_37_sv2v_reg;
  assign data_o[36] = data_o_36_sv2v_reg;
  assign data_o[35] = data_o_35_sv2v_reg;
  assign data_o[34] = data_o_34_sv2v_reg;
  assign data_o[33] = data_o_33_sv2v_reg;
  assign data_o[32] = data_o_32_sv2v_reg;
  assign data_o[31] = data_o_31_sv2v_reg;
  assign data_o[30] = data_o_30_sv2v_reg;
  assign data_o[29] = data_o_29_sv2v_reg;
  assign data_o[28] = data_o_28_sv2v_reg;
  assign data_o[27] = data_o_27_sv2v_reg;
  assign data_o[26] = data_o_26_sv2v_reg;
  assign data_o[25] = data_o_25_sv2v_reg;
  assign data_o[24] = data_o_24_sv2v_reg;
  assign data_o[23] = data_o_23_sv2v_reg;
  assign data_o[22] = data_o_22_sv2v_reg;
  assign data_o[21] = data_o_21_sv2v_reg;
  assign data_o[20] = data_o_20_sv2v_reg;
  assign data_o[19] = data_o_19_sv2v_reg;
  assign data_o[18] = data_o_18_sv2v_reg;
  assign data_o[17] = data_o_17_sv2v_reg;
  assign data_o[16] = data_o_16_sv2v_reg;
  assign data_o[15] = data_o_15_sv2v_reg;
  assign data_o[14] = data_o_14_sv2v_reg;
  assign data_o[13] = data_o_13_sv2v_reg;
  assign data_o[12] = data_o_12_sv2v_reg;
  assign data_o[11] = data_o_11_sv2v_reg;
  assign data_o[10] = data_o_10_sv2v_reg;
  assign data_o[9] = data_o_9_sv2v_reg;
  assign data_o[8] = data_o_8_sv2v_reg;
  assign data_o[7] = data_o_7_sv2v_reg;
  assign data_o[6] = data_o_6_sv2v_reg;
  assign data_o[5] = data_o_5_sv2v_reg;
  assign data_o[4] = data_o_4_sv2v_reg;
  assign data_o[3] = data_o_3_sv2v_reg;
  assign data_o[2] = data_o_2_sv2v_reg;
  assign data_o[1] = data_o_1_sv2v_reg;
  assign data_o[0] = data_o_0_sv2v_reg;

  always @(posedge clk_i) begin
    if(N3) begin
      data_o_172_sv2v_reg <= N177;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_171_sv2v_reg <= N176;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_170_sv2v_reg <= N175;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_169_sv2v_reg <= N174;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_168_sv2v_reg <= N173;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_167_sv2v_reg <= N172;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_166_sv2v_reg <= N171;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_165_sv2v_reg <= N170;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_164_sv2v_reg <= N169;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_163_sv2v_reg <= N168;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_162_sv2v_reg <= N167;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_161_sv2v_reg <= N166;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_160_sv2v_reg <= N165;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_159_sv2v_reg <= N164;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_158_sv2v_reg <= N163;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_157_sv2v_reg <= N162;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_156_sv2v_reg <= N161;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_155_sv2v_reg <= N160;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_154_sv2v_reg <= N159;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_153_sv2v_reg <= N158;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_152_sv2v_reg <= N157;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_151_sv2v_reg <= N156;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_150_sv2v_reg <= N155;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_149_sv2v_reg <= N154;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_148_sv2v_reg <= N153;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_147_sv2v_reg <= N152;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_146_sv2v_reg <= N151;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_145_sv2v_reg <= N150;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_144_sv2v_reg <= N149;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_143_sv2v_reg <= N148;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_142_sv2v_reg <= N147;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_141_sv2v_reg <= N146;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_140_sv2v_reg <= N145;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_139_sv2v_reg <= N144;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_138_sv2v_reg <= N143;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_137_sv2v_reg <= N142;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_136_sv2v_reg <= N141;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_135_sv2v_reg <= N140;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_134_sv2v_reg <= N139;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_133_sv2v_reg <= N138;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_132_sv2v_reg <= N137;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_131_sv2v_reg <= N136;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_130_sv2v_reg <= N135;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_129_sv2v_reg <= N134;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_128_sv2v_reg <= N133;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_127_sv2v_reg <= N132;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_126_sv2v_reg <= N131;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_125_sv2v_reg <= N130;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_124_sv2v_reg <= N129;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_123_sv2v_reg <= N128;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_122_sv2v_reg <= N127;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_121_sv2v_reg <= N126;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_120_sv2v_reg <= N125;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_119_sv2v_reg <= N124;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_118_sv2v_reg <= N123;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_117_sv2v_reg <= N122;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_116_sv2v_reg <= N121;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_115_sv2v_reg <= N120;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_114_sv2v_reg <= N119;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_113_sv2v_reg <= N118;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_112_sv2v_reg <= N117;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_111_sv2v_reg <= N116;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_110_sv2v_reg <= N115;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_109_sv2v_reg <= N114;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_108_sv2v_reg <= N113;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_107_sv2v_reg <= N112;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_106_sv2v_reg <= N111;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_105_sv2v_reg <= N110;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_104_sv2v_reg <= N109;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_103_sv2v_reg <= N108;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_102_sv2v_reg <= N107;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_101_sv2v_reg <= N106;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_100_sv2v_reg <= N105;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_99_sv2v_reg <= N104;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_98_sv2v_reg <= N103;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_97_sv2v_reg <= N102;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_96_sv2v_reg <= N101;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_95_sv2v_reg <= N100;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_94_sv2v_reg <= N99;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_93_sv2v_reg <= N98;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_92_sv2v_reg <= N97;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_91_sv2v_reg <= N96;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_90_sv2v_reg <= N95;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_89_sv2v_reg <= N94;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_88_sv2v_reg <= N93;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_87_sv2v_reg <= N92;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_86_sv2v_reg <= N91;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_85_sv2v_reg <= N90;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_84_sv2v_reg <= N89;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_83_sv2v_reg <= N88;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_82_sv2v_reg <= N87;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_81_sv2v_reg <= N86;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_80_sv2v_reg <= N85;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_79_sv2v_reg <= N84;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_78_sv2v_reg <= N83;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_77_sv2v_reg <= N82;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_76_sv2v_reg <= N81;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_75_sv2v_reg <= N80;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_74_sv2v_reg <= N79;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_73_sv2v_reg <= N78;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_72_sv2v_reg <= N77;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_71_sv2v_reg <= N76;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_70_sv2v_reg <= N75;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_69_sv2v_reg <= N74;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_68_sv2v_reg <= N73;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_67_sv2v_reg <= N72;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_66_sv2v_reg <= N71;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_65_sv2v_reg <= N70;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_64_sv2v_reg <= N69;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_63_sv2v_reg <= N68;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_62_sv2v_reg <= N67;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_61_sv2v_reg <= N66;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_60_sv2v_reg <= N65;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_59_sv2v_reg <= N64;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_58_sv2v_reg <= N63;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_57_sv2v_reg <= N62;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_56_sv2v_reg <= N61;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_55_sv2v_reg <= N60;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_54_sv2v_reg <= N59;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_53_sv2v_reg <= N58;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_52_sv2v_reg <= N57;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_51_sv2v_reg <= N56;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_50_sv2v_reg <= N55;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_49_sv2v_reg <= N54;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_48_sv2v_reg <= N53;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_47_sv2v_reg <= N52;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_46_sv2v_reg <= N51;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_45_sv2v_reg <= N50;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_44_sv2v_reg <= N49;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_43_sv2v_reg <= N48;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_42_sv2v_reg <= N47;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_41_sv2v_reg <= N46;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_40_sv2v_reg <= N45;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_39_sv2v_reg <= N44;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_38_sv2v_reg <= N43;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_37_sv2v_reg <= N42;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_36_sv2v_reg <= N41;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_35_sv2v_reg <= N40;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_34_sv2v_reg <= N39;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_33_sv2v_reg <= N38;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_32_sv2v_reg <= N37;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_31_sv2v_reg <= N36;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_30_sv2v_reg <= N35;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_29_sv2v_reg <= N34;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_28_sv2v_reg <= N33;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_27_sv2v_reg <= N32;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_26_sv2v_reg <= N31;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_25_sv2v_reg <= N30;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_24_sv2v_reg <= N29;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_23_sv2v_reg <= N28;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_22_sv2v_reg <= N27;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_21_sv2v_reg <= N26;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_20_sv2v_reg <= N25;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_19_sv2v_reg <= N24;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_18_sv2v_reg <= N23;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_17_sv2v_reg <= N22;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_16_sv2v_reg <= N21;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_15_sv2v_reg <= N20;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_14_sv2v_reg <= N19;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_13_sv2v_reg <= N18;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_12_sv2v_reg <= N17;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_11_sv2v_reg <= N16;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_10_sv2v_reg <= N15;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_9_sv2v_reg <= N14;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_8_sv2v_reg <= N13;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_7_sv2v_reg <= N12;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_6_sv2v_reg <= N11;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_5_sv2v_reg <= N10;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_4_sv2v_reg <= N9;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_3_sv2v_reg <= N8;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_2_sv2v_reg <= N7;
    end 
  end


  always @(posedge clk_i) begin
    if(N5) begin
      data_o_1_sv2v_reg <= N6;
    end 
  end


  always @(posedge clk_i) begin
    if(N3) begin
      data_o_0_sv2v_reg <= N4;
    end 
  end

  assign { N5, N3 } = (N0)? { 1'b1, 1'b1 } : 
                      (N179)? { 1'b1, 1'b1 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N0 = reset_i;
  assign { N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N4 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        (N179)? data_i : 1'b0;
  assign N1 = en_i | reset_i;
  assign N2 = ~N1;
  assign N178 = ~reset_i;
  assign N179 = en_i & N178;

endmodule