module mmu(clk, rst, \l_in.valid , \l_in.tlbie , \l_in.slbia , \l_in.mtspr , \l_in.iside , \l_in.load , \l_in.priv , \l_in.sprn , \l_in.addr , \l_in.rs , \d_in.stall , \d_in.done , \d_in.err , \d_in.data , \l_out.done , \l_out.err , \l_out.invalid , \l_out.badtree , \l_out.segerr , \l_out.perm_error , \l_out.rc_error , \l_out.sprval , \d_out.valid , \d_out.tlbie , \d_out.doall , \d_out.tlbld , \d_out.addr , \d_out.pte , \i_out.tlbld , \i_out.tlbie , \i_out.doall , \i_out.addr , \i_out.pte );
  wire [63:0] _000_;
  wire _001_;
  wire [67:0] _002_;
  wire [99:0] _003_;
  wire [65:0] _004_;
  wire _005_;
  wire [63:0] _006_;
  wire _007_;
  wire [63:0] _008_;
  wire _009_;
  wire [135:0] _010_;
  reg [501:0] _011_;
  wire _012_;
  wire _013_;
  wire [30:0] _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire [18:0] _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire [15:0] _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire [63:0] _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire [3:0] _149_;
  wire _150_;
  wire [3:0] _151_;
  wire [5:0] _152_;
  wire _153_;
  wire [3:0] _154_;
  wire [5:0] _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire [3:0] _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire [5:0] _163_;
  wire _164_;
  wire [3:0] _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire [63:0] _170_;
  wire [31:0] _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire [100:0] _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire [67:0] _181_;
  wire [5:0] _182_;
  wire _183_;
  wire _184_;
  wire [3:0] _185_;
  wire _186_;
  wire _187_;
  wire [3:0] _188_;
  wire [64:0] _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire [64:0] _193_;
  wire [64:0] _194_;
  wire _195_;
  wire [3:0] _196_;
  wire _197_;
  wire [3:0] _198_;
  wire [196:0] _199_;
  wire _200_;
  wire [3:0] _201_;
  wire _202_;
  wire _203_;
  wire [5:0] _204_;
  wire [5:0] _205_;
  wire [30:0] _206_;
  wire [30:0] _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire [5:0] _214_;
  wire _215_;
  wire _216_;
  wire [3:0] _217_;
  wire _218_;
  wire [3:0] _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire [3:0] _239_;
  wire [1:0] _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire [5:0] _246_;
  wire [3:0] _247_;
  wire [66:0] _248_;
  wire _249_;
  wire [3:0] _250_;
  wire [66:0] _251_;
  wire _252_;
  wire [1:0] _253_;
  wire [3:0] _254_;
  wire [66:0] _255_;
  wire _256_;
  wire _257_;
  wire [1:0] _258_;
  wire [3:0] _259_;
  wire [1:0] _260_;
  wire [3:0] _261_;
  wire _262_;
  wire _263_;
  wire [131:0] _264_;
  wire _265_;
  wire _266_;
  wire [3:0] _267_;
  wire _268_;
  wire _269_;
  wire _270_;
  wire _271_;
  wire [67:0] _272_;
  wire [96:0] _273_;
  wire [3:0] _274_;
  wire [63:0] _275_;
  wire _276_;
  wire [63:0] _277_;
  wire _278_;
  wire [63:0] _279_;
  wire _280_;
  wire [5:0] _281_;
  wire [4:0] _282_;
  wire [55:0] _283_;
  wire [63:0] _284_;
  wire _285_;
  wire _286_;
  wire _287_;
  wire [1:0] _288_;
  wire _289_;
  wire _290_;
  wire _291_;
  wire _292_;
  wire _293_;
  wire _294_;
  wire _295_;
  wire _296_;
  wire _297_;
  wire _298_;
  wire _299_;
  wire _300_;
  wire _301_;
  wire _302_;
  wire _303_;
  wire [1:0] _304_;
  wire [31:0] _305_;
  wire [23:0] _306_;
  wire [23:0] _307_;
  wire [23:0] _308_;
  wire [23:0] _309_;
  wire [15:0] _310_;
  wire [15:0] _311_;
  wire [15:0] _312_;
  wire [15:0] _313_;
  wire [43:0] _314_;
  wire [43:0] _315_;
  wire [43:0] _316_;
  wire [43:0] _317_;
  wire [63:0] _318_;
  wire [63:0] _319_;
  wire [63:0] _320_;
  wire [63:0] _321_;
  wire [63:0] _322_;
  wire [63:0] _323_;
  wire [15:0] addrsh;
  input clk;
  wire clk;
  input [63:0] \d_in.data ;
  wire [63:0] \d_in.data ;
  input \d_in.done ;
  wire \d_in.done ;
  input \d_in.err ;
  wire \d_in.err ;
  input \d_in.stall ;
  wire \d_in.stall ;
  output [63:0] \d_out.addr ;
  wire [63:0] \d_out.addr ;
  output \d_out.doall ;
  wire \d_out.doall ;
  output [63:0] \d_out.pte ;
  wire [63:0] \d_out.pte ;
  output \d_out.tlbie ;
  wire \d_out.tlbie ;
  output \d_out.tlbld ;
  wire \d_out.tlbld ;
  output \d_out.valid ;
  wire \d_out.valid ;
  wire [43:0] finalmask;
  output [63:0] \i_out.addr ;
  wire [63:0] \i_out.addr ;
  output \i_out.doall ;
  wire \i_out.doall ;
  output [63:0] \i_out.pte ;
  wire [63:0] \i_out.pte ;
  output \i_out.tlbie ;
  wire \i_out.tlbie ;
  output \i_out.tlbld ;
  wire \i_out.tlbld ;
  input [63:0] \l_in.addr ;
  wire [63:0] \l_in.addr ;
  input \l_in.iside ;
  wire \l_in.iside ;
  input \l_in.load ;
  wire \l_in.load ;
  input \l_in.mtspr ;
  wire \l_in.mtspr ;
  input \l_in.priv ;
  wire \l_in.priv ;
  input [63:0] \l_in.rs ;
  wire [63:0] \l_in.rs ;
  input \l_in.slbia ;
  wire \l_in.slbia ;
  input [9:0] \l_in.sprn ;
  wire [9:0] \l_in.sprn ;
  input \l_in.tlbie ;
  wire \l_in.tlbie ;
  input \l_in.valid ;
  wire \l_in.valid ;
  output \l_out.badtree ;
  wire \l_out.badtree ;
  output \l_out.done ;
  wire \l_out.done ;
  output \l_out.err ;
  wire \l_out.err ;
  output \l_out.invalid ;
  wire \l_out.invalid ;
  output \l_out.perm_error ;
  wire \l_out.perm_error ;
  output \l_out.rc_error ;
  wire \l_out.rc_error ;
  output \l_out.segerr ;
  wire \l_out.segerr ;
  output [63:0] \l_out.sprval ;
  wire [63:0] \l_out.sprval ;
  wire [15:0] mask;
  wire [501:0] r;
  wire [501:0] rin;
  input rst;
  wire rst;
  assign _000_ = \l_in.sprn [8] ? r[132:69] : { 32'h00000000, r[164:133] };
  assign _001_ = rst ? 1'h0 : rin[0];
  assign _002_ = rst ? r[68:1] : rin[68:1];
  assign _003_ = rst ? 100'h0000000000000000000000000 : rin[168:69];
  assign _004_ = rst ? r[234:169] : rin[234:169];
  assign _005_ = rst ? 1'h0 : rin[235];
  assign _006_ = rst ? r[299:236] : rin[299:236];
  assign _007_ = rst ? 1'h0 : rin[300];
  assign _008_ = rst ? r[364:301] : rin[364:301];
  assign _009_ = rst ? 1'h0 : rin[365];
  assign _010_ = rst ? r[501:366] : rin[501:366];
  always @(posedge clk)
    _011_ <= { _010_, _009_, _008_, _007_, _006_, _005_, _004_, _003_, _002_, _001_ };
  assign _012_ = r[371:370] == 2'h0;
  assign _013_ = r[371:370] == 2'h1;
  function [30:0] \22555 ;
    input [30:0] a;
    input [61:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \22555  = b[30:0];
      2'b1?:
        \22555  = b[61:31];
      default:
        \22555  = a;
    endcase
  endfunction
  assign _014_ = \22555 ({ 13'h0000, r[65:48] }, { r[62:32], r[46:16] }, { _013_, _012_ });
  assign _015_ = r[369:368] == 2'h0;
  assign _016_ = r[369:368] == 2'h1;
  assign _017_ = r[369:368] == 2'h2;
  function [18:0] \22568 ;
    input [18:0] a;
    input [56:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \22568  = b[18:0];
      3'b?1?:
        \22568  = b[37:19];
      3'b1??:
        \22568  = b[56:38];
      default:
        \22568  = a;
    endcase
  endfunction
  assign _018_ = \22568 (_014_[30:12], { _014_[26:8], _014_[22:4], _014_[18:0] }, { _017_, _016_, _015_ });
  assign _019_ = r[367:366] == 2'h0;
  assign _020_ = r[367:366] == 2'h1;
  assign _021_ = r[367:366] == 2'h2;
  function [15:0] \22581 ;
    input [15:0] a;
    input [47:0] b;
    input [2:0] s;
    (* parallel_case *)
    casez (s)
      3'b??1:
        \22581  = b[15:0];
      3'b?1?:
        \22581  = b[31:16];
      3'b1??:
        \22581  = b[47:32];
      default:
        \22581  = a;
    endcase
  endfunction
  assign _022_ = \22581 (_018_[18:3], { _018_[17:2], _018_[16:1], _018_[15:0] }, { _021_, _020_, _019_ });
  assign _023_ = $signed(32'd5) < $signed({ 27'h0000000, r[376:372] });
  assign _024_ = _023_ ? 1'h1 : 1'h0;
  assign _025_ = $signed(32'd6) < $signed({ 27'h0000000, r[376:372] });
  assign _026_ = _025_ ? 1'h1 : 1'h0;
  assign _027_ = $signed(32'd7) < $signed({ 27'h0000000, r[376:372] });
  assign _028_ = _027_ ? 1'h1 : 1'h0;
  assign _029_ = $signed(32'd8) < $signed({ 27'h0000000, r[376:372] });
  assign _030_ = _029_ ? 1'h1 : 1'h0;
  assign _031_ = $signed(32'd9) < $signed({ 27'h0000000, r[376:372] });
  assign _032_ = _031_ ? 1'h1 : 1'h0;
  assign _033_ = $signed(32'd10) < $signed({ 27'h0000000, r[376:372] });
  assign _034_ = _033_ ? 1'h1 : 1'h0;
  assign _035_ = $signed(32'd11) < $signed({ 27'h0000000, r[376:372] });
  assign _036_ = _035_ ? 1'h1 : 1'h0;
  assign _037_ = $signed(32'd12) < $signed({ 27'h0000000, r[376:372] });
  assign _038_ = _037_ ? 1'h1 : 1'h0;
  assign _039_ = $signed(32'd13) < $signed({ 27'h0000000, r[376:372] });
  assign _040_ = _039_ ? 1'h1 : 1'h0;
  assign _041_ = $signed(32'd14) < $signed({ 27'h0000000, r[376:372] });
  assign _042_ = _041_ ? 1'h1 : 1'h0;
  assign _043_ = $signed(32'd15) < $signed({ 27'h0000000, r[376:372] });
  assign _044_ = _043_ ? 1'h1 : 1'h0;
  assign _045_ = $signed(32'd0) < $signed({ 26'h0000000, r[371:366] });
  assign _046_ = _045_ ? 1'h1 : 1'h0;
  assign _047_ = $signed(32'd1) < $signed({ 26'h0000000, r[371:366] });
  assign _048_ = _047_ ? 1'h1 : 1'h0;
  assign _049_ = $signed(32'd2) < $signed({ 26'h0000000, r[371:366] });
  assign _050_ = _049_ ? 1'h1 : 1'h0;
  assign _051_ = $signed(32'd3) < $signed({ 26'h0000000, r[371:366] });
  assign _052_ = _051_ ? 1'h1 : 1'h0;
  assign _053_ = $signed(32'd4) < $signed({ 26'h0000000, r[371:366] });
  assign _054_ = _053_ ? 1'h1 : 1'h0;
  assign _055_ = $signed(32'd5) < $signed({ 26'h0000000, r[371:366] });
  assign _056_ = _055_ ? 1'h1 : 1'h0;
  assign _057_ = $signed(32'd6) < $signed({ 26'h0000000, r[371:366] });
  assign _058_ = _057_ ? 1'h1 : 1'h0;
  assign _059_ = $signed(32'd7) < $signed({ 26'h0000000, r[371:366] });
  assign _060_ = _059_ ? 1'h1 : 1'h0;
  assign _061_ = $signed(32'd8) < $signed({ 26'h0000000, r[371:366] });
  assign _062_ = _061_ ? 1'h1 : 1'h0;
  assign _063_ = $signed(32'd9) < $signed({ 26'h0000000, r[371:366] });
  assign _064_ = _063_ ? 1'h1 : 1'h0;
  assign _065_ = $signed(32'd10) < $signed({ 26'h0000000, r[371:366] });
  assign _066_ = _065_ ? 1'h1 : 1'h0;
  assign _067_ = $signed(32'd11) < $signed({ 26'h0000000, r[371:366] });
  assign _068_ = _067_ ? 1'h1 : 1'h0;
  assign _069_ = $signed(32'd12) < $signed({ 26'h0000000, r[371:366] });
  assign _070_ = _069_ ? 1'h1 : 1'h0;
  assign _071_ = $signed(32'd13) < $signed({ 26'h0000000, r[371:366] });
  assign _072_ = _071_ ? 1'h1 : 1'h0;
  assign _073_ = $signed(32'd14) < $signed({ 26'h0000000, r[371:366] });
  assign _074_ = _073_ ? 1'h1 : 1'h0;
  assign _075_ = $signed(32'd15) < $signed({ 26'h0000000, r[371:366] });
  assign _076_ = _075_ ? 1'h1 : 1'h0;
  assign _077_ = $signed(32'd16) < $signed({ 26'h0000000, r[371:366] });
  assign _078_ = _077_ ? 1'h1 : 1'h0;
  assign _079_ = $signed(32'd17) < $signed({ 26'h0000000, r[371:366] });
  assign _080_ = _079_ ? 1'h1 : 1'h0;
  assign _081_ = $signed(32'd18) < $signed({ 26'h0000000, r[371:366] });
  assign _082_ = _081_ ? 1'h1 : 1'h0;
  assign _083_ = $signed(32'd19) < $signed({ 26'h0000000, r[371:366] });
  assign _084_ = _083_ ? 1'h1 : 1'h0;
  assign _085_ = $signed(32'd20) < $signed({ 26'h0000000, r[371:366] });
  assign _086_ = _085_ ? 1'h1 : 1'h0;
  assign _087_ = $signed(32'd21) < $signed({ 26'h0000000, r[371:366] });
  assign _088_ = _087_ ? 1'h1 : 1'h0;
  assign _089_ = $signed(32'd22) < $signed({ 26'h0000000, r[371:366] });
  assign _090_ = _089_ ? 1'h1 : 1'h0;
  assign _091_ = $signed(32'd23) < $signed({ 26'h0000000, r[371:366] });
  assign _092_ = _091_ ? 1'h1 : 1'h0;
  assign _093_ = $signed(32'd24) < $signed({ 26'h0000000, r[371:366] });
  assign _094_ = _093_ ? 1'h1 : 1'h0;
  assign _095_ = $signed(32'd25) < $signed({ 26'h0000000, r[371:366] });
  assign _096_ = _095_ ? 1'h1 : 1'h0;
  assign _097_ = $signed(32'd26) < $signed({ 26'h0000000, r[371:366] });
  assign _098_ = _097_ ? 1'h1 : 1'h0;
  assign _099_ = $signed(32'd27) < $signed({ 26'h0000000, r[371:366] });
  assign _100_ = _099_ ? 1'h1 : 1'h0;
  assign _101_ = $signed(32'd28) < $signed({ 26'h0000000, r[371:366] });
  assign _102_ = _101_ ? 1'h1 : 1'h0;
  assign _103_ = $signed(32'd29) < $signed({ 26'h0000000, r[371:366] });
  assign _104_ = _103_ ? 1'h1 : 1'h0;
  assign _105_ = $signed(32'd30) < $signed({ 26'h0000000, r[371:366] });
  assign _106_ = _105_ ? 1'h1 : 1'h0;
  assign _107_ = $signed(32'd31) < $signed({ 26'h0000000, r[371:366] });
  assign _108_ = _107_ ? 1'h1 : 1'h0;
  assign _109_ = $signed(32'd32) < $signed({ 26'h0000000, r[371:366] });
  assign _110_ = _109_ ? 1'h1 : 1'h0;
  assign _111_ = $signed(32'd33) < $signed({ 26'h0000000, r[371:366] });
  assign _112_ = _111_ ? 1'h1 : 1'h0;
  assign _113_ = $signed(32'd34) < $signed({ 26'h0000000, r[371:366] });
  assign _114_ = _113_ ? 1'h1 : 1'h0;
  assign _115_ = $signed(32'd35) < $signed({ 26'h0000000, r[371:366] });
  assign _116_ = _115_ ? 1'h1 : 1'h0;
  assign _117_ = $signed(32'd36) < $signed({ 26'h0000000, r[371:366] });
  assign _118_ = _117_ ? 1'h1 : 1'h0;
  assign _119_ = $signed(32'd37) < $signed({ 26'h0000000, r[371:366] });
  assign _120_ = _119_ ? 1'h1 : 1'h0;
  assign _121_ = $signed(32'd38) < $signed({ 26'h0000000, r[371:366] });
  assign _122_ = _121_ ? 1'h1 : 1'h0;
  assign _123_ = $signed(32'd39) < $signed({ 26'h0000000, r[371:366] });
  assign _124_ = _123_ ? 1'h1 : 1'h0;
  assign _125_ = $signed(32'd40) < $signed({ 26'h0000000, r[371:366] });
  assign _126_ = _125_ ? 1'h1 : 1'h0;
  assign _127_ = $signed(32'd41) < $signed({ 26'h0000000, r[371:366] });
  assign _128_ = _127_ ? 1'h1 : 1'h0;
  assign _129_ = $signed(32'd42) < $signed({ 26'h0000000, r[371:366] });
  assign _130_ = _129_ ? 1'h1 : 1'h0;
  assign _131_ = $signed(32'd43) < $signed({ 26'h0000000, r[371:366] });
  assign _132_ = _131_ ? 1'h1 : 1'h0;
  assign _133_ = ~ \l_in.addr [63];
  assign _134_ = _133_ ? r[300] : r[365];
  assign _135_ = _133_ ? r[299:236] : r[364:301];
  assign _136_ = \l_in.load  | \l_in.iside ;
  assign _137_ = ~ _136_;
  assign _138_ = \l_in.slbia  | \l_in.addr [11];
  assign _139_ = _138_ | \l_in.addr [10];
  assign _140_ = _139_ | \l_in.addr [7];
  assign _141_ = _140_ | \l_in.addr [6];
  assign _142_ = _141_ | \l_in.addr [5];
  assign _143_ = _166_ ? 1'h0 : r[235];
  assign _144_ = _167_ ? 1'h0 : r[300];
  assign _145_ = _162_ ? 1'h0 : r[365];
  assign _146_ = ~ r[235];
  assign _147_ = ~ _134_;
  assign _148_ = { 1'h0, _135_[4:0] } == 6'h00;
  assign _149_ = _148_ ? 4'hc : 4'h8;
  assign _150_ = _148_ ? 1'h1 : 1'h0;
  assign _151_ = _147_ ? 4'h6 : _149_;
  assign _152_ = _147_ ? { 1'h0, r[175:171] } : { 1'h0, _135_[62:61], _135_[7:5] };
  assign _153_ = _147_ ? 1'h0 : _150_;
  assign _154_ = _146_ ? 4'h3 : _151_;
  assign _155_ = _146_ ? { 1'h0, _135_[62:61], _135_[7:5] } : _152_;
  assign _156_ = _146_ ? 1'h0 : _153_;
  assign _157_ = \l_in.tlbie  ? 1'h0 : 1'h1;
  assign _158_ = \l_in.tlbie  ? _142_ : 1'h0;
  assign _159_ = \l_in.tlbie  ? 4'h1 : _154_;
  assign _160_ = \l_in.tlbie  & \l_in.sprn [3];
  assign _161_ = \l_in.tlbie  & \l_in.sprn [3];
  assign _162_ = \l_in.tlbie  & \l_in.sprn [3];
  assign _163_ = \l_in.tlbie  ? { 1'h0, _135_[62:61], _135_[7:5] } : _155_;
  assign _164_ = \l_in.tlbie  ? 1'h0 : _156_;
  assign _165_ = \l_in.valid  ? _159_ : r[168:165];
  assign _166_ = \l_in.valid  & _160_;
  assign _167_ = \l_in.valid  & _161_;
  assign _168_ = \l_in.valid  ? _164_ : 1'h0;
  assign _169_ = ~ \l_in.sprn [8];
  assign _170_ = _169_ ? r[132:69] : \l_in.rs ;
  assign _171_ = _169_ ? \l_in.rs [31:0] : r[164:133];
  assign _172_ = _169_ ? _143_ : 1'h0;
  assign _173_ = \l_in.valid  ? _145_ : r[365];
  assign _174_ = _169_ ? _173_ : 1'h0;
  assign _175_ = \l_in.valid  ? _158_ : 1'h0;
  assign _176_ = \l_in.mtspr  ? { 4'h1, _171_, _170_, 1'h1 } : { _165_, r[164:69], _175_ };
  assign _177_ = \l_in.mtspr  ? _172_ : _143_;
  assign _178_ = \l_in.mtspr  ? 1'h0 : _144_;
  assign _179_ = \l_in.valid  ? _145_ : r[365];
  assign _180_ = \l_in.mtspr  ? _174_ : _179_;
  assign _181_ = \l_in.valid  ? { \l_in.addr , \l_in.priv , _137_, \l_in.iside , _157_ } : { r[67:1], 1'h0 };
  assign _182_ = \l_in.valid  ? _163_ : { 1'h0, _135_[62:61], _135_[7:5] };
  assign _183_ = r[168:165] == 4'h0;
  assign _184_ = r[168:165] == 4'h1;
  assign _185_ = \d_in.done  ? 4'hc : r[168:165];
  assign _186_ = r[168:165] == 4'h2;
  assign _187_ = r[168:165] == 4'h3;
  assign _188_ = \d_in.done  ? 4'h5 : r[168:165];
  assign _189_ = \d_in.done  ? { 1'h1, \d_in.data [7:0], \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], \d_in.data [63:56] } : r[235:171];
  assign _190_ = r[168:165] == 4'h4;
  assign _191_ = r[168:165] == 4'h5;
  assign _192_ = r[168:165] == 4'h6;
  assign _193_ = r[67] ? r[300:236] : { 1'h1, \d_in.data [7:0], \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], \d_in.data [63:56] };
  assign _194_ = r[67] ? { 1'h1, \d_in.data [7:0], \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], \d_in.data [63:56] } : r[365:301];
  assign _195_ = { 1'h0, \d_in.data [60:56] } == 6'h00;
  assign _196_ = _195_ ? 4'hc : 4'h8;
  assign _197_ = _200_ ? 1'h1 : 1'h0;
  assign _198_ = \d_in.done  ? _196_ : r[168:165];
  assign _199_ = \d_in.done  ? { \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], 8'h00, \d_in.data [60:56], 1'h0, \d_in.data [6:5], \d_in.data [63:61], _194_, _193_ } : r[432:236];
  assign _200_ = \d_in.done  & _195_;
  assign _201_ = \d_in.err  ? 4'hc : _198_;
  assign _202_ = \d_in.err  ? 1'h1 : 1'h0;
  assign _203_ = r[168:165] == 4'h7;
  assign _204_ = r[371:366] + 6'h13;
  assign _205_ = _204_ - { 1'h0, r[376:372] };
  assign _206_ = ~ finalmask[30:0];
  assign _207_ = r[65:35] & _206_;
  assign _208_ = | _207_;
  assign _209_ = r[67] != r[66];
  assign _210_ = _209_ | _208_;
  assign _211_ = { 1'h0, r[376:372] } < 6'h05;
  assign _212_ = { 1'h0, r[376:372] } > 6'h10;
  assign _213_ = _211_ | _212_;
  assign _214_ = r[371:366] + 6'h13;
  assign _215_ = { 1'h0, r[376:372] } > _214_;
  assign _216_ = _213_ | _215_;
  assign _217_ = _216_ ? 4'hc : 4'h9;
  assign _218_ = _216_ ? 1'h1 : 1'h0;
  assign _219_ = _210_ ? 4'hc : _217_;
  assign _220_ = _210_ ? 1'h0 : _218_;
  assign _221_ = _210_ ? 1'h1 : 1'h0;
  assign _222_ = r[168:165] == 4'h8;
  assign _223_ = r[168:165] == 4'h9;
  assign _224_ = ~ \d_in.data [59];
  assign _225_ = r[3] | _224_;
  assign _226_ = ~ r[1];
  assign _227_ = ~ r[2];
  assign _228_ = \d_in.data [58] & _227_;
  assign _229_ = \d_in.data [57] | _228_;
  assign _230_ = ~ \d_in.data [61];
  assign _231_ = \d_in.data [56] & _230_;
  assign _232_ = _226_ ? _229_ : _231_;
  assign _233_ = _225_ ? _232_ : 1'h0;
  assign _234_ = ~ r[2];
  assign _235_ = \d_in.data [63] | _234_;
  assign _236_ = \d_in.data [48] & _235_;
  assign _237_ = _233_ & _236_;
  assign _238_ = ~ _233_;
  assign _239_ = _237_ ? 4'hb : 4'hc;
  assign _240_ = _237_ ? 2'h0 : { _233_, _238_ };
  assign _241_ = { 1'h0, \d_in.data [60:56] } < 6'h05;
  assign _242_ = { 1'h0, \d_in.data [60:56] } > 6'h10;
  assign _243_ = _241_ | _242_;
  assign _244_ = { 1'h0, \d_in.data [60:56] } > r[371:366];
  assign _245_ = _243_ | _244_;
  assign _246_ = r[371:366] - { 1'h0, \d_in.data [60:56] };
  assign _247_ = _245_ ? 4'hc : 4'h9;
  assign _248_ = _245_ ? r[432:366] : { \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], 8'h00, \d_in.data [60:56], _246_ };
  assign _249_ = _245_ ? 1'h1 : 1'h0;
  assign _250_ = \d_in.data [6] ? _239_ : _247_;
  assign _251_ = \d_in.data [6] ? r[432:366] : _248_;
  assign _252_ = \d_in.data [6] ? 1'h0 : _249_;
  assign _253_ = \d_in.data [6] ? _240_ : 2'h0;
  assign _254_ = \d_in.data [7] ? _250_ : 4'hc;
  assign _255_ = \d_in.data [7] ? _251_ : r[432:366];
  assign _256_ = \d_in.data [7] ? 1'h0 : 1'h1;
  assign _257_ = \d_in.data [7] ? _252_ : 1'h0;
  assign _258_ = \d_in.data [7] ? _253_ : 2'h0;
  assign _259_ = \d_in.done  ? _254_ : r[168:165];
  assign _260_ = \d_in.done  ? _258_ : 2'h0;
  assign _261_ = \d_in.err  ? 4'hc : _259_;
  assign _262_ = \d_in.done  ? _257_ : 1'h0;
  assign _263_ = \d_in.err  ? 1'h1 : _262_;
  assign _264_ = \d_in.done  ? { _256_, \d_in.data [7:0], \d_in.data [15:8], \d_in.data [23:16], \d_in.data [31:24], \d_in.data [39:32], \d_in.data [47:40], \d_in.data [55:48], \d_in.data [63:56], _255_ } : { 1'h0, r[496:366] };
  assign _265_ = r[168:165] == 4'ha;
  assign _266_ = ~ r[1];
  assign _267_ = _266_ ? 4'h2 : 4'h0;
  assign _268_ = _266_ ? 1'h1 : 1'h0;
  assign _269_ = _266_ ? 1'h0 : 1'h1;
  assign _270_ = r[168:165] == 4'hb;
  assign _271_ = r[168:165] == 4'hc;
  function [67:0] \23539 ;
    input [67:0] a;
    input [883:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23539  = b[67:0];
      13'b???????????1?:
        \23539  = b[135:68];
      13'b??????????1??:
        \23539  = b[203:136];
      13'b?????????1???:
        \23539  = b[271:204];
      13'b????????1????:
        \23539  = b[339:272];
      13'b???????1?????:
        \23539  = b[407:340];
      13'b??????1??????:
        \23539  = b[475:408];
      13'b?????1???????:
        \23539  = b[543:476];
      13'b????1????????:
        \23539  = b[611:544];
      13'b???1?????????:
        \23539  = b[679:612];
      13'b??1??????????:
        \23539  = b[747:680];
      13'b?1???????????:
        \23539  = b[815:748];
      13'b1????????????:
        \23539  = b[883:816];
      default:
        \23539  = a;
    endcase
  endfunction
  assign _272_ = \23539 (68'hxxxxxxxxxxxxxxxxx, { r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, r[67:1], 1'h0, _181_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [96:0] \23544 ;
    input [96:0] a;
    input [1260:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23544  = b[96:0];
      13'b???????????1?:
        \23544  = b[193:97];
      13'b??????????1??:
        \23544  = b[290:194];
      13'b?????????1???:
        \23544  = b[387:291];
      13'b????????1????:
        \23544  = b[484:388];
      13'b???????1?????:
        \23544  = b[581:485];
      13'b??????1??????:
        \23544  = b[678:582];
      13'b?????1???????:
        \23544  = b[775:679];
      13'b????1????????:
        \23544  = b[872:776];
      13'b???1?????????:
        \23544  = b[969:873];
      13'b??1??????????:
        \23544  = b[1066:970];
      13'b?1???????????:
        \23544  = b[1163:1067];
      13'b1????????????:
        \23544  = b[1260:1164];
      default:
        \23544  = a;
    endcase
  endfunction
  assign _273_ = \23544 (97'hxxxxxxxxxxxxxxxxxxxxxxxxx, { r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, r[164:69], 1'h0, _176_[96:0] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [3:0] \23547 ;
    input [3:0] a;
    input [51:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23547  = b[3:0];
      13'b???????????1?:
        \23547  = b[7:4];
      13'b??????????1??:
        \23547  = b[11:8];
      13'b?????????1???:
        \23547  = b[15:12];
      13'b????????1????:
        \23547  = b[19:16];
      13'b???????1?????:
        \23547  = b[23:20];
      13'b??????1??????:
        \23547  = b[27:24];
      13'b?????1???????:
        \23547  = b[31:28];
      13'b????1????????:
        \23547  = b[35:32];
      13'b???1?????????:
        \23547  = b[39:36];
      13'b??1??????????:
        \23547  = b[43:40];
      13'b?1???????????:
        \23547  = b[47:44];
      13'b1????????????:
        \23547  = b[51:48];
      default:
        \23547  = a;
    endcase
  endfunction
  assign _274_ = \23547 (4'hx, { 4'h0, _267_, _261_, 4'ha, _219_, _201_, 8'h76, _188_, 4'h4, _185_, 4'h2, _176_[100:97] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [63:0] \23551 ;
    input [63:0] a;
    input [831:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23551  = b[63:0];
      13'b???????????1?:
        \23551  = b[127:64];
      13'b??????????1??:
        \23551  = b[191:128];
      13'b?????????1???:
        \23551  = b[255:192];
      13'b????????1????:
        \23551  = b[319:256];
      13'b???????1?????:
        \23551  = b[383:320];
      13'b??????1??????:
        \23551  = b[447:384];
      13'b?????1???????:
        \23551  = b[511:448];
      13'b????1????????:
        \23551  = b[575:512];
      13'b???1?????????:
        \23551  = b[639:576];
      13'b??1??????????:
        \23551  = b[703:640];
      13'b?1???????????:
        \23551  = b[767:704];
      13'b1????????????:
        \23551  = b[831:768];
      default:
        \23551  = a;
    endcase
  endfunction
  assign _275_ = \23551 (64'hxxxxxxxxxxxxxxxx, { r[234:171], r[234:171], r[234:171], r[234:171], r[234:171], r[234:171], r[234:171], r[234:171], _189_[63:0], r[234:171], r[234:171], r[234:171], r[234:171] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23555 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23555  = b[0:0];
      13'b???????????1?:
        \23555  = b[1:1];
      13'b??????????1??:
        \23555  = b[2:2];
      13'b?????????1???:
        \23555  = b[3:3];
      13'b????????1????:
        \23555  = b[4:4];
      13'b???????1?????:
        \23555  = b[5:5];
      13'b??????1??????:
        \23555  = b[6:6];
      13'b?????1???????:
        \23555  = b[7:7];
      13'b????1????????:
        \23555  = b[8:8];
      13'b???1?????????:
        \23555  = b[9:9];
      13'b??1??????????:
        \23555  = b[10:10];
      13'b?1???????????:
        \23555  = b[11:11];
      13'b1????????????:
        \23555  = b[12:12];
      default:
        \23555  = a;
    endcase
  endfunction
  assign _276_ = \23555 (1'hx, { r[235], r[235], r[235], r[235], r[235], r[235], r[235], r[235], _189_[64], r[235], r[235], r[235], _177_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [63:0] \23559 ;
    input [63:0] a;
    input [831:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23559  = b[63:0];
      13'b???????????1?:
        \23559  = b[127:64];
      13'b??????????1??:
        \23559  = b[191:128];
      13'b?????????1???:
        \23559  = b[255:192];
      13'b????????1????:
        \23559  = b[319:256];
      13'b???????1?????:
        \23559  = b[383:320];
      13'b??????1??????:
        \23559  = b[447:384];
      13'b?????1???????:
        \23559  = b[511:448];
      13'b????1????????:
        \23559  = b[575:512];
      13'b???1?????????:
        \23559  = b[639:576];
      13'b??1??????????:
        \23559  = b[703:640];
      13'b?1???????????:
        \23559  = b[767:704];
      13'b1????????????:
        \23559  = b[831:768];
      default:
        \23559  = a;
    endcase
  endfunction
  assign _277_ = \23559 (64'hxxxxxxxxxxxxxxxx, { r[299:236], r[299:236], r[299:236], r[299:236], r[299:236], _199_[63:0], r[299:236], r[299:236], r[299:236], r[299:236], r[299:236], r[299:236], r[299:236] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23563 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23563  = b[0:0];
      13'b???????????1?:
        \23563  = b[1:1];
      13'b??????????1??:
        \23563  = b[2:2];
      13'b?????????1???:
        \23563  = b[3:3];
      13'b????????1????:
        \23563  = b[4:4];
      13'b???????1?????:
        \23563  = b[5:5];
      13'b??????1??????:
        \23563  = b[6:6];
      13'b?????1???????:
        \23563  = b[7:7];
      13'b????1????????:
        \23563  = b[8:8];
      13'b???1?????????:
        \23563  = b[9:9];
      13'b??1??????????:
        \23563  = b[10:10];
      13'b?1???????????:
        \23563  = b[11:11];
      13'b1????????????:
        \23563  = b[12:12];
      default:
        \23563  = a;
    endcase
  endfunction
  assign _278_ = \23563 (1'hx, { r[300], r[300], r[300], r[300], r[300], _199_[64], r[300], r[300], r[300], r[300], r[300], r[300], _178_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [63:0] \23567 ;
    input [63:0] a;
    input [831:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23567  = b[63:0];
      13'b???????????1?:
        \23567  = b[127:64];
      13'b??????????1??:
        \23567  = b[191:128];
      13'b?????????1???:
        \23567  = b[255:192];
      13'b????????1????:
        \23567  = b[319:256];
      13'b???????1?????:
        \23567  = b[383:320];
      13'b??????1??????:
        \23567  = b[447:384];
      13'b?????1???????:
        \23567  = b[511:448];
      13'b????1????????:
        \23567  = b[575:512];
      13'b???1?????????:
        \23567  = b[639:576];
      13'b??1??????????:
        \23567  = b[703:640];
      13'b?1???????????:
        \23567  = b[767:704];
      13'b1????????????:
        \23567  = b[831:768];
      default:
        \23567  = a;
    endcase
  endfunction
  assign _279_ = \23567 (64'hxxxxxxxxxxxxxxxx, { r[364:301], r[364:301], r[364:301], r[364:301], r[364:301], _199_[128:65], r[364:301], r[364:301], r[364:301], r[364:301], r[364:301], r[364:301], r[364:301] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23571 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23571  = b[0:0];
      13'b???????????1?:
        \23571  = b[1:1];
      13'b??????????1??:
        \23571  = b[2:2];
      13'b?????????1???:
        \23571  = b[3:3];
      13'b????????1????:
        \23571  = b[4:4];
      13'b???????1?????:
        \23571  = b[5:5];
      13'b??????1??????:
        \23571  = b[6:6];
      13'b?????1???????:
        \23571  = b[7:7];
      13'b????1????????:
        \23571  = b[8:8];
      13'b???1?????????:
        \23571  = b[9:9];
      13'b??1??????????:
        \23571  = b[10:10];
      13'b?1???????????:
        \23571  = b[11:11];
      13'b1????????????:
        \23571  = b[12:12];
      default:
        \23571  = a;
    endcase
  endfunction
  assign _280_ = \23571 (1'hx, { r[365], r[365], r[365], r[365], r[365], _199_[129], r[365], r[365], r[365], r[365], r[365], r[365], _180_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [5:0] \23576 ;
    input [5:0] a;
    input [77:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23576  = b[5:0];
      13'b???????????1?:
        \23576  = b[11:6];
      13'b??????????1??:
        \23576  = b[17:12];
      13'b?????????1???:
        \23576  = b[23:18];
      13'b????????1????:
        \23576  = b[29:24];
      13'b???????1?????:
        \23576  = b[35:30];
      13'b??????1??????:
        \23576  = b[41:36];
      13'b?????1???????:
        \23576  = b[47:42];
      13'b????1????????:
        \23576  = b[53:48];
      13'b???1?????????:
        \23576  = b[59:54];
      13'b??1??????????:
        \23576  = b[65:60];
      13'b?1???????????:
        \23576  = b[71:66];
      13'b1????????????:
        \23576  = b[77:72];
      default:
        \23576  = a;
    endcase
  endfunction
  assign _281_ = \23576 (6'hxx, { r[371:366], r[371:366], _264_[5:0], r[371:366], _205_, _199_[135:130], r[371:366], 1'h0, r[175:171], r[371:366], r[371:366], r[371:366], r[371:366], _182_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [4:0] \23581 ;
    input [4:0] a;
    input [64:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23581  = b[4:0];
      13'b???????????1?:
        \23581  = b[9:5];
      13'b??????????1??:
        \23581  = b[14:10];
      13'b?????????1???:
        \23581  = b[19:15];
      13'b????????1????:
        \23581  = b[24:20];
      13'b???????1?????:
        \23581  = b[29:25];
      13'b??????1??????:
        \23581  = b[34:30];
      13'b?????1???????:
        \23581  = b[39:35];
      13'b????1????????:
        \23581  = b[44:40];
      13'b???1?????????:
        \23581  = b[49:45];
      13'b??1??????????:
        \23581  = b[54:50];
      13'b?1???????????:
        \23581  = b[59:55];
      13'b1????????????:
        \23581  = b[64:60];
      default:
        \23581  = a;
    endcase
  endfunction
  assign _282_ = \23581 (5'hxx, { r[376:372], r[376:372], _264_[10:6], r[376:372], r[376:372], _199_[140:136], r[376:372], r[376:372], r[376:372], r[376:372], r[376:372], r[376:372], _135_[4:0] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [55:0] \23586 ;
    input [55:0] a;
    input [727:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23586  = b[55:0];
      13'b???????????1?:
        \23586  = b[111:56];
      13'b??????????1??:
        \23586  = b[167:112];
      13'b?????????1???:
        \23586  = b[223:168];
      13'b????????1????:
        \23586  = b[279:224];
      13'b???????1?????:
        \23586  = b[335:280];
      13'b??????1??????:
        \23586  = b[391:336];
      13'b?????1???????:
        \23586  = b[447:392];
      13'b????1????????:
        \23586  = b[503:448];
      13'b???1?????????:
        \23586  = b[559:504];
      13'b??1??????????:
        \23586  = b[615:560];
      13'b?1???????????:
        \23586  = b[671:616];
      13'b1????????????:
        \23586  = b[727:672];
      default:
        \23586  = a;
    endcase
  endfunction
  assign _283_ = \23586 (56'hxxxxxxxxxxxxxx, { r[432:377], r[432:377], _264_[66:11], r[432:377], r[432:377], _199_[196:141], r[432:377], r[432:377], r[432:377], r[432:377], r[432:377], r[432:377], _135_[55:8], 8'h00 }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [63:0] \23590 ;
    input [63:0] a;
    input [831:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23590  = b[63:0];
      13'b???????????1?:
        \23590  = b[127:64];
      13'b??????????1??:
        \23590  = b[191:128];
      13'b?????????1???:
        \23590  = b[255:192];
      13'b????????1????:
        \23590  = b[319:256];
      13'b???????1?????:
        \23590  = b[383:320];
      13'b??????1??????:
        \23590  = b[447:384];
      13'b?????1???????:
        \23590  = b[511:448];
      13'b????1????????:
        \23590  = b[575:512];
      13'b???1?????????:
        \23590  = b[639:576];
      13'b??1??????????:
        \23590  = b[703:640];
      13'b?1???????????:
        \23590  = b[767:704];
      13'b1????????????:
        \23590  = b[831:768];
      default:
        \23590  = a;
    endcase
  endfunction
  assign _284_ = \23590 (64'hxxxxxxxxxxxxxxxx, { r[496:433], r[496:433], _264_[130:67], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433], r[496:433] }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23593 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23593  = b[0:0];
      13'b???????????1?:
        \23593  = b[1:1];
      13'b??????????1??:
        \23593  = b[2:2];
      13'b?????????1???:
        \23593  = b[3:3];
      13'b????????1????:
        \23593  = b[4:4];
      13'b???????1?????:
        \23593  = b[5:5];
      13'b??????1??????:
        \23593  = b[6:6];
      13'b?????1???????:
        \23593  = b[7:7];
      13'b????1????????:
        \23593  = b[8:8];
      13'b???1?????????:
        \23593  = b[9:9];
      13'b??1??????????:
        \23593  = b[10:10];
      13'b?1???????????:
        \23593  = b[11:11];
      13'b1????????????:
        \23593  = b[12:12];
      default:
        \23593  = a;
    endcase
  endfunction
  assign _285_ = \23593 (1'hx, { 2'h0, _264_[131], 2'h0, _197_, 6'h00, _168_ }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23595 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23595  = b[0:0];
      13'b???????????1?:
        \23595  = b[1:1];
      13'b??????????1??:
        \23595  = b[2:2];
      13'b?????????1???:
        \23595  = b[3:3];
      13'b????????1????:
        \23595  = b[4:4];
      13'b???????1?????:
        \23595  = b[5:5];
      13'b??????1??????:
        \23595  = b[6:6];
      13'b?????1???????:
        \23595  = b[7:7];
      13'b????1????????:
        \23595  = b[8:8];
      13'b???1?????????:
        \23595  = b[9:9];
      13'b??1??????????:
        \23595  = b[10:10];
      13'b?1???????????:
        \23595  = b[11:11];
      13'b1????????????:
        \23595  = b[12:12];
      default:
        \23595  = a;
    endcase
  endfunction
  assign _286_ = \23595 (1'hx, { 2'h0, _263_, 1'h0, _220_, _202_, 7'h00 }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23597 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23597  = b[0:0];
      13'b???????????1?:
        \23597  = b[1:1];
      13'b??????????1??:
        \23597  = b[2:2];
      13'b?????????1???:
        \23597  = b[3:3];
      13'b????????1????:
        \23597  = b[4:4];
      13'b???????1?????:
        \23597  = b[5:5];
      13'b??????1??????:
        \23597  = b[6:6];
      13'b?????1???????:
        \23597  = b[7:7];
      13'b????1????????:
        \23597  = b[8:8];
      13'b???1?????????:
        \23597  = b[9:9];
      13'b??1??????????:
        \23597  = b[10:10];
      13'b?1???????????:
        \23597  = b[11:11];
      13'b1????????????:
        \23597  = b[12:12];
      default:
        \23597  = a;
    endcase
  endfunction
  assign _287_ = \23597 (1'hx, { 4'h0, _221_, 8'h00 }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [1:0] \23600 ;
    input [1:0] a;
    input [25:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23600  = b[1:0];
      13'b???????????1?:
        \23600  = b[3:2];
      13'b??????????1??:
        \23600  = b[5:4];
      13'b?????????1???:
        \23600  = b[7:6];
      13'b????????1????:
        \23600  = b[9:8];
      13'b???????1?????:
        \23600  = b[11:10];
      13'b??????1??????:
        \23600  = b[13:12];
      13'b?????1???????:
        \23600  = b[15:14];
      13'b????1????????:
        \23600  = b[17:16];
      13'b???1?????????:
        \23600  = b[19:18];
      13'b??1??????????:
        \23600  = b[21:20];
      13'b?1???????????:
        \23600  = b[23:22];
      13'b1????????????:
        \23600  = b[25:24];
      default:
        \23600  = a;
    endcase
  endfunction
  assign _288_ = \23600 (2'hx, { 4'h0, _260_, 20'h00000 }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23617 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23617  = b[0:0];
      13'b???????????1?:
        \23617  = b[1:1];
      13'b??????????1??:
        \23617  = b[2:2];
      13'b?????????1???:
        \23617  = b[3:3];
      13'b????????1????:
        \23617  = b[4:4];
      13'b???????1?????:
        \23617  = b[5:5];
      13'b??????1??????:
        \23617  = b[6:6];
      13'b?????1???????:
        \23617  = b[7:7];
      13'b????1????????:
        \23617  = b[8:8];
      13'b???1?????????:
        \23617  = b[9:9];
      13'b??1??????????:
        \23617  = b[10:10];
      13'b?1???????????:
        \23617  = b[11:11];
      13'b1????????????:
        \23617  = b[12:12];
      default:
        \23617  = a;
    endcase
  endfunction
  assign _289_ = \23617 (1'hx, { 1'h0, _268_, 11'h24a }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23622 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23622  = b[0:0];
      13'b???????????1?:
        \23622  = b[1:1];
      13'b??????????1??:
        \23622  = b[2:2];
      13'b?????????1???:
        \23622  = b[3:3];
      13'b????????1????:
        \23622  = b[4:4];
      13'b???????1?????:
        \23622  = b[5:5];
      13'b??????1??????:
        \23622  = b[6:6];
      13'b?????1???????:
        \23622  = b[7:7];
      13'b????1????????:
        \23622  = b[8:8];
      13'b???1?????????:
        \23622  = b[9:9];
      13'b??1??????????:
        \23622  = b[10:10];
      13'b?1???????????:
        \23622  = b[11:11];
      13'b1????????????:
        \23622  = b[12:12];
      default:
        \23622  = a;
    endcase
  endfunction
  assign _290_ = \23622 (1'hx, 13'h0800, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23626 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23626  = b[0:0];
      13'b???????????1?:
        \23626  = b[1:1];
      13'b??????????1??:
        \23626  = b[2:2];
      13'b?????????1???:
        \23626  = b[3:3];
      13'b????????1????:
        \23626  = b[4:4];
      13'b???????1?????:
        \23626  = b[5:5];
      13'b??????1??????:
        \23626  = b[6:6];
      13'b?????1???????:
        \23626  = b[7:7];
      13'b????1????????:
        \23626  = b[8:8];
      13'b???1?????????:
        \23626  = b[9:9];
      13'b??1??????????:
        \23626  = b[10:10];
      13'b?1???????????:
        \23626  = b[11:11];
      13'b1????????????:
        \23626  = b[12:12];
      default:
        \23626  = a;
    endcase
  endfunction
  assign _291_ = \23626 (1'hx, { 1'h0, _269_, 11'h000 }, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23631 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23631  = b[0:0];
      13'b???????????1?:
        \23631  = b[1:1];
      13'b??????????1??:
        \23631  = b[2:2];
      13'b?????????1???:
        \23631  = b[3:3];
      13'b????????1????:
        \23631  = b[4:4];
      13'b???????1?????:
        \23631  = b[5:5];
      13'b??????1??????:
        \23631  = b[6:6];
      13'b?????1???????:
        \23631  = b[7:7];
      13'b????1????????:
        \23631  = b[8:8];
      13'b???1?????????:
        \23631  = b[9:9];
      13'b??1??????????:
        \23631  = b[10:10];
      13'b?1???????????:
        \23631  = b[11:11];
      13'b1????????????:
        \23631  = b[12:12];
      default:
        \23631  = a;
    endcase
  endfunction
  assign _292_ = \23631 (1'hx, 13'h0002, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23636 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23636  = b[0:0];
      13'b???????????1?:
        \23636  = b[1:1];
      13'b??????????1??:
        \23636  = b[2:2];
      13'b?????????1???:
        \23636  = b[3:3];
      13'b????????1????:
        \23636  = b[4:4];
      13'b???????1?????:
        \23636  = b[5:5];
      13'b??????1??????:
        \23636  = b[6:6];
      13'b?????1???????:
        \23636  = b[7:7];
      13'b????1????????:
        \23636  = b[8:8];
      13'b???1?????????:
        \23636  = b[9:9];
      13'b??1??????????:
        \23636  = b[10:10];
      13'b?1???????????:
        \23636  = b[11:11];
      13'b1????????????:
        \23636  = b[12:12];
      default:
        \23636  = a;
    endcase
  endfunction
  assign _293_ = \23636 (1'hx, 13'h0008, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  function [0:0] \23641 ;
    input [0:0] a;
    input [12:0] b;
    input [12:0] s;
    (* parallel_case *)
    casez (s)
      13'b????????????1:
        \23641  = b[0:0];
      13'b???????????1?:
        \23641  = b[1:1];
      13'b??????????1??:
        \23641  = b[2:2];
      13'b?????????1???:
        \23641  = b[3:3];
      13'b????????1????:
        \23641  = b[4:4];
      13'b???????1?????:
        \23641  = b[5:5];
      13'b??????1??????:
        \23641  = b[6:6];
      13'b?????1???????:
        \23641  = b[7:7];
      13'b????1????????:
        \23641  = b[8:8];
      13'b???1?????????:
        \23641  = b[9:9];
      13'b??1??????????:
        \23641  = b[10:10];
      13'b?1???????????:
        \23641  = b[11:11];
      13'b1????????????:
        \23641  = b[12:12];
      default:
        \23641  = a;
    endcase
  endfunction
  assign _294_ = \23641 (1'hx, 13'h0040, { _271_, _270_, _265_, _223_, _222_, _203_, _192_, _191_, _190_, _187_, _186_, _184_, _183_ });
  assign _295_ = _274_ == 4'hc;
  assign _296_ = _274_ == 4'hb;
  assign _297_ = _296_ & r[1];
  assign _298_ = _295_ | _297_;
  assign _299_ = _285_ | _286_;
  assign _300_ = _299_ | _287_;
  assign _301_ = _300_ | _288_[0];
  assign _302_ = _301_ | _288_[1];
  assign _303_ = ~ _302_;
  assign _304_ = _298_ ? { _302_, _303_ } : 2'h0;
  assign _305_ = r[67] ? 32'd0 : r[164:133];
  assign _306_ = ~ finalmask[23:0];
  assign _307_ = r[206:183] & _306_;
  assign _308_ = _305_[31:8] & finalmask[23:0];
  assign _309_ = _307_ | _308_;
  assign _310_ = ~ mask;
  assign _311_ = r[395:380] & _310_;
  assign _312_ = addrsh & mask;
  assign _313_ = _311_ | _312_;
  assign _314_ = ~ finalmask;
  assign _315_ = r[488:445] & _314_;
  assign _316_ = r[59:16] & finalmask;
  assign _317_ = _315_ | _316_;
  assign _318_ = _294_ ? { 8'h00, r[226:207], _309_, _305_[7:0], 4'h0 } : { 8'h00, r[432:396], _313_, 3'h0 };
  assign _319_ = _293_ ? { 8'h00, r[124:81], 12'h008 } : _318_;
  assign _320_ = _290_ ? { 8'h00, _317_, r[444:433] } : 64'h0000000000000000;
  assign _321_ = _290_ ? { r[67:16], 12'h000 } : _319_;
  assign _322_ = _292_ ? 64'h0000000000000000 : _320_;
  assign _323_ = _292_ ? r[67:4] : _321_;
  assign r = _011_;
  assign rin = { _288_, _287_, _286_, _285_, _284_, _283_, _282_, _281_, _280_, _279_, _278_, _277_, _276_, _275_, _304_, _274_, _273_, _272_ };
  assign addrsh = _022_;
  assign mask = { _044_, _042_, _040_, _038_, _036_, _034_, _032_, _030_, _028_, _026_, _024_, 5'h1f };
  assign finalmask = { _132_, _130_, _128_, _126_, _124_, _122_, _120_, _118_, _116_, _114_, _112_, _110_, _108_, _106_, _104_, _102_, _100_, _098_, _096_, _094_, _092_, _090_, _088_, _086_, _084_, _082_, _080_, _078_, _076_, _074_, _072_, _070_, _068_, _066_, _064_, _062_, _060_, _058_, _056_, _054_, _052_, _050_, _048_, _046_ };
  assign \l_out.done  = r[169];
  assign \l_out.err  = r[170];
  assign \l_out.invalid  = r[497];
  assign \l_out.badtree  = r[498];
  assign \l_out.segerr  = r[499];
  assign \l_out.perm_error  = r[500];
  assign \l_out.rc_error  = r[501];
  assign \l_out.sprval  = _000_;
  assign \d_out.valid  = _289_;
  assign \d_out.tlbie  = _292_;
  assign \d_out.doall  = r[68];
  assign \d_out.tlbld  = _290_;
  assign \d_out.addr  = _323_;
  assign \d_out.pte  = _322_;
  assign \i_out.tlbld  = _291_;
  assign \i_out.tlbie  = _292_;
  assign \i_out.doall  = r[68];
  assign \i_out.addr  = _323_;
  assign \i_out.pte  = _322_;
endmodule