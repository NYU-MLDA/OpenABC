module logical(rs, rb, op, invert_in, invert_out, datalen, result);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire [63:0] _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire [15:0] _0913_;
  wire _0914_;
  wire [7:0] _0915_;
  wire _0916_;
  wire [7:0] _0917_;
  wire [7:0] _0918_;
  wire [15:0] _0919_;
  wire [31:0] _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire [5:0] _1099_;
  wire _1100_;
  wire _1101_;
  wire [5:0] _1102_;
  wire _1103_;
  wire _1104_;
  wire [5:0] _1105_;
  wire _1106_;
  wire _1107_;
  wire [5:0] _1108_;
  wire _1109_;
  wire _1110_;
  wire [5:0] _1111_;
  wire _1112_;
  wire _1113_;
  wire [5:0] _1114_;
  wire _1115_;
  wire _1116_;
  wire [5:0] _1117_;
  wire _1118_;
  wire _1119_;
  wire [5:0] _1120_;
  wire _1121_;
  wire [63:0] _1122_;
  wire [63:0] _1123_;
  wire [63:0] _1124_;
  wire _1125_;
  wire [63:0] _1126_;
  wire _1127_;
  wire [63:0] _1128_;
  wire [63:0] _1129_;
  wire [63:0] _1130_;
  wire [63:0] _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire [7:0] _1139_;
  wire _1140_;
  wire [7:0] _1141_;
  wire _1142_;
  wire [7:0] _1143_;
  wire _1144_;
  wire [7:0] _1145_;
  wire _1146_;
  wire [7:0] _1147_;
  wire _1148_;
  wire [7:0] _1149_;
  wire _1150_;
  wire [7:0] _1151_;
  wire _1152_;
  wire [7:0] _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  input [3:0] datalen;
  wire [3:0] datalen;
  input invert_in;
  wire invert_in;
  input invert_out;
  wire invert_out;
  input [5:0] op;
  wire [5:0] op;
  wire par0;
  wire par1;
  wire [63:0] parity;
  wire [7:0] permute;
  input [63:0] rb;
  wire [63:0] rb;
  output [63:0] result;
  wire [63:0] result;
  input [63:0] rs;
  wire [63:0] rs;
  assign _0000_ = _1099_[0] ? rb[1] : rb[0];
  assign _0001_ = _1099_[0] ? rb[5] : rb[4];
  assign _0002_ = _1099_[0] ? rb[9] : rb[8];
  assign _0003_ = _1099_[0] ? rb[13] : rb[12];
  assign _0004_ = _1099_[0] ? rb[17] : rb[16];
  assign _0005_ = _1099_[0] ? rb[21] : rb[20];
  assign _0006_ = _1099_[0] ? rb[25] : rb[24];
  assign _0007_ = _1099_[0] ? rb[29] : rb[28];
  assign _0008_ = _1099_[0] ? rb[33] : rb[32];
  assign _0009_ = _1099_[0] ? rb[37] : rb[36];
  assign _0010_ = _1099_[0] ? rb[41] : rb[40];
  assign _0011_ = _1099_[0] ? rb[45] : rb[44];
  assign _0012_ = _1099_[0] ? rb[49] : rb[48];
  assign _0013_ = _1099_[0] ? rb[53] : rb[52];
  assign _0014_ = _1099_[0] ? rb[57] : rb[56];
  assign _0015_ = _1099_[0] ? rb[61] : rb[60];
  assign _0016_ = _1099_[2] ? _0922_ : _0921_;
  assign _0017_ = _1099_[2] ? _0926_ : _0925_;
  assign _0018_ = _1099_[2] ? _0930_ : _0929_;
  assign _0019_ = _1099_[2] ? _0934_ : _0933_;
  assign _0020_ = _1099_[4] ? _0938_ : _0937_;
  assign _0021_ = _1102_[0] ? rb[1] : rb[0];
  assign _0022_ = _1102_[0] ? rb[5] : rb[4];
  assign _0023_ = _1102_[0] ? rb[9] : rb[8];
  assign _0024_ = _1102_[0] ? rb[13] : rb[12];
  assign _0025_ = _1102_[0] ? rb[17] : rb[16];
  assign _0026_ = _1102_[0] ? rb[21] : rb[20];
  assign _0027_ = _1102_[0] ? rb[25] : rb[24];
  assign _0028_ = _1102_[0] ? rb[29] : rb[28];
  assign _0029_ = _1102_[0] ? rb[33] : rb[32];
  assign _0030_ = _1102_[0] ? rb[37] : rb[36];
  assign _0031_ = _1102_[0] ? rb[41] : rb[40];
  assign _0032_ = _1102_[0] ? rb[45] : rb[44];
  assign _0033_ = _1102_[0] ? rb[49] : rb[48];
  assign _0034_ = _1102_[0] ? rb[53] : rb[52];
  assign _0035_ = _1102_[0] ? rb[57] : rb[56];
  assign _0036_ = _1102_[0] ? rb[61] : rb[60];
  assign _0037_ = _1102_[2] ? _0943_ : _0942_;
  assign _0038_ = _1102_[2] ? _0947_ : _0946_;
  assign _0039_ = _1102_[2] ? _0951_ : _0950_;
  assign _0040_ = _1102_[2] ? _0955_ : _0954_;
  assign _0041_ = _1102_[4] ? _0959_ : _0958_;
  assign _0042_ = _1105_[0] ? rb[1] : rb[0];
  assign _0043_ = _1105_[0] ? rb[5] : rb[4];
  assign _0044_ = _1105_[0] ? rb[9] : rb[8];
  assign _0045_ = _1105_[0] ? rb[13] : rb[12];
  assign _0046_ = _1105_[0] ? rb[17] : rb[16];
  assign _0047_ = _1105_[0] ? rb[21] : rb[20];
  assign _0048_ = _1105_[0] ? rb[25] : rb[24];
  assign _0049_ = _1105_[0] ? rb[29] : rb[28];
  assign _0050_ = _1105_[0] ? rb[33] : rb[32];
  assign _0051_ = _1105_[0] ? rb[37] : rb[36];
  assign _0052_ = _1105_[0] ? rb[41] : rb[40];
  assign _0053_ = _1105_[0] ? rb[45] : rb[44];
  assign _0054_ = _1105_[0] ? rb[49] : rb[48];
  assign _0055_ = _1105_[0] ? rb[53] : rb[52];
  assign _0056_ = _1105_[0] ? rb[57] : rb[56];
  assign _0057_ = _1105_[0] ? rb[61] : rb[60];
  assign _0058_ = _1105_[2] ? _0964_ : _0963_;
  assign _0059_ = _1105_[2] ? _0968_ : _0967_;
  assign _0060_ = _1105_[2] ? _0972_ : _0971_;
  assign _0061_ = _1105_[2] ? _0976_ : _0975_;
  assign _0062_ = _1105_[4] ? _0980_ : _0979_;
  assign _0063_ = _1108_[0] ? rb[1] : rb[0];
  assign _0064_ = _1108_[0] ? rb[5] : rb[4];
  assign _0065_ = _1108_[0] ? rb[9] : rb[8];
  assign _0066_ = _1108_[0] ? rb[13] : rb[12];
  assign _0067_ = _1108_[0] ? rb[17] : rb[16];
  assign _0068_ = _1108_[0] ? rb[21] : rb[20];
  assign _0069_ = _1108_[0] ? rb[25] : rb[24];
  assign _0070_ = _1108_[0] ? rb[29] : rb[28];
  assign _0071_ = _1108_[0] ? rb[33] : rb[32];
  assign _0072_ = _1108_[0] ? rb[37] : rb[36];
  assign _0073_ = _1108_[0] ? rb[41] : rb[40];
  assign _0074_ = _1108_[0] ? rb[45] : rb[44];
  assign _0075_ = _1108_[0] ? rb[49] : rb[48];
  assign _0076_ = _1108_[0] ? rb[53] : rb[52];
  assign _0077_ = _1108_[0] ? rb[57] : rb[56];
  assign _0078_ = _1108_[0] ? rb[61] : rb[60];
  assign _0079_ = _1108_[2] ? _0985_ : _0984_;
  assign _0080_ = _1108_[2] ? _0989_ : _0988_;
  assign _0081_ = _1108_[2] ? _0993_ : _0992_;
  assign _0082_ = _1108_[2] ? _0997_ : _0996_;
  assign _0083_ = _1108_[4] ? _1001_ : _1000_;
  assign _0084_ = _1111_[0] ? rb[1] : rb[0];
  assign _0085_ = _1111_[0] ? rb[5] : rb[4];
  assign _0086_ = _1111_[0] ? rb[9] : rb[8];
  assign _0087_ = _1111_[0] ? rb[13] : rb[12];
  assign _0088_ = _1111_[0] ? rb[17] : rb[16];
  assign _0089_ = _1111_[0] ? rb[21] : rb[20];
  assign _0090_ = _1111_[0] ? rb[25] : rb[24];
  assign _0091_ = _1111_[0] ? rb[29] : rb[28];
  assign _0092_ = _1111_[0] ? rb[33] : rb[32];
  assign _0093_ = _1111_[0] ? rb[37] : rb[36];
  assign _0094_ = _1111_[0] ? rb[41] : rb[40];
  assign _0095_ = _1111_[0] ? rb[45] : rb[44];
  assign _0096_ = _1111_[0] ? rb[49] : rb[48];
  assign _0097_ = _1111_[0] ? rb[53] : rb[52];
  assign _0098_ = _1111_[0] ? rb[57] : rb[56];
  assign _0099_ = _1111_[0] ? rb[61] : rb[60];
  assign _0100_ = _1111_[2] ? _1006_ : _1005_;
  assign _0101_ = _1111_[2] ? _1010_ : _1009_;
  assign _0102_ = _1111_[2] ? _1014_ : _1013_;
  assign _0103_ = _1111_[2] ? _1018_ : _1017_;
  assign _0104_ = _1111_[4] ? _1022_ : _1021_;
  assign _0105_ = _1114_[0] ? rb[1] : rb[0];
  assign _0106_ = _1114_[0] ? rb[5] : rb[4];
  assign _0107_ = _1114_[0] ? rb[9] : rb[8];
  assign _0108_ = _1114_[0] ? rb[13] : rb[12];
  assign _0109_ = _1114_[0] ? rb[17] : rb[16];
  assign _0110_ = _1114_[0] ? rb[21] : rb[20];
  assign _0111_ = _1114_[0] ? rb[25] : rb[24];
  assign _0112_ = _1114_[0] ? rb[29] : rb[28];
  assign _0113_ = _1114_[0] ? rb[33] : rb[32];
  assign _0114_ = _1114_[0] ? rb[37] : rb[36];
  assign _0115_ = _1114_[0] ? rb[41] : rb[40];
  assign _0116_ = _1114_[0] ? rb[45] : rb[44];
  assign _0117_ = _1114_[0] ? rb[49] : rb[48];
  assign _0118_ = _1114_[0] ? rb[53] : rb[52];
  assign _0119_ = _1114_[0] ? rb[57] : rb[56];
  assign _0120_ = _1114_[0] ? rb[61] : rb[60];
  assign _0121_ = _1114_[2] ? _1027_ : _1026_;
  assign _0122_ = _1114_[2] ? _1031_ : _1030_;
  assign _0123_ = _1114_[2] ? _1035_ : _1034_;
  assign _0124_ = _1114_[2] ? _1039_ : _1038_;
  assign _0125_ = _1114_[4] ? _1043_ : _1042_;
  assign _0126_ = _1117_[0] ? rb[1] : rb[0];
  assign _0127_ = _1117_[0] ? rb[5] : rb[4];
  assign _0128_ = _1117_[0] ? rb[9] : rb[8];
  assign _0129_ = _1117_[0] ? rb[13] : rb[12];
  assign _0130_ = _1117_[0] ? rb[17] : rb[16];
  assign _0131_ = _1117_[0] ? rb[21] : rb[20];
  assign _0132_ = _1117_[0] ? rb[25] : rb[24];
  assign _0133_ = _1117_[0] ? rb[29] : rb[28];
  assign _0134_ = _1117_[0] ? rb[33] : rb[32];
  assign _0135_ = _1117_[0] ? rb[37] : rb[36];
  assign _0136_ = _1117_[0] ? rb[41] : rb[40];
  assign _0137_ = _1117_[0] ? rb[45] : rb[44];
  assign _0138_ = _1117_[0] ? rb[49] : rb[48];
  assign _0139_ = _1117_[0] ? rb[53] : rb[52];
  assign _0140_ = _1117_[0] ? rb[57] : rb[56];
  assign _0141_ = _1117_[0] ? rb[61] : rb[60];
  assign _0142_ = _1117_[2] ? _1048_ : _1047_;
  assign _0143_ = _1117_[2] ? _1052_ : _1051_;
  assign _0144_ = _1117_[2] ? _1056_ : _1055_;
  assign _0145_ = _1117_[2] ? _1060_ : _1059_;
  assign _0146_ = _1117_[4] ? _1064_ : _1063_;
  assign _0147_ = _1120_[0] ? rb[1] : rb[0];
  assign _0148_ = _1120_[0] ? rb[5] : rb[4];
  assign _0149_ = _1120_[0] ? rb[9] : rb[8];
  assign _0150_ = _1120_[0] ? rb[13] : rb[12];
  assign _0151_ = _1120_[0] ? rb[17] : rb[16];
  assign _0152_ = _1120_[0] ? rb[21] : rb[20];
  assign _0153_ = _1120_[0] ? rb[25] : rb[24];
  assign _0154_ = _1120_[0] ? rb[29] : rb[28];
  assign _0155_ = _1120_[0] ? rb[33] : rb[32];
  assign _0156_ = _1120_[0] ? rb[37] : rb[36];
  assign _0157_ = _1120_[0] ? rb[41] : rb[40];
  assign _0158_ = _1120_[0] ? rb[45] : rb[44];
  assign _0159_ = _1120_[0] ? rb[49] : rb[48];
  assign _0160_ = _1120_[0] ? rb[53] : rb[52];
  assign _0161_ = _1120_[0] ? rb[57] : rb[56];
  assign _0162_ = _1120_[0] ? rb[61] : rb[60];
  assign _0163_ = _1120_[2] ? _1069_ : _1068_;
  assign _0164_ = _1120_[2] ? _1073_ : _1072_;
  assign _0165_ = _1120_[2] ? _1077_ : _1076_;
  assign _0166_ = _1120_[2] ? _1081_ : _1080_;
  assign _0167_ = _1120_[4] ? _1085_ : _1084_;
  assign _0168_ = _1099_[0] ? rb[3] : rb[2];
  assign _0169_ = _1099_[0] ? rb[7] : rb[6];
  assign _0170_ = _1099_[0] ? rb[11] : rb[10];
  assign _0171_ = _1099_[0] ? rb[15] : rb[14];
  assign _0172_ = _1099_[0] ? rb[19] : rb[18];
  assign _0173_ = _1099_[0] ? rb[23] : rb[22];
  assign _0174_ = _1099_[0] ? rb[27] : rb[26];
  assign _0175_ = _1099_[0] ? rb[31] : rb[30];
  assign _0176_ = _1099_[0] ? rb[35] : rb[34];
  assign _0177_ = _1099_[0] ? rb[39] : rb[38];
  assign _0178_ = _1099_[0] ? rb[43] : rb[42];
  assign _0179_ = _1099_[0] ? rb[47] : rb[46];
  assign _0180_ = _1099_[0] ? rb[51] : rb[50];
  assign _0181_ = _1099_[0] ? rb[55] : rb[54];
  assign _0182_ = _1099_[0] ? rb[59] : rb[58];
  assign _0183_ = _1099_[0] ? rb[63] : rb[62];
  assign _0184_ = _1099_[2] ? _0924_ : _0923_;
  assign _0185_ = _1099_[2] ? _0928_ : _0927_;
  assign _0186_ = _1099_[2] ? _0932_ : _0931_;
  assign _0187_ = _1099_[2] ? _0936_ : _0935_;
  assign _0188_ = _1099_[4] ? _0940_ : _0939_;
  assign _0189_ = _1102_[0] ? rb[3] : rb[2];
  assign _0190_ = _1102_[0] ? rb[7] : rb[6];
  assign _0191_ = _1102_[0] ? rb[11] : rb[10];
  assign _0192_ = _1102_[0] ? rb[15] : rb[14];
  assign _0193_ = _1102_[0] ? rb[19] : rb[18];
  assign _0194_ = _1102_[0] ? rb[23] : rb[22];
  assign _0195_ = _1102_[0] ? rb[27] : rb[26];
  assign _0196_ = _1102_[0] ? rb[31] : rb[30];
  assign _0197_ = _1102_[0] ? rb[35] : rb[34];
  assign _0198_ = _1102_[0] ? rb[39] : rb[38];
  assign _0199_ = _1102_[0] ? rb[43] : rb[42];
  assign _0200_ = _1102_[0] ? rb[47] : rb[46];
  assign _0201_ = _1102_[0] ? rb[51] : rb[50];
  assign _0202_ = _1102_[0] ? rb[55] : rb[54];
  assign _0203_ = _1102_[0] ? rb[59] : rb[58];
  assign _0204_ = _1102_[0] ? rb[63] : rb[62];
  assign _0205_ = _1102_[2] ? _0945_ : _0944_;
  assign _0206_ = _1102_[2] ? _0949_ : _0948_;
  assign _0207_ = _1102_[2] ? _0953_ : _0952_;
  assign _0208_ = _1102_[2] ? _0957_ : _0956_;
  assign _0209_ = _1102_[4] ? _0961_ : _0960_;
  assign _0210_ = _1105_[0] ? rb[3] : rb[2];
  assign _0211_ = _1105_[0] ? rb[7] : rb[6];
  assign _0212_ = _1105_[0] ? rb[11] : rb[10];
  assign _0213_ = _1105_[0] ? rb[15] : rb[14];
  assign _0214_ = _1105_[0] ? rb[19] : rb[18];
  assign _0215_ = _1105_[0] ? rb[23] : rb[22];
  assign _0216_ = _1105_[0] ? rb[27] : rb[26];
  assign _0217_ = _1105_[0] ? rb[31] : rb[30];
  assign _0218_ = _1105_[0] ? rb[35] : rb[34];
  assign _0219_ = _1105_[0] ? rb[39] : rb[38];
  assign _0220_ = _1105_[0] ? rb[43] : rb[42];
  assign _0221_ = _1105_[0] ? rb[47] : rb[46];
  assign _0222_ = _1105_[0] ? rb[51] : rb[50];
  assign _0223_ = _1105_[0] ? rb[55] : rb[54];
  assign _0224_ = _1105_[0] ? rb[59] : rb[58];
  assign _0225_ = _1105_[0] ? rb[63] : rb[62];
  assign _0226_ = _1105_[2] ? _0966_ : _0965_;
  assign _0227_ = _1105_[2] ? _0970_ : _0969_;
  assign _0228_ = _1105_[2] ? _0974_ : _0973_;
  assign _0229_ = _1105_[2] ? _0978_ : _0977_;
  assign _0230_ = _1105_[4] ? _0982_ : _0981_;
  assign _0231_ = _1108_[0] ? rb[3] : rb[2];
  assign _0232_ = _1108_[0] ? rb[7] : rb[6];
  assign _0233_ = _1108_[0] ? rb[11] : rb[10];
  assign _0234_ = _1108_[0] ? rb[15] : rb[14];
  assign _0235_ = _1108_[0] ? rb[19] : rb[18];
  assign _0236_ = _1108_[0] ? rb[23] : rb[22];
  assign _0237_ = _1108_[0] ? rb[27] : rb[26];
  assign _0238_ = _1108_[0] ? rb[31] : rb[30];
  assign _0239_ = _1108_[0] ? rb[35] : rb[34];
  assign _0240_ = _1108_[0] ? rb[39] : rb[38];
  assign _0241_ = _1108_[0] ? rb[43] : rb[42];
  assign _0242_ = _1108_[0] ? rb[47] : rb[46];
  assign _0243_ = _1108_[0] ? rb[51] : rb[50];
  assign _0244_ = _1108_[0] ? rb[55] : rb[54];
  assign _0245_ = _1108_[0] ? rb[59] : rb[58];
  assign _0246_ = _1108_[0] ? rb[63] : rb[62];
  assign _0247_ = _1108_[2] ? _0987_ : _0986_;
  assign _0248_ = _1108_[2] ? _0991_ : _0990_;
  assign _0249_ = _1108_[2] ? _0995_ : _0994_;
  assign _0250_ = _1108_[2] ? _0999_ : _0998_;
  assign _0251_ = _1108_[4] ? _1003_ : _1002_;
  assign _0252_ = _1111_[0] ? rb[3] : rb[2];
  assign _0253_ = _1111_[0] ? rb[7] : rb[6];
  assign _0254_ = _1111_[0] ? rb[11] : rb[10];
  assign _0255_ = _1111_[0] ? rb[15] : rb[14];
  assign _0256_ = _1111_[0] ? rb[19] : rb[18];
  assign _0257_ = _1111_[0] ? rb[23] : rb[22];
  assign _0258_ = _1111_[0] ? rb[27] : rb[26];
  assign _0259_ = _1111_[0] ? rb[31] : rb[30];
  assign _0260_ = _1111_[0] ? rb[35] : rb[34];
  assign _0261_ = _1111_[0] ? rb[39] : rb[38];
  assign _0262_ = _1111_[0] ? rb[43] : rb[42];
  assign _0263_ = _1111_[0] ? rb[47] : rb[46];
  assign _0264_ = _1111_[0] ? rb[51] : rb[50];
  assign _0265_ = _1111_[0] ? rb[55] : rb[54];
  assign _0266_ = _1111_[0] ? rb[59] : rb[58];
  assign _0267_ = _1111_[0] ? rb[63] : rb[62];
  assign _0268_ = _1111_[2] ? _1008_ : _1007_;
  assign _0269_ = _1111_[2] ? _1012_ : _1011_;
  assign _0270_ = _1111_[2] ? _1016_ : _1015_;
  assign _0271_ = _1111_[2] ? _1020_ : _1019_;
  assign _0272_ = _1111_[4] ? _1024_ : _1023_;
  assign _0273_ = _1114_[0] ? rb[3] : rb[2];
  assign _0274_ = _1114_[0] ? rb[7] : rb[6];
  assign _0275_ = _1114_[0] ? rb[11] : rb[10];
  assign _0276_ = _1114_[0] ? rb[15] : rb[14];
  assign _0277_ = _1114_[0] ? rb[19] : rb[18];
  assign _0278_ = _1114_[0] ? rb[23] : rb[22];
  assign _0279_ = _1114_[0] ? rb[27] : rb[26];
  assign _0280_ = _1114_[0] ? rb[31] : rb[30];
  assign _0281_ = _1114_[0] ? rb[35] : rb[34];
  assign _0282_ = _1114_[0] ? rb[39] : rb[38];
  assign _0283_ = _1114_[0] ? rb[43] : rb[42];
  assign _0284_ = _1114_[0] ? rb[47] : rb[46];
  assign _0285_ = _1114_[0] ? rb[51] : rb[50];
  assign _0286_ = _1114_[0] ? rb[55] : rb[54];
  assign _0287_ = _1114_[0] ? rb[59] : rb[58];
  assign _0288_ = _1114_[0] ? rb[63] : rb[62];
  assign _0289_ = _1114_[2] ? _1029_ : _1028_;
  assign _0290_ = _1114_[2] ? _1033_ : _1032_;
  assign _0291_ = _1114_[2] ? _1037_ : _1036_;
  assign _0292_ = _1114_[2] ? _1041_ : _1040_;
  assign _0293_ = _1114_[4] ? _1045_ : _1044_;
  assign _0294_ = _1117_[0] ? rb[3] : rb[2];
  assign _0295_ = _1117_[0] ? rb[7] : rb[6];
  assign _0296_ = _1117_[0] ? rb[11] : rb[10];
  assign _0297_ = _1117_[0] ? rb[15] : rb[14];
  assign _0298_ = _1117_[0] ? rb[19] : rb[18];
  assign _0299_ = _1117_[0] ? rb[23] : rb[22];
  assign _0300_ = _1117_[0] ? rb[27] : rb[26];
  assign _0301_ = _1117_[0] ? rb[31] : rb[30];
  assign _0302_ = _1117_[0] ? rb[35] : rb[34];
  assign _0303_ = _1117_[0] ? rb[39] : rb[38];
  assign _0304_ = _1117_[0] ? rb[43] : rb[42];
  assign _0305_ = _1117_[0] ? rb[47] : rb[46];
  assign _0306_ = _1117_[0] ? rb[51] : rb[50];
  assign _0307_ = _1117_[0] ? rb[55] : rb[54];
  assign _0308_ = _1117_[0] ? rb[59] : rb[58];
  assign _0309_ = _1117_[0] ? rb[63] : rb[62];
  assign _0310_ = _1117_[2] ? _1050_ : _1049_;
  assign _0311_ = _1117_[2] ? _1054_ : _1053_;
  assign _0312_ = _1117_[2] ? _1058_ : _1057_;
  assign _0313_ = _1117_[2] ? _1062_ : _1061_;
  assign _0314_ = _1117_[4] ? _1066_ : _1065_;
  assign _0315_ = _1120_[0] ? rb[3] : rb[2];
  assign _0316_ = _1120_[0] ? rb[7] : rb[6];
  assign _0317_ = _1120_[0] ? rb[11] : rb[10];
  assign _0318_ = _1120_[0] ? rb[15] : rb[14];
  assign _0319_ = _1120_[0] ? rb[19] : rb[18];
  assign _0320_ = _1120_[0] ? rb[23] : rb[22];
  assign _0321_ = _1120_[0] ? rb[27] : rb[26];
  assign _0322_ = _1120_[0] ? rb[31] : rb[30];
  assign _0323_ = _1120_[0] ? rb[35] : rb[34];
  assign _0324_ = _1120_[0] ? rb[39] : rb[38];
  assign _0325_ = _1120_[0] ? rb[43] : rb[42];
  assign _0326_ = _1120_[0] ? rb[47] : rb[46];
  assign _0327_ = _1120_[0] ? rb[51] : rb[50];
  assign _0328_ = _1120_[0] ? rb[55] : rb[54];
  assign _0329_ = _1120_[0] ? rb[59] : rb[58];
  assign _0330_ = _1120_[0] ? rb[63] : rb[62];
  assign _0331_ = _1120_[2] ? _1071_ : _1070_;
  assign _0332_ = _1120_[2] ? _1075_ : _1074_;
  assign _0333_ = _1120_[2] ? _1079_ : _1078_;
  assign _0334_ = _1120_[2] ? _1083_ : _1082_;
  assign _0335_ = _1120_[4] ? _1087_ : _1086_;
  assign _0921_ = _1099_[1] ? _0168_ : _0000_;
  assign _0922_ = _1099_[1] ? _0169_ : _0001_;
  assign _0923_ = _1099_[1] ? _0170_ : _0002_;
  assign _0924_ = _1099_[1] ? _0171_ : _0003_;
  assign _0925_ = _1099_[1] ? _0172_ : _0004_;
  assign _0926_ = _1099_[1] ? _0173_ : _0005_;
  assign _0927_ = _1099_[1] ? _0174_ : _0006_;
  assign _0928_ = _1099_[1] ? _0175_ : _0007_;
  assign _0929_ = _1099_[1] ? _0176_ : _0008_;
  assign _0930_ = _1099_[1] ? _0177_ : _0009_;
  assign _0931_ = _1099_[1] ? _0178_ : _0010_;
  assign _0932_ = _1099_[1] ? _0179_ : _0011_;
  assign _0933_ = _1099_[1] ? _0180_ : _0012_;
  assign _0934_ = _1099_[1] ? _0181_ : _0013_;
  assign _0935_ = _1099_[1] ? _0182_ : _0014_;
  assign _0936_ = _1099_[1] ? _0183_ : _0015_;
  assign _0937_ = _1099_[3] ? _0184_ : _0016_;
  assign _0938_ = _1099_[3] ? _0185_ : _0017_;
  assign _0939_ = _1099_[3] ? _0186_ : _0018_;
  assign _0940_ = _1099_[3] ? _0187_ : _0019_;
  assign _0941_ = _1099_[5] ? _0188_ : _0020_;
  assign _0942_ = _1102_[1] ? _0189_ : _0021_;
  assign _0943_ = _1102_[1] ? _0190_ : _0022_;
  assign _0944_ = _1102_[1] ? _0191_ : _0023_;
  assign _0945_ = _1102_[1] ? _0192_ : _0024_;
  assign _0946_ = _1102_[1] ? _0193_ : _0025_;
  assign _0947_ = _1102_[1] ? _0194_ : _0026_;
  assign _0948_ = _1102_[1] ? _0195_ : _0027_;
  assign _0949_ = _1102_[1] ? _0196_ : _0028_;
  assign _0950_ = _1102_[1] ? _0197_ : _0029_;
  assign _0951_ = _1102_[1] ? _0198_ : _0030_;
  assign _0952_ = _1102_[1] ? _0199_ : _0031_;
  assign _0953_ = _1102_[1] ? _0200_ : _0032_;
  assign _0954_ = _1102_[1] ? _0201_ : _0033_;
  assign _0955_ = _1102_[1] ? _0202_ : _0034_;
  assign _0956_ = _1102_[1] ? _0203_ : _0035_;
  assign _0957_ = _1102_[1] ? _0204_ : _0036_;
  assign _0958_ = _1102_[3] ? _0205_ : _0037_;
  assign _0959_ = _1102_[3] ? _0206_ : _0038_;
  assign _0960_ = _1102_[3] ? _0207_ : _0039_;
  assign _0961_ = _1102_[3] ? _0208_ : _0040_;
  assign _0962_ = _1102_[5] ? _0209_ : _0041_;
  assign _0963_ = _1105_[1] ? _0210_ : _0042_;
  assign _0964_ = _1105_[1] ? _0211_ : _0043_;
  assign _0965_ = _1105_[1] ? _0212_ : _0044_;
  assign _0966_ = _1105_[1] ? _0213_ : _0045_;
  assign _0967_ = _1105_[1] ? _0214_ : _0046_;
  assign _0968_ = _1105_[1] ? _0215_ : _0047_;
  assign _0969_ = _1105_[1] ? _0216_ : _0048_;
  assign _0970_ = _1105_[1] ? _0217_ : _0049_;
  assign _0971_ = _1105_[1] ? _0218_ : _0050_;
  assign _0972_ = _1105_[1] ? _0219_ : _0051_;
  assign _0973_ = _1105_[1] ? _0220_ : _0052_;
  assign _0974_ = _1105_[1] ? _0221_ : _0053_;
  assign _0975_ = _1105_[1] ? _0222_ : _0054_;
  assign _0976_ = _1105_[1] ? _0223_ : _0055_;
  assign _0977_ = _1105_[1] ? _0224_ : _0056_;
  assign _0978_ = _1105_[1] ? _0225_ : _0057_;
  assign _0979_ = _1105_[3] ? _0226_ : _0058_;
  assign _0980_ = _1105_[3] ? _0227_ : _0059_;
  assign _0981_ = _1105_[3] ? _0228_ : _0060_;
  assign _0982_ = _1105_[3] ? _0229_ : _0061_;
  assign _0983_ = _1105_[5] ? _0230_ : _0062_;
  assign _0984_ = _1108_[1] ? _0231_ : _0063_;
  assign _0985_ = _1108_[1] ? _0232_ : _0064_;
  assign _0986_ = _1108_[1] ? _0233_ : _0065_;
  assign _0987_ = _1108_[1] ? _0234_ : _0066_;
  assign _0988_ = _1108_[1] ? _0235_ : _0067_;
  assign _0989_ = _1108_[1] ? _0236_ : _0068_;
  assign _0990_ = _1108_[1] ? _0237_ : _0069_;
  assign _0991_ = _1108_[1] ? _0238_ : _0070_;
  assign _0992_ = _1108_[1] ? _0239_ : _0071_;
  assign _0993_ = _1108_[1] ? _0240_ : _0072_;
  assign _0994_ = _1108_[1] ? _0241_ : _0073_;
  assign _0995_ = _1108_[1] ? _0242_ : _0074_;
  assign _0996_ = _1108_[1] ? _0243_ : _0075_;
  assign _0997_ = _1108_[1] ? _0244_ : _0076_;
  assign _0998_ = _1108_[1] ? _0245_ : _0077_;
  assign _0999_ = _1108_[1] ? _0246_ : _0078_;
  assign _1000_ = _1108_[3] ? _0247_ : _0079_;
  assign _1001_ = _1108_[3] ? _0248_ : _0080_;
  assign _1002_ = _1108_[3] ? _0249_ : _0081_;
  assign _1003_ = _1108_[3] ? _0250_ : _0082_;
  assign _1004_ = _1108_[5] ? _0251_ : _0083_;
  assign _1005_ = _1111_[1] ? _0252_ : _0084_;
  assign _1006_ = _1111_[1] ? _0253_ : _0085_;
  assign _1007_ = _1111_[1] ? _0254_ : _0086_;
  assign _1008_ = _1111_[1] ? _0255_ : _0087_;
  assign _1009_ = _1111_[1] ? _0256_ : _0088_;
  assign _1010_ = _1111_[1] ? _0257_ : _0089_;
  assign _1011_ = _1111_[1] ? _0258_ : _0090_;
  assign _1012_ = _1111_[1] ? _0259_ : _0091_;
  assign _1013_ = _1111_[1] ? _0260_ : _0092_;
  assign _1014_ = _1111_[1] ? _0261_ : _0093_;
  assign _1015_ = _1111_[1] ? _0262_ : _0094_;
  assign _1016_ = _1111_[1] ? _0263_ : _0095_;
  assign _1017_ = _1111_[1] ? _0264_ : _0096_;
  assign _1018_ = _1111_[1] ? _0265_ : _0097_;
  assign _1019_ = _1111_[1] ? _0266_ : _0098_;
  assign _1020_ = _1111_[1] ? _0267_ : _0099_;
  assign _1021_ = _1111_[3] ? _0268_ : _0100_;
  assign _1022_ = _1111_[3] ? _0269_ : _0101_;
  assign _1023_ = _1111_[3] ? _0270_ : _0102_;
  assign _1024_ = _1111_[3] ? _0271_ : _0103_;
  assign _1025_ = _1111_[5] ? _0272_ : _0104_;
  assign _1026_ = _1114_[1] ? _0273_ : _0105_;
  assign _1027_ = _1114_[1] ? _0274_ : _0106_;
  assign _1028_ = _1114_[1] ? _0275_ : _0107_;
  assign _1029_ = _1114_[1] ? _0276_ : _0108_;
  assign _1030_ = _1114_[1] ? _0277_ : _0109_;
  assign _1031_ = _1114_[1] ? _0278_ : _0110_;
  assign _1032_ = _1114_[1] ? _0279_ : _0111_;
  assign _1033_ = _1114_[1] ? _0280_ : _0112_;
  assign _1034_ = _1114_[1] ? _0281_ : _0113_;
  assign _1035_ = _1114_[1] ? _0282_ : _0114_;
  assign _1036_ = _1114_[1] ? _0283_ : _0115_;
  assign _1037_ = _1114_[1] ? _0284_ : _0116_;
  assign _1038_ = _1114_[1] ? _0285_ : _0117_;
  assign _1039_ = _1114_[1] ? _0286_ : _0118_;
  assign _1040_ = _1114_[1] ? _0287_ : _0119_;
  assign _1041_ = _1114_[1] ? _0288_ : _0120_;
  assign _1042_ = _1114_[3] ? _0289_ : _0121_;
  assign _1043_ = _1114_[3] ? _0290_ : _0122_;
  assign _1044_ = _1114_[3] ? _0291_ : _0123_;
  assign _1045_ = _1114_[3] ? _0292_ : _0124_;
  assign _1046_ = _1114_[5] ? _0293_ : _0125_;
  assign _1047_ = _1117_[1] ? _0294_ : _0126_;
  assign _1048_ = _1117_[1] ? _0295_ : _0127_;
  assign _1049_ = _1117_[1] ? _0296_ : _0128_;
  assign _1050_ = _1117_[1] ? _0297_ : _0129_;
  assign _1051_ = _1117_[1] ? _0298_ : _0130_;
  assign _1052_ = _1117_[1] ? _0299_ : _0131_;
  assign _1053_ = _1117_[1] ? _0300_ : _0132_;
  assign _1054_ = _1117_[1] ? _0301_ : _0133_;
  assign _1055_ = _1117_[1] ? _0302_ : _0134_;
  assign _1056_ = _1117_[1] ? _0303_ : _0135_;
  assign _1057_ = _1117_[1] ? _0304_ : _0136_;
  assign _1058_ = _1117_[1] ? _0305_ : _0137_;
  assign _1059_ = _1117_[1] ? _0306_ : _0138_;
  assign _1060_ = _1117_[1] ? _0307_ : _0139_;
  assign _1061_ = _1117_[1] ? _0308_ : _0140_;
  assign _1062_ = _1117_[1] ? _0309_ : _0141_;
  assign _1063_ = _1117_[3] ? _0310_ : _0142_;
  assign _1064_ = _1117_[3] ? _0311_ : _0143_;
  assign _1065_ = _1117_[3] ? _0312_ : _0144_;
  assign _1066_ = _1117_[3] ? _0313_ : _0145_;
  assign _1067_ = _1117_[5] ? _0314_ : _0146_;
  assign _1068_ = _1120_[1] ? _0315_ : _0147_;
  assign _1069_ = _1120_[1] ? _0316_ : _0148_;
  assign _1070_ = _1120_[1] ? _0317_ : _0149_;
  assign _1071_ = _1120_[1] ? _0318_ : _0150_;
  assign _1072_ = _1120_[1] ? _0319_ : _0151_;
  assign _1073_ = _1120_[1] ? _0320_ : _0152_;
  assign _1074_ = _1120_[1] ? _0321_ : _0153_;
  assign _1075_ = _1120_[1] ? _0322_ : _0154_;
  assign _1076_ = _1120_[1] ? _0323_ : _0155_;
  assign _1077_ = _1120_[1] ? _0324_ : _0156_;
  assign _1078_ = _1120_[1] ? _0325_ : _0157_;
  assign _1079_ = _1120_[1] ? _0326_ : _0158_;
  assign _1080_ = _1120_[1] ? _0327_ : _0159_;
  assign _1081_ = _1120_[1] ? _0328_ : _0160_;
  assign _1082_ = _1120_[1] ? _0329_ : _0161_;
  assign _1083_ = _1120_[1] ? _0330_ : _0162_;
  assign _1084_ = _1120_[3] ? _0331_ : _0163_;
  assign _1085_ = _1120_[3] ? _0332_ : _0164_;
  assign _1086_ = _1120_[3] ? _0333_ : _0165_;
  assign _1087_ = _1120_[3] ? _0334_ : _0166_;
  assign _1088_ = _1120_[5] ? _0335_ : _0167_;
  assign _1089_ = rs[0] ^ rs[8];
  assign _1090_ = _1089_ ^ rs[16];
  assign _1091_ = _1090_ ^ rs[24];
  assign _1092_ = rs[32] ^ rs[40];
  assign _1093_ = _1092_ ^ rs[48];
  assign _1094_ = _1093_ ^ rs[56];
  assign _1095_ = par0 ^ par1;
  assign _1096_ = datalen[3] ? _1095_ : par0;
  assign _1097_ = datalen[3] ? 1'h0 : par1;
  assign _1098_ = rs[7:6] == 2'h0;
  assign _1099_ = ~ rs[5:0];
  assign _1100_ = _1098_ ? _0941_ : 1'h0;
  assign _1101_ = rs[15:14] == 2'h0;
  assign _1102_ = ~ rs[13:8];
  assign _1103_ = _1101_ ? _0962_ : 1'h0;
  assign _1104_ = rs[23:22] == 2'h0;
  assign _1105_ = ~ rs[21:16];
  assign _1106_ = _1104_ ? _0983_ : 1'h0;
  assign _1107_ = rs[31:30] == 2'h0;
  assign _1108_ = ~ rs[29:24];
  assign _1109_ = _1107_ ? _1004_ : 1'h0;
  assign _1110_ = rs[39:38] == 2'h0;
  assign _1111_ = ~ rs[37:32];
  assign _1112_ = _1110_ ? _1025_ : 1'h0;
  assign _1113_ = rs[47:46] == 2'h0;
  assign _1114_ = ~ rs[45:40];
  assign _1115_ = _1113_ ? _1046_ : 1'h0;
  assign _1116_ = rs[55:54] == 2'h0;
  assign _1117_ = ~ rs[53:48];
  assign _1118_ = _1116_ ? _1067_ : 1'h0;
  assign _1119_ = rs[63:62] == 2'h0;
  assign _1120_ = ~ rs[61:56];
  assign _1121_ = _1119_ ? _1088_ : 1'h0;
  assign _1122_ = ~ rb;
  assign _1123_ = invert_in ? _1122_ : rb;
  assign _1124_ = rs & _1123_;
  assign _1125_ = op == 6'h03;
  assign _1126_ = rs | _1123_;
  assign _1127_ = op == 6'h2c;
  assign _1128_ = rs ^ _1123_;
  function [63:0] \29091 ;
    input [63:0] a;
    input [127:0] b;
    input [1:0] s;
    (* parallel_case *)
    casez (s)
      2'b?1:
        \29091  = b[63:0];
      2'b1?:
        \29091  = b[127:64];
      default:
        \29091  = a;
    endcase
  endfunction
  assign _1129_ = \29091 (_1128_, { _1126_, _1124_ }, { _1127_, _1125_ });
  assign _1130_ = ~ _1129_;
  assign _1131_ = invert_out ? _1130_ : _1129_;
  assign _1132_ = op == 6'h03;
  assign _1133_ = op == 6'h2c;
  assign _1134_ = _1132_ | _1133_;
  assign _1135_ = op == 6'h3a;
  assign _1136_ = _1134_ | _1135_;
  assign _1137_ = op == 6'h2e;
  assign _1138_ = rs[7:0] == rb[7:0];
  assign _1139_ = _1138_ ? 8'hff : 8'h00;
  assign _1140_ = rs[15:8] == rb[15:8];
  assign _1141_ = _1140_ ? 8'hff : 8'h00;
  assign _1142_ = rs[23:16] == rb[23:16];
  assign _1143_ = _1142_ ? 8'hff : 8'h00;
  assign _1144_ = rs[31:24] == rb[31:24];
  assign _1145_ = _1144_ ? 8'hff : 8'h00;
  assign _1146_ = rs[39:32] == rb[39:32];
  assign _1147_ = _1146_ ? 8'hff : 8'h00;
  assign _1148_ = rs[47:40] == rb[47:40];
  assign _1149_ = _1148_ ? 8'hff : 8'h00;
  assign _1150_ = rs[55:48] == rb[55:48];
  assign _1151_ = _1150_ ? 8'hff : 8'h00;
  assign _1152_ = rs[63:56] == rb[63:56];
  assign _1153_ = _1152_ ? 8'hff : 8'h00;
  assign _1154_ = op == 6'h0a;
  assign _1155_ = op == 6'h08;
  assign _1156_ = ~ invert_in;
  assign _1157_ = rs[50] & rs[55];
  assign _1158_ = _1157_ & rs[47];
  assign _1159_ = ~ rs[51];
  assign _1160_ = _1158_ & _1159_;
  assign _1161_ = rs[46] & rs[55];
  assign _1162_ = ~ rs[47];
  assign _1163_ = _1161_ & _1162_;
  assign _1164_ = _1160_ | _1163_;
  assign _1165_ = ~ rs[55];
  assign _1166_ = rs[54] & _1165_;
  assign _1167_ = _1164_ | _1166_;
  assign _1168_ = rs[49] & rs[55];
  assign _1169_ = _1168_ & rs[47];
  assign _1170_ = ~ rs[51];
  assign _1171_ = _1169_ & _1170_;
  assign _1172_ = rs[45] & rs[55];
  assign _1173_ = ~ rs[47];
  assign _1174_ = _1172_ & _1173_;
  assign _1175_ = _1171_ | _1174_;
  assign _1176_ = ~ rs[55];
  assign _1177_ = rs[53] & _1176_;
  assign _1178_ = _1175_ | _1177_;
  assign _1179_ = ~ rs[55];
  assign _1180_ = rs[46] & _1179_;
  assign _1181_ = _1180_ & rs[51];
  assign _1182_ = ~ rs[47];
  assign _1183_ = _1181_ & _1182_;
  assign _1184_ = ~ rs[47];
  assign _1185_ = rs[50] & _1184_;
  assign _1186_ = ~ rs[51];
  assign _1187_ = _1185_ & _1186_;
  assign _1188_ = _1183_ | _1187_;
  assign _1189_ = ~ rs[55];
  assign _1190_ = rs[50] & _1189_;
  assign _1191_ = ~ rs[51];
  assign _1192_ = _1190_ & _1191_;
  assign _1193_ = _1188_ | _1192_;
  assign _1194_ = rs[51] & rs[47];
  assign _1195_ = _1193_ | _1194_;
  assign _1196_ = ~ rs[55];
  assign _1197_ = rs[45] & _1196_;
  assign _1198_ = _1197_ & rs[51];
  assign _1199_ = ~ rs[47];
  assign _1200_ = _1198_ & _1199_;
  assign _1201_ = ~ rs[47];
  assign _1202_ = rs[49] & _1201_;
  assign _1203_ = ~ rs[51];
  assign _1204_ = _1202_ & _1203_;
  assign _1205_ = _1200_ | _1204_;
  assign _1206_ = ~ rs[55];
  assign _1207_ = rs[49] & _1206_;
  assign _1208_ = ~ rs[51];
  assign _1209_ = _1207_ & _1208_;
  assign _1210_ = _1205_ | _1209_;
  assign _1211_ = rs[55] & rs[47];
  assign _1212_ = _1210_ | _1211_;
  assign _1213_ = rs[55] | rs[51];
  assign _1214_ = _1213_ | rs[47];
  assign _1215_ = ~ rs[51];
  assign _1216_ = _1215_ & rs[46];
  assign _1217_ = ~ rs[47];
  assign _1218_ = _1216_ & _1217_;
  assign _1219_ = rs[51] & rs[47];
  assign _1220_ = _1218_ | _1219_;
  assign _1221_ = _1220_ | rs[55];
  assign _1222_ = ~ rs[55];
  assign _1223_ = _1222_ & rs[45];
  assign _1224_ = ~ rs[47];
  assign _1225_ = _1223_ & _1224_;
  assign _1226_ = rs[55] & rs[47];
  assign _1227_ = _1225_ | _1226_;
  assign _1228_ = _1227_ | rs[51];
  assign _1229_ = rs[38] & rs[43];
  assign _1230_ = _1229_ & rs[35];
  assign _1231_ = ~ rs[39];
  assign _1232_ = _1230_ & _1231_;
  assign _1233_ = rs[34] & rs[43];
  assign _1234_ = ~ rs[35];
  assign _1235_ = _1233_ & _1234_;
  assign _1236_ = _1232_ | _1235_;
  assign _1237_ = ~ rs[43];
  assign _1238_ = rs[42] & _1237_;
  assign _1239_ = _1236_ | _1238_;
  assign _1240_ = rs[37] & rs[43];
  assign _1241_ = _1240_ & rs[35];
  assign _1242_ = ~ rs[39];
  assign _1243_ = _1241_ & _1242_;
  assign _1244_ = rs[33] & rs[43];
  assign _1245_ = ~ rs[35];
  assign _1246_ = _1244_ & _1245_;
  assign _1247_ = _1243_ | _1246_;
  assign _1248_ = ~ rs[43];
  assign _1249_ = rs[41] & _1248_;
  assign _1250_ = _1247_ | _1249_;
  assign _1251_ = ~ rs[43];
  assign _1252_ = rs[34] & _1251_;
  assign _1253_ = _1252_ & rs[39];
  assign _1254_ = ~ rs[35];
  assign _1255_ = _1253_ & _1254_;
  assign _1256_ = ~ rs[35];
  assign _1257_ = rs[38] & _1256_;
  assign _1258_ = ~ rs[39];
  assign _1259_ = _1257_ & _1258_;
  assign _1260_ = _1255_ | _1259_;
  assign _1261_ = ~ rs[43];
  assign _1262_ = rs[38] & _1261_;
  assign _1263_ = ~ rs[39];
  assign _1264_ = _1262_ & _1263_;
  assign _1265_ = _1260_ | _1264_;
  assign _1266_ = rs[39] & rs[35];
  assign _1267_ = _1265_ | _1266_;
  assign _1268_ = ~ rs[43];
  assign _1269_ = rs[33] & _1268_;
  assign _1270_ = _1269_ & rs[39];
  assign _1271_ = ~ rs[35];
  assign _1272_ = _1270_ & _1271_;
  assign _1273_ = ~ rs[35];
  assign _1274_ = rs[37] & _1273_;
  assign _1275_ = ~ rs[39];
  assign _1276_ = _1274_ & _1275_;
  assign _1277_ = _1272_ | _1276_;
  assign _1278_ = ~ rs[43];
  assign _1279_ = rs[37] & _1278_;
  assign _1280_ = ~ rs[39];
  assign _1281_ = _1279_ & _1280_;
  assign _1282_ = _1277_ | _1281_;
  assign _1283_ = rs[43] & rs[35];
  assign _1284_ = _1282_ | _1283_;
  assign _1285_ = rs[43] | rs[39];
  assign _1286_ = _1285_ | rs[35];
  assign _1287_ = ~ rs[39];
  assign _1288_ = _1287_ & rs[34];
  assign _1289_ = ~ rs[35];
  assign _1290_ = _1288_ & _1289_;
  assign _1291_ = rs[39] & rs[35];
  assign _1292_ = _1290_ | _1291_;
  assign _1293_ = _1292_ | rs[43];
  assign _1294_ = ~ rs[43];
  assign _1295_ = _1294_ & rs[33];
  assign _1296_ = ~ rs[35];
  assign _1297_ = _1295_ & _1296_;
  assign _1298_ = rs[43] & rs[35];
  assign _1299_ = _1297_ | _1298_;
  assign _1300_ = _1299_ | rs[39];
  assign _1301_ = rs[18] & rs[23];
  assign _1302_ = _1301_ & rs[15];
  assign _1303_ = ~ rs[19];
  assign _1304_ = _1302_ & _1303_;
  assign _1305_ = rs[14] & rs[23];
  assign _1306_ = ~ rs[15];
  assign _1307_ = _1305_ & _1306_;
  assign _1308_ = _1304_ | _1307_;
  assign _1309_ = ~ rs[23];
  assign _1310_ = rs[22] & _1309_;
  assign _1311_ = _1308_ | _1310_;
  assign _1312_ = rs[17] & rs[23];
  assign _1313_ = _1312_ & rs[15];
  assign _1314_ = ~ rs[19];
  assign _1315_ = _1313_ & _1314_;
  assign _1316_ = rs[13] & rs[23];
  assign _1317_ = ~ rs[15];
  assign _1318_ = _1316_ & _1317_;
  assign _1319_ = _1315_ | _1318_;
  assign _1320_ = ~ rs[23];
  assign _1321_ = rs[21] & _1320_;
  assign _1322_ = _1319_ | _1321_;
  assign _1323_ = ~ rs[23];
  assign _1324_ = rs[14] & _1323_;
  assign _1325_ = _1324_ & rs[19];
  assign _1326_ = ~ rs[15];
  assign _1327_ = _1325_ & _1326_;
  assign _1328_ = ~ rs[15];
  assign _1329_ = rs[18] & _1328_;
  assign _1330_ = ~ rs[19];
  assign _1331_ = _1329_ & _1330_;
  assign _1332_ = _1327_ | _1331_;
  assign _1333_ = ~ rs[23];
  assign _1334_ = rs[18] & _1333_;
  assign _1335_ = ~ rs[19];
  assign _1336_ = _1334_ & _1335_;
  assign _1337_ = _1332_ | _1336_;
  assign _1338_ = rs[19] & rs[15];
  assign _1339_ = _1337_ | _1338_;
  assign _1340_ = ~ rs[23];
  assign _1341_ = rs[13] & _1340_;
  assign _1342_ = _1341_ & rs[19];
  assign _1343_ = ~ rs[15];
  assign _1344_ = _1342_ & _1343_;
  assign _1345_ = ~ rs[15];
  assign _1346_ = rs[17] & _1345_;
  assign _1347_ = ~ rs[19];
  assign _1348_ = _1346_ & _1347_;
  assign _1349_ = _1344_ | _1348_;
  assign _1350_ = ~ rs[23];
  assign _0336_ = rs[17] & _1350_;
  assign _0337_ = ~ rs[19];
  assign _0338_ = _0336_ & _0337_;
  assign _0339_ = _1349_ | _0338_;
  assign _0340_ = rs[23] & rs[15];
  assign _0341_ = _0339_ | _0340_;
  assign _0342_ = rs[23] | rs[19];
  assign _0343_ = _0342_ | rs[15];
  assign _0344_ = ~ rs[19];
  assign _0345_ = _0344_ & rs[14];
  assign _0346_ = ~ rs[15];
  assign _0347_ = _0345_ & _0346_;
  assign _0348_ = rs[19] & rs[15];
  assign _0349_ = _0347_ | _0348_;
  assign _0350_ = _0349_ | rs[23];
  assign _0351_ = ~ rs[23];
  assign _0352_ = _0351_ & rs[13];
  assign _0353_ = ~ rs[15];
  assign _0354_ = _0352_ & _0353_;
  assign _0355_ = rs[23] & rs[15];
  assign _0356_ = _0354_ | _0355_;
  assign _0357_ = _0356_ | rs[19];
  assign _0358_ = rs[6] & rs[11];
  assign _0359_ = _0358_ & rs[3];
  assign _0360_ = ~ rs[7];
  assign _0361_ = _0359_ & _0360_;
  assign _0362_ = rs[2] & rs[11];
  assign _0363_ = ~ rs[3];
  assign _0364_ = _0362_ & _0363_;
  assign _0365_ = _0361_ | _0364_;
  assign _0366_ = ~ rs[11];
  assign _0367_ = rs[10] & _0366_;
  assign _0368_ = _0365_ | _0367_;
  assign _0369_ = rs[5] & rs[11];
  assign _0370_ = _0369_ & rs[3];
  assign _0371_ = ~ rs[7];
  assign _0372_ = _0370_ & _0371_;
  assign _0373_ = rs[1] & rs[11];
  assign _0374_ = ~ rs[3];
  assign _0375_ = _0373_ & _0374_;
  assign _0376_ = _0372_ | _0375_;
  assign _0377_ = ~ rs[11];
  assign _0378_ = rs[9] & _0377_;
  assign _0379_ = _0376_ | _0378_;
  assign _0380_ = ~ rs[11];
  assign _0381_ = rs[2] & _0380_;
  assign _0382_ = _0381_ & rs[7];
  assign _0383_ = ~ rs[3];
  assign _0384_ = _0382_ & _0383_;
  assign _0385_ = ~ rs[3];
  assign _0386_ = rs[6] & _0385_;
  assign _0387_ = ~ rs[7];
  assign _0388_ = _0386_ & _0387_;
  assign _0389_ = _0384_ | _0388_;
  assign _0390_ = ~ rs[11];
  assign _0391_ = rs[6] & _0390_;
  assign _0392_ = ~ rs[7];
  assign _0393_ = _0391_ & _0392_;
  assign _0394_ = _0389_ | _0393_;
  assign _0395_ = rs[7] & rs[3];
  assign _0396_ = _0394_ | _0395_;
  assign _0397_ = ~ rs[11];
  assign _0398_ = rs[1] & _0397_;
  assign _0399_ = _0398_ & rs[7];
  assign _0400_ = ~ rs[3];
  assign _0401_ = _0399_ & _0400_;
  assign _0402_ = ~ rs[3];
  assign _0403_ = rs[5] & _0402_;
  assign _0404_ = ~ rs[7];
  assign _0405_ = _0403_ & _0404_;
  assign _0406_ = _0401_ | _0405_;
  assign _0407_ = ~ rs[11];
  assign _0408_ = rs[5] & _0407_;
  assign _0409_ = ~ rs[7];
  assign _0410_ = _0408_ & _0409_;
  assign _0411_ = _0406_ | _0410_;
  assign _0412_ = rs[11] & rs[3];
  assign _0413_ = _0411_ | _0412_;
  assign _0414_ = rs[11] | rs[7];
  assign _0415_ = _0414_ | rs[3];
  assign _0416_ = ~ rs[7];
  assign _0417_ = _0416_ & rs[2];
  assign _0418_ = ~ rs[3];
  assign _0419_ = _0417_ & _0418_;
  assign _0420_ = rs[7] & rs[3];
  assign _0421_ = _0419_ | _0420_;
  assign _0422_ = _0421_ | rs[11];
  assign _0423_ = ~ rs[11];
  assign _0424_ = _0423_ & rs[1];
  assign _0425_ = ~ rs[3];
  assign _0426_ = _0424_ & _0425_;
  assign _0427_ = rs[11] & rs[3];
  assign _0428_ = _0426_ | _0427_;
  assign _0429_ = _0428_ | rs[7];
  assign _0430_ = ~ rs[48];
  assign _0431_ = _0430_ & rs[45];
  assign _0432_ = _0431_ & rs[44];
  assign _0433_ = rs[47] & rs[45];
  assign _0434_ = _0433_ & rs[44];
  assign _0435_ = _0434_ & rs[48];
  assign _0436_ = _0432_ | _0435_;
  assign _0437_ = rs[45] & rs[44];
  assign _0438_ = ~ rs[43];
  assign _0439_ = _0437_ & _0438_;
  assign _0440_ = _0436_ | _0439_;
  assign _0441_ = rs[51] & rs[48];
  assign _0442_ = _0441_ & rs[43];
  assign _0443_ = ~ rs[47];
  assign _0444_ = _0442_ & _0443_;
  assign _0445_ = ~ rs[44];
  assign _0446_ = rs[51] & _0445_;
  assign _0447_ = _0444_ | _0446_;
  assign _0448_ = ~ rs[45];
  assign _0449_ = rs[51] & _0448_;
  assign _0450_ = _0447_ | _0449_;
  assign _0451_ = rs[50] & rs[48];
  assign _0452_ = _0451_ & rs[43];
  assign _0453_ = ~ rs[47];
  assign _0454_ = _0452_ & _0453_;
  assign _0455_ = ~ rs[44];
  assign _0456_ = rs[50] & _0455_;
  assign _0457_ = _0454_ | _0456_;
  assign _0458_ = ~ rs[45];
  assign _0459_ = rs[50] & _0458_;
  assign _0460_ = _0457_ | _0459_;
  assign _0461_ = ~ rs[44];
  assign _0462_ = rs[45] & _0461_;
  assign _0463_ = _0462_ & rs[43];
  assign _0464_ = rs[48] & rs[45];
  assign _0465_ = _0464_ & rs[44];
  assign _0466_ = _0465_ & rs[43];
  assign _0467_ = _0463_ | _0466_;
  assign _0468_ = ~ rs[47];
  assign _0469_ = _0468_ & rs[45];
  assign _0470_ = _0469_ & rs[44];
  assign _0471_ = _0470_ & rs[43];
  assign _0472_ = _0467_ | _0471_;
  assign _0473_ = rs[51] & rs[47];
  assign _0474_ = _0473_ & rs[45];
  assign _0475_ = _0474_ & rs[44];
  assign _0476_ = _0475_ & rs[43];
  assign _0477_ = ~ rs[48];
  assign _0478_ = _0476_ & _0477_;
  assign _0479_ = ~ rs[43];
  assign _0480_ = rs[48] & _0479_;
  assign _0481_ = _0480_ & rs[45];
  assign _0482_ = _0478_ | _0481_;
  assign _0483_ = ~ rs[45];
  assign _0484_ = rs[48] & _0483_;
  assign _0485_ = _0482_ | _0484_;
  assign _0486_ = rs[50] & rs[47];
  assign _0487_ = _0486_ & rs[44];
  assign _0488_ = _0487_ & rs[45];
  assign _0489_ = _0488_ & rs[43];
  assign _0490_ = ~ rs[48];
  assign _0491_ = _0489_ & _0490_;
  assign _0492_ = ~ rs[43];
  assign _0493_ = rs[47] & _0492_;
  assign _0494_ = _0493_ & rs[45];
  assign _0495_ = _0491_ | _0494_;
  assign _0496_ = ~ rs[45];
  assign _0497_ = rs[47] & _0496_;
  assign _0498_ = _0495_ | _0497_;
  assign _0499_ = rs[47] & rs[45];
  assign _0500_ = _0499_ & rs[44];
  assign _0501_ = _0500_ & rs[43];
  assign _0502_ = rs[48] & rs[45];
  assign _0503_ = _0502_ & rs[44];
  assign _0504_ = _0503_ & rs[43];
  assign _0505_ = _0501_ | _0504_;
  assign _0506_ = ~ rs[44];
  assign _0507_ = rs[45] & _0506_;
  assign _0508_ = ~ rs[43];
  assign _0509_ = _0507_ & _0508_;
  assign _0510_ = _0505_ | _0509_;
  assign _0511_ = ~ rs[48];
  assign _0512_ = rs[51] & _0511_;
  assign _0513_ = ~ rs[47];
  assign _0514_ = _0512_ & _0513_;
  assign _0515_ = _0514_ & rs[44];
  assign _0516_ = _0515_ & rs[45];
  assign _0517_ = rs[48] & rs[45];
  assign _0518_ = ~ rs[44];
  assign _0519_ = _0517_ & _0518_;
  assign _0520_ = _0519_ & rs[43];
  assign _0521_ = _0516_ | _0520_;
  assign _0522_ = rs[51] & rs[44];
  assign _0523_ = ~ rs[43];
  assign _0524_ = _0522_ & _0523_;
  assign _0525_ = _0524_ & rs[45];
  assign _0526_ = _0521_ | _0525_;
  assign _0527_ = ~ rs[45];
  assign _0528_ = rs[44] & _0527_;
  assign _0529_ = _0526_ | _0528_;
  assign _0530_ = ~ rs[48];
  assign _0531_ = rs[50] & _0530_;
  assign _0532_ = ~ rs[47];
  assign _0533_ = _0531_ & _0532_;
  assign _0534_ = _0533_ & rs[45];
  assign _0535_ = _0534_ & rs[44];
  assign _0536_ = rs[47] & rs[45];
  assign _0537_ = ~ rs[44];
  assign _0538_ = _0536_ & _0537_;
  assign _0539_ = _0538_ & rs[43];
  assign _0540_ = _0535_ | _0539_;
  assign _0541_ = rs[50] & rs[45];
  assign _0542_ = _0541_ & rs[44];
  assign _0543_ = ~ rs[43];
  assign _0544_ = _0542_ & _0543_;
  assign _0545_ = _0540_ | _0544_;
  assign _0546_ = ~ rs[45];
  assign _0547_ = rs[43] & _0546_;
  assign _0548_ = _0545_ | _0547_;
  assign _0549_ = ~ rs[38];
  assign _0550_ = _0549_ & rs[35];
  assign _0551_ = _0550_ & rs[34];
  assign _0552_ = rs[37] & rs[35];
  assign _0553_ = _0552_ & rs[34];
  assign _0554_ = _0553_ & rs[38];
  assign _0555_ = _0551_ | _0554_;
  assign _0556_ = rs[35] & rs[34];
  assign _0557_ = ~ rs[33];
  assign _0558_ = _0556_ & _0557_;
  assign _0559_ = _0555_ | _0558_;
  assign _0560_ = rs[41] & rs[38];
  assign _0561_ = _0560_ & rs[33];
  assign _0562_ = ~ rs[37];
  assign _0563_ = _0561_ & _0562_;
  assign _0564_ = ~ rs[34];
  assign _0565_ = rs[41] & _0564_;
  assign _0566_ = _0563_ | _0565_;
  assign _0567_ = ~ rs[35];
  assign _0568_ = rs[41] & _0567_;
  assign _0569_ = _0566_ | _0568_;
  assign _0570_ = rs[40] & rs[38];
  assign _0571_ = _0570_ & rs[33];
  assign _0572_ = ~ rs[37];
  assign _0573_ = _0571_ & _0572_;
  assign _0574_ = ~ rs[34];
  assign _0575_ = rs[40] & _0574_;
  assign _0576_ = _0573_ | _0575_;
  assign _0577_ = ~ rs[35];
  assign _0578_ = rs[40] & _0577_;
  assign _0579_ = _0576_ | _0578_;
  assign _0580_ = ~ rs[34];
  assign _0581_ = rs[35] & _0580_;
  assign _0582_ = _0581_ & rs[33];
  assign _0583_ = rs[38] & rs[35];
  assign _0584_ = _0583_ & rs[34];
  assign _0585_ = _0584_ & rs[33];
  assign _0586_ = _0582_ | _0585_;
  assign _0587_ = ~ rs[37];
  assign _0588_ = _0587_ & rs[35];
  assign _0589_ = _0588_ & rs[34];
  assign _0590_ = _0589_ & rs[33];
  assign _0591_ = _0586_ | _0590_;
  assign _0592_ = rs[41] & rs[37];
  assign _0593_ = _0592_ & rs[35];
  assign _0594_ = _0593_ & rs[34];
  assign _0595_ = _0594_ & rs[33];
  assign _0596_ = ~ rs[38];
  assign _0597_ = _0595_ & _0596_;
  assign _0598_ = ~ rs[33];
  assign _0599_ = rs[38] & _0598_;
  assign _0600_ = _0599_ & rs[35];
  assign _0601_ = _0597_ | _0600_;
  assign _0602_ = ~ rs[35];
  assign _0603_ = rs[38] & _0602_;
  assign _0604_ = _0601_ | _0603_;
  assign _0605_ = rs[40] & rs[37];
  assign _0606_ = _0605_ & rs[34];
  assign _0607_ = _0606_ & rs[35];
  assign _0608_ = _0607_ & rs[33];
  assign _0609_ = ~ rs[38];
  assign _0610_ = _0608_ & _0609_;
  assign _0611_ = ~ rs[33];
  assign _0612_ = rs[37] & _0611_;
  assign _0613_ = _0612_ & rs[35];
  assign _0614_ = _0610_ | _0613_;
  assign _0615_ = ~ rs[35];
  assign _0616_ = rs[37] & _0615_;
  assign _0617_ = _0614_ | _0616_;
  assign _0618_ = rs[37] & rs[35];
  assign _0619_ = _0618_ & rs[34];
  assign _0620_ = _0619_ & rs[33];
  assign _0621_ = rs[38] & rs[35];
  assign _0622_ = _0621_ & rs[34];
  assign _0623_ = _0622_ & rs[33];
  assign _0624_ = _0620_ | _0623_;
  assign _0625_ = ~ rs[34];
  assign _0626_ = rs[35] & _0625_;
  assign _0627_ = ~ rs[33];
  assign _0628_ = _0626_ & _0627_;
  assign _0629_ = _0624_ | _0628_;
  assign _0630_ = ~ rs[38];
  assign _0631_ = rs[41] & _0630_;
  assign _0632_ = ~ rs[37];
  assign _0633_ = _0631_ & _0632_;
  assign _0634_ = _0633_ & rs[34];
  assign _0635_ = _0634_ & rs[35];
  assign _0636_ = rs[38] & rs[35];
  assign _0637_ = ~ rs[34];
  assign _0638_ = _0636_ & _0637_;
  assign _0639_ = _0638_ & rs[33];
  assign _0640_ = _0635_ | _0639_;
  assign _0641_ = rs[41] & rs[34];
  assign _0642_ = ~ rs[33];
  assign _0643_ = _0641_ & _0642_;
  assign _0644_ = _0643_ & rs[35];
  assign _0645_ = _0640_ | _0644_;
  assign _0646_ = ~ rs[35];
  assign _0647_ = rs[34] & _0646_;
  assign _0648_ = _0645_ | _0647_;
  assign _0649_ = ~ rs[38];
  assign _0650_ = rs[40] & _0649_;
  assign _0651_ = ~ rs[37];
  assign _0652_ = _0650_ & _0651_;
  assign _0653_ = _0652_ & rs[35];
  assign _0654_ = _0653_ & rs[34];
  assign _0655_ = rs[37] & rs[35];
  assign _0656_ = ~ rs[34];
  assign _0657_ = _0655_ & _0656_;
  assign _0658_ = _0657_ & rs[33];
  assign _0659_ = _0654_ | _0658_;
  assign _0660_ = rs[40] & rs[35];
  assign _0661_ = _0660_ & rs[34];
  assign _0662_ = ~ rs[33];
  assign _0663_ = _0661_ & _0662_;
  assign _0664_ = _0659_ | _0663_;
  assign _0665_ = ~ rs[35];
  assign _0666_ = rs[33] & _0665_;
  assign _0667_ = _0664_ | _0666_;
  assign _0668_ = ~ rs[16];
  assign _0669_ = _0668_ & rs[13];
  assign _0670_ = _0669_ & rs[12];
  assign _0671_ = rs[15] & rs[13];
  assign _0672_ = _0671_ & rs[12];
  assign _0673_ = _0672_ & rs[16];
  assign _0674_ = _0670_ | _0673_;
  assign _0675_ = rs[13] & rs[12];
  assign _0676_ = ~ rs[11];
  assign _0677_ = _0675_ & _0676_;
  assign _0678_ = _0674_ | _0677_;
  assign _0679_ = rs[19] & rs[16];
  assign _0680_ = _0679_ & rs[11];
  assign _0681_ = ~ rs[15];
  assign _0682_ = _0680_ & _0681_;
  assign _0683_ = ~ rs[12];
  assign _0684_ = rs[19] & _0683_;
  assign _0685_ = _0682_ | _0684_;
  assign _0686_ = ~ rs[13];
  assign _0687_ = rs[19] & _0686_;
  assign _0688_ = _0685_ | _0687_;
  assign _0689_ = rs[18] & rs[16];
  assign _0690_ = _0689_ & rs[11];
  assign _0691_ = ~ rs[15];
  assign _0692_ = _0690_ & _0691_;
  assign _0693_ = ~ rs[12];
  assign _0694_ = rs[18] & _0693_;
  assign _0695_ = _0692_ | _0694_;
  assign _0696_ = ~ rs[13];
  assign _0697_ = rs[18] & _0696_;
  assign _0698_ = _0695_ | _0697_;
  assign _0699_ = ~ rs[12];
  assign _0700_ = rs[13] & _0699_;
  assign _0701_ = _0700_ & rs[11];
  assign _0702_ = rs[16] & rs[13];
  assign _0703_ = _0702_ & rs[12];
  assign _0704_ = _0703_ & rs[11];
  assign _0705_ = _0701_ | _0704_;
  assign _0706_ = ~ rs[15];
  assign _0707_ = _0706_ & rs[13];
  assign _0708_ = _0707_ & rs[12];
  assign _0709_ = _0708_ & rs[11];
  assign _0710_ = _0705_ | _0709_;
  assign _0711_ = rs[19] & rs[15];
  assign _0712_ = _0711_ & rs[13];
  assign _0713_ = _0712_ & rs[12];
  assign _0714_ = _0713_ & rs[11];
  assign _0715_ = ~ rs[16];
  assign _0716_ = _0714_ & _0715_;
  assign _0717_ = ~ rs[11];
  assign _0718_ = rs[16] & _0717_;
  assign _0719_ = _0718_ & rs[13];
  assign _0720_ = _0716_ | _0719_;
  assign _0721_ = ~ rs[13];
  assign _0722_ = rs[16] & _0721_;
  assign _0723_ = _0720_ | _0722_;
  assign _0724_ = rs[18] & rs[15];
  assign _0725_ = _0724_ & rs[12];
  assign _0726_ = _0725_ & rs[13];
  assign _0727_ = _0726_ & rs[11];
  assign _0728_ = ~ rs[16];
  assign _0729_ = _0727_ & _0728_;
  assign _0730_ = ~ rs[11];
  assign _0731_ = rs[15] & _0730_;
  assign _0732_ = _0731_ & rs[13];
  assign _0733_ = _0729_ | _0732_;
  assign _0734_ = ~ rs[13];
  assign _0735_ = rs[15] & _0734_;
  assign _0736_ = _0733_ | _0735_;
  assign _0737_ = rs[15] & rs[13];
  assign _0738_ = _0737_ & rs[12];
  assign _0739_ = _0738_ & rs[11];
  assign _0740_ = rs[16] & rs[13];
  assign _0741_ = _0740_ & rs[12];
  assign _0742_ = _0741_ & rs[11];
  assign _0743_ = _0739_ | _0742_;
  assign _0744_ = ~ rs[12];
  assign _0745_ = rs[13] & _0744_;
  assign _0746_ = ~ rs[11];
  assign _0747_ = _0745_ & _0746_;
  assign _0748_ = _0743_ | _0747_;
  assign _0749_ = ~ rs[16];
  assign _0750_ = rs[19] & _0749_;
  assign _0751_ = ~ rs[15];
  assign _0752_ = _0750_ & _0751_;
  assign _0753_ = _0752_ & rs[12];
  assign _0754_ = _0753_ & rs[13];
  assign _0755_ = rs[16] & rs[13];
  assign _0756_ = ~ rs[12];
  assign _0757_ = _0755_ & _0756_;
  assign _0758_ = _0757_ & rs[11];
  assign _0759_ = _0754_ | _0758_;
  assign _0760_ = rs[19] & rs[12];
  assign _0761_ = ~ rs[11];
  assign _0762_ = _0760_ & _0761_;
  assign _0763_ = _0762_ & rs[13];
  assign _0764_ = _0759_ | _0763_;
  assign _0765_ = ~ rs[13];
  assign _0766_ = rs[12] & _0765_;
  assign _0767_ = _0764_ | _0766_;
  assign _0768_ = ~ rs[16];
  assign _0769_ = rs[18] & _0768_;
  assign _0770_ = ~ rs[15];
  assign _0771_ = _0769_ & _0770_;
  assign _0772_ = _0771_ & rs[13];
  assign _0773_ = _0772_ & rs[12];
  assign _0774_ = rs[15] & rs[13];
  assign _0775_ = ~ rs[12];
  assign _0776_ = _0774_ & _0775_;
  assign _0777_ = _0776_ & rs[11];
  assign _0778_ = _0773_ | _0777_;
  assign _0779_ = rs[18] & rs[13];
  assign _0780_ = _0779_ & rs[12];
  assign _0781_ = ~ rs[11];
  assign _0782_ = _0780_ & _0781_;
  assign _0783_ = _0778_ | _0782_;
  assign _0784_ = ~ rs[13];
  assign _0785_ = rs[11] & _0784_;
  assign _0786_ = _0783_ | _0785_;
  assign _0787_ = ~ rs[6];
  assign _0788_ = _0787_ & rs[3];
  assign _0789_ = _0788_ & rs[2];
  assign _0790_ = rs[5] & rs[3];
  assign _0791_ = _0790_ & rs[2];
  assign _0792_ = _0791_ & rs[6];
  assign _0793_ = _0789_ | _0792_;
  assign _0794_ = rs[3] & rs[2];
  assign _0795_ = ~ rs[1];
  assign _0796_ = _0794_ & _0795_;
  assign _0797_ = _0793_ | _0796_;
  assign _0798_ = rs[9] & rs[6];
  assign _0799_ = _0798_ & rs[1];
  assign _0800_ = ~ rs[5];
  assign _0801_ = _0799_ & _0800_;
  assign _0802_ = ~ rs[2];
  assign _0803_ = rs[9] & _0802_;
  assign _0804_ = _0801_ | _0803_;
  assign _0805_ = ~ rs[3];
  assign _0806_ = rs[9] & _0805_;
  assign _0807_ = _0804_ | _0806_;
  assign _0808_ = rs[8] & rs[6];
  assign _0809_ = _0808_ & rs[1];
  assign _0810_ = ~ rs[5];
  assign _0811_ = _0809_ & _0810_;
  assign _0812_ = ~ rs[2];
  assign _0813_ = rs[8] & _0812_;
  assign _0814_ = _0811_ | _0813_;
  assign _0815_ = ~ rs[3];
  assign _0816_ = rs[8] & _0815_;
  assign _0817_ = _0814_ | _0816_;
  assign _0818_ = ~ rs[2];
  assign _0819_ = rs[3] & _0818_;
  assign _0820_ = _0819_ & rs[1];
  assign _0821_ = rs[6] & rs[3];
  assign _0822_ = _0821_ & rs[2];
  assign _0823_ = _0822_ & rs[1];
  assign _0824_ = _0820_ | _0823_;
  assign _0825_ = ~ rs[5];
  assign _0826_ = _0825_ & rs[3];
  assign _0827_ = _0826_ & rs[2];
  assign _0828_ = _0827_ & rs[1];
  assign _0829_ = _0824_ | _0828_;
  assign _0830_ = rs[9] & rs[5];
  assign _0831_ = _0830_ & rs[3];
  assign _0832_ = _0831_ & rs[2];
  assign _0833_ = _0832_ & rs[1];
  assign _0834_ = ~ rs[6];
  assign _0835_ = _0833_ & _0834_;
  assign _0836_ = ~ rs[1];
  assign _0837_ = rs[6] & _0836_;
  assign _0838_ = _0837_ & rs[3];
  assign _0839_ = _0835_ | _0838_;
  assign _0840_ = ~ rs[3];
  assign _0841_ = rs[6] & _0840_;
  assign _0842_ = _0839_ | _0841_;
  assign _0843_ = rs[8] & rs[5];
  assign _0844_ = _0843_ & rs[2];
  assign _0845_ = _0844_ & rs[3];
  assign _0846_ = _0845_ & rs[1];
  assign _0847_ = ~ rs[6];
  assign _0848_ = _0846_ & _0847_;
  assign _0849_ = ~ rs[1];
  assign _0850_ = rs[5] & _0849_;
  assign _0851_ = _0850_ & rs[3];
  assign _0852_ = _0848_ | _0851_;
  assign _0853_ = ~ rs[3];
  assign _0854_ = rs[5] & _0853_;
  assign _0855_ = _0852_ | _0854_;
  assign _0856_ = rs[5] & rs[3];
  assign _0857_ = _0856_ & rs[2];
  assign _0858_ = _0857_ & rs[1];
  assign _0859_ = rs[6] & rs[3];
  assign _0860_ = _0859_ & rs[2];
  assign _0861_ = _0860_ & rs[1];
  assign _0862_ = _0858_ | _0861_;
  assign _0863_ = ~ rs[2];
  assign _0864_ = rs[3] & _0863_;
  assign _0865_ = ~ rs[1];
  assign _0866_ = _0864_ & _0865_;
  assign _0867_ = _0862_ | _0866_;
  assign _0868_ = ~ rs[6];
  assign _0869_ = rs[9] & _0868_;
  assign _0870_ = ~ rs[5];
  assign _0871_ = _0869_ & _0870_;
  assign _0872_ = _0871_ & rs[2];
  assign _0873_ = _0872_ & rs[3];
  assign _0874_ = rs[6] & rs[3];
  assign _0875_ = ~ rs[2];
  assign _0876_ = _0874_ & _0875_;
  assign _0877_ = _0876_ & rs[1];
  assign _0878_ = _0873_ | _0877_;
  assign _0879_ = rs[9] & rs[2];
  assign _0880_ = ~ rs[1];
  assign _0881_ = _0879_ & _0880_;
  assign _0882_ = _0881_ & rs[3];
  assign _0883_ = _0878_ | _0882_;
  assign _0884_ = ~ rs[3];
  assign _0885_ = rs[2] & _0884_;
  assign _0886_ = _0883_ | _0885_;
  assign _0887_ = ~ rs[6];
  assign _0888_ = rs[8] & _0887_;
  assign _0889_ = ~ rs[5];
  assign _0890_ = _0888_ & _0889_;
  assign _0891_ = _0890_ & rs[3];
  assign _0892_ = _0891_ & rs[2];
  assign _0893_ = rs[5] & rs[3];
  assign _0894_ = ~ rs[2];
  assign _0895_ = _0893_ & _0894_;
  assign _0896_ = _0895_ & rs[1];
  assign _0897_ = _0892_ | _0896_;
  assign _0898_ = rs[8] & rs[3];
  assign _0899_ = _0898_ & rs[2];
  assign _0900_ = ~ rs[1];
  assign _0901_ = _0899_ & _0900_;
  assign _0902_ = _0897_ | _0901_;
  assign _0903_ = ~ rs[3];
  assign _0904_ = rs[1] & _0903_;
  assign _0905_ = _0902_ | _0904_;
  assign _0906_ = _1156_ ? { 12'h000, _1167_, _1178_, rs[52], _1195_, _1212_, rs[48], _1214_, _1221_, _1228_, rs[44], _1239_, _1250_, rs[40], _1267_, _1284_, rs[36], _1286_, _1293_, _1300_, rs[32], 12'h000, _1311_, _1322_, rs[20], _1339_, _0341_, rs[16], _0343_, _0350_, _0357_, rs[12], _0368_, _0379_, rs[8], _0396_, _0413_, rs[4], _0415_, _0422_, _0429_, rs[0] } : { 8'h00, _0440_, _0450_, _0460_, rs[49], _0472_, _0485_, _0498_, rs[46], _0510_, _0529_, _0548_, rs[42], _0559_, _0569_, _0579_, rs[39], _0591_, _0604_, _0617_, rs[36], _0629_, _0648_, _0667_, rs[32], 8'h00, _0678_, _0688_, _0698_, rs[17], _0710_, _0723_, _0736_, rs[14], _0748_, _0767_, _0786_, rs[10], _0797_, _0807_, _0817_, rs[7], _0829_, _0842_, _0855_, rs[4], _0867_, _0886_, _0905_, rs[0] };
  assign _0907_ = op == 6'h3b;
  assign _0908_ = datalen[0] & rs[7];
  assign _0909_ = datalen[1] & rs[15];
  assign _0910_ = _0908_ | _0909_;
  assign _0911_ = datalen[2] & rs[31];
  assign _0912_ = _0910_ | _0911_;
  assign _0913_ = datalen[2] ? rs[31:16] : { _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_ };
  assign _0914_ = datalen[2] | datalen[1];
  assign _0915_ = _0914_ ? rs[15:8] : { _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_ };
  assign _0916_ = op == 6'h17;
  function [7:0] \30483 ;
    input [7:0] a;
    input [47:0] b;
    input [5:0] s;
    (* parallel_case *)
    casez (s)
      6'b?????1:
        \30483  = b[7:0];
      6'b????1?:
        \30483  = b[15:8];
      6'b???1??:
        \30483  = b[23:16];
      6'b??1???:
        \30483  = b[31:24];
      6'b?1????:
        \30483  = b[39:32];
      6'b1?????:
        \30483  = b[47:40];
      default:
        \30483  = a;
    endcase
  endfunction
  assign _0917_ = \30483 (rs[7:0], { rs[7:0], _0906_[7:0], permute, _1139_, parity[7:0], _1131_[7:0] }, { _0916_, _0907_, _1155_, _1154_, _1137_, _1136_ });
  function [7:0] \30490 ;
    input [7:0] a;
    input [47:0] b;
    input [5:0] s;
    (* parallel_case *)
    casez (s)
      6'b?????1:
        \30490  = b[7:0];
      6'b????1?:
        \30490  = b[15:8];
      6'b???1??:
        \30490  = b[23:16];
      6'b??1???:
        \30490  = b[31:24];
      6'b?1????:
        \30490  = b[39:32];
      6'b1?????:
        \30490  = b[47:40];
      default:
        \30490  = a;
    endcase
  endfunction
  assign _0918_ = \30490 (rs[15:8], { _0915_, _0906_[15:8], 8'h00, _1141_, parity[15:8], _1131_[15:8] }, { _0916_, _0907_, _1155_, _1154_, _1137_, _1136_ });
  function [15:0] \30497 ;
    input [15:0] a;
    input [95:0] b;
    input [5:0] s;
    (* parallel_case *)
    casez (s)
      6'b?????1:
        \30497  = b[15:0];
      6'b????1?:
        \30497  = b[31:16];
      6'b???1??:
        \30497  = b[47:32];
      6'b??1???:
        \30497  = b[63:48];
      6'b?1????:
        \30497  = b[79:64];
      6'b1?????:
        \30497  = b[95:80];
      default:
        \30497  = a;
    endcase
  endfunction
  assign _0919_ = \30497 (rs[31:16], { _0913_, _0906_[31:16], 16'h0000, _1145_, _1143_, parity[31:16], _1131_[31:16] }, { _0916_, _0907_, _1155_, _1154_, _1137_, _1136_ });
  function [31:0] \30504 ;
    input [31:0] a;
    input [191:0] b;
    input [5:0] s;
    (* parallel_case *)
    casez (s)
      6'b?????1:
        \30504  = b[31:0];
      6'b????1?:
        \30504  = b[63:32];
      6'b???1??:
        \30504  = b[95:64];
      6'b??1???:
        \30504  = b[127:96];
      6'b?1????:
        \30504  = b[159:128];
      6'b1?????:
        \30504  = b[191:160];
      default:
        \30504  = a;
    endcase
  endfunction
  assign _0920_ = \30504 (rs[63:32], { _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0912_, _0906_[63:32], 32'h00000000, _1153_, _1151_, _1149_, _1147_, parity[63:32], _1131_[63:32] }, { _0916_, _0907_, _1155_, _1154_, _1137_, _1136_ });
  assign par0 = _1091_;
  assign par1 = _1094_;
  assign parity = { 31'h00000000, _1097_, 31'h00000000, _1096_ };
  assign permute = { _1121_, _1118_, _1115_, _1112_, _1109_, _1106_, _1103_, _1100_ };
  assign result = { _0920_, _0919_, _0918_, _0917_ };
endmodule