module BTB
(
  clk,
  reset,
  io_req_valid,
  io_req_bits_addr,
  io_resp_valid,
  io_resp_bits_taken,
  io_resp_bits_mask,
  io_resp_bits_bridx,
  io_resp_bits_target,
  io_resp_bits_entry,
  io_resp_bits_bht_history,
  io_resp_bits_bht_value,
  io_btb_update_valid,
  io_btb_update_bits_prediction_valid,
  io_btb_update_bits_prediction_bits_taken,
  io_btb_update_bits_prediction_bits_mask,
  io_btb_update_bits_prediction_bits_bridx,
  io_btb_update_bits_prediction_bits_target,
  io_btb_update_bits_prediction_bits_entry,
  io_btb_update_bits_prediction_bits_bht_history,
  io_btb_update_bits_prediction_bits_bht_value,
  io_btb_update_bits_pc,
  io_btb_update_bits_target,
  io_btb_update_bits_taken,
  io_btb_update_bits_isJump,
  io_btb_update_bits_isReturn,
  io_btb_update_bits_br_pc,
  io_bht_update_valid,
  io_bht_update_bits_prediction_valid,
  io_bht_update_bits_prediction_bits_taken,
  io_bht_update_bits_prediction_bits_mask,
  io_bht_update_bits_prediction_bits_bridx,
  io_bht_update_bits_prediction_bits_target,
  io_bht_update_bits_prediction_bits_entry,
  io_bht_update_bits_prediction_bits_bht_history,
  io_bht_update_bits_prediction_bits_bht_value,
  io_bht_update_bits_pc,
  io_bht_update_bits_taken,
  io_bht_update_bits_mispredict,
  io_ras_update_valid,
  io_ras_update_bits_isCall,
  io_ras_update_bits_isReturn,
  io_ras_update_bits_returnAddr,
  io_ras_update_bits_prediction_valid,
  io_ras_update_bits_prediction_bits_taken,
  io_ras_update_bits_prediction_bits_mask,
  io_ras_update_bits_prediction_bits_bridx,
  io_ras_update_bits_prediction_bits_target,
  io_ras_update_bits_prediction_bits_entry,
  io_ras_update_bits_prediction_bits_bht_history,
  io_ras_update_bits_prediction_bits_bht_value,
  io_invalidate
);

  input [38:0] io_req_bits_addr;
  output [38:0] io_resp_bits_target;
  output [5:0] io_resp_bits_entry;
  output [6:0] io_resp_bits_bht_history;
  output [1:0] io_resp_bits_bht_value;
  input [38:0] io_btb_update_bits_prediction_bits_target;
  input [5:0] io_btb_update_bits_prediction_bits_entry;
  input [6:0] io_btb_update_bits_prediction_bits_bht_history;
  input [1:0] io_btb_update_bits_prediction_bits_bht_value;
  input [38:0] io_btb_update_bits_pc;
  input [38:0] io_btb_update_bits_target;
  input [38:0] io_btb_update_bits_br_pc;
  input [38:0] io_bht_update_bits_prediction_bits_target;
  input [5:0] io_bht_update_bits_prediction_bits_entry;
  input [6:0] io_bht_update_bits_prediction_bits_bht_history;
  input [1:0] io_bht_update_bits_prediction_bits_bht_value;
  input [38:0] io_bht_update_bits_pc;
  input [38:0] io_ras_update_bits_returnAddr;
  input [38:0] io_ras_update_bits_prediction_bits_target;
  input [5:0] io_ras_update_bits_prediction_bits_entry;
  input [6:0] io_ras_update_bits_prediction_bits_bht_history;
  input [1:0] io_ras_update_bits_prediction_bits_bht_value;
  input clk;
  input reset;
  input io_req_valid;
  input io_btb_update_valid;
  input io_btb_update_bits_prediction_valid;
  input io_btb_update_bits_prediction_bits_taken;
  input io_btb_update_bits_prediction_bits_mask;
  input io_btb_update_bits_prediction_bits_bridx;
  input io_btb_update_bits_taken;
  input io_btb_update_bits_isJump;
  input io_btb_update_bits_isReturn;
  input io_bht_update_valid;
  input io_bht_update_bits_prediction_valid;
  input io_bht_update_bits_prediction_bits_taken;
  input io_bht_update_bits_prediction_bits_mask;
  input io_bht_update_bits_prediction_bits_bridx;
  input io_bht_update_bits_taken;
  input io_bht_update_bits_mispredict;
  input io_ras_update_valid;
  input io_ras_update_bits_isCall;
  input io_ras_update_bits_isReturn;
  input io_ras_update_bits_prediction_valid;
  input io_ras_update_bits_prediction_bits_taken;
  input io_ras_update_bits_prediction_bits_mask;
  input io_ras_update_bits_prediction_bits_bridx;
  input io_invalidate;
  output io_resp_valid;
  output io_resp_bits_taken;
  output io_resp_bits_mask;
  output io_resp_bits_bridx;
  wire [38:0] io_resp_bits_target,T1535,T1995,T1536;
  wire [5:0] io_resp_bits_entry,T169,T172,T173,T189,idxPagesOH_0,pageHit,T266,T192,
  pageReplEn,idxPageReplEn,tgtPageReplEn,tgtPageRepl,T193,updatePageHit,idxPageRepl,T204,
  T262,T263,T291,idxPagesOH_1,T296,idxPagesOH_2,T300,idxPagesOH_3,T306,idxPagesOH_4,
  T310,idxPagesOH_5,T315,idxPagesOH_6,T319,idxPagesOH_7,T326,idxPagesOH_8,T330,
  idxPagesOH_9,T335,idxPagesOH_10,T339,idxPagesOH_11,T345,idxPagesOH_12,T349,
  idxPagesOH_13,T354,idxPagesOH_14,T358,idxPagesOH_15,T366,idxPagesOH_16,T370,
  idxPagesOH_17,T375,idxPagesOH_18,T379,idxPagesOH_19,T385,idxPagesOH_20,T389,idxPagesOH_21,
  T394,idxPagesOH_22,T398,idxPagesOH_23,T405,idxPagesOH_24,T409,idxPagesOH_25,T414,
  idxPagesOH_26,T418,idxPagesOH_27,T424,idxPagesOH_28,T428,idxPagesOH_29,T432,
  idxPagesOH_30,T441,idxPagesOH_31,T445,idxPagesOH_32,T450,idxPagesOH_33,T454,
  idxPagesOH_34,T460,idxPagesOH_35,T464,idxPagesOH_36,T469,idxPagesOH_37,T473,idxPagesOH_38,
  T480,idxPagesOH_39,T484,idxPagesOH_40,T489,idxPagesOH_41,T493,idxPagesOH_42,
  T499,idxPagesOH_43,T503,idxPagesOH_44,T508,idxPagesOH_45,T512,idxPagesOH_46,T520,
  idxPagesOH_47,T524,idxPagesOH_48,T529,idxPagesOH_49,T533,idxPagesOH_50,T539,
  idxPagesOH_51,T543,idxPagesOH_52,T548,idxPagesOH_53,T552,idxPagesOH_54,T559,
  idxPagesOH_55,T563,idxPagesOH_56,T568,idxPagesOH_57,T572,idxPagesOH_58,T578,idxPagesOH_59,
  T582,idxPagesOH_60,T586,idxPagesOH_61,T794,T795,tgtPagesOH_0,T803,T804,
  tgtPagesOH_1,T809,T810,tgtPagesOH_2,T814,T815,tgtPagesOH_3,T821,T822,tgtPagesOH_4,T826,
  T827,tgtPagesOH_5,T832,T833,tgtPagesOH_6,T837,T838,tgtPagesOH_7,T845,T846,
  tgtPagesOH_8,T850,T851,tgtPagesOH_9,T856,T857,tgtPagesOH_10,T861,T862,tgtPagesOH_11,T868,
  T869,tgtPagesOH_12,T873,T874,tgtPagesOH_13,T879,T880,tgtPagesOH_14,T884,T885,
  tgtPagesOH_15,T893,T894,tgtPagesOH_16,T898,T899,tgtPagesOH_17,T904,T905,
  tgtPagesOH_18,T909,T910,tgtPagesOH_19,T916,T917,tgtPagesOH_20,T921,T922,tgtPagesOH_21,T927,
  T928,tgtPagesOH_22,T932,T933,tgtPagesOH_23,T940,T941,tgtPagesOH_24,T945,T946,
  tgtPagesOH_25,T951,T952,tgtPagesOH_26,T956,T957,tgtPagesOH_27,T963,T964,
  tgtPagesOH_28,T968,T969,tgtPagesOH_29,T973,T974,tgtPagesOH_30,T983,T984,tgtPagesOH_31,T988,
  T989,tgtPagesOH_32,T994,T995,tgtPagesOH_33,T999,T1000,tgtPagesOH_34,T1006,T1007,
  tgtPagesOH_35,T1011,T1012,tgtPagesOH_36,T1017,T1018,tgtPagesOH_37,T1022,T1023,
  tgtPagesOH_38,T1030,T1031,tgtPagesOH_39,T1035,T1036,tgtPagesOH_40,T1041,T1042,
  tgtPagesOH_41,T1046,T1047,tgtPagesOH_42,T1053,T1054,tgtPagesOH_43,T1058,T1059,
  tgtPagesOH_44,T1064,T1065,tgtPagesOH_45,T1069,T1070,tgtPagesOH_46,T1078,T1079,
  tgtPagesOH_47,T1083,T1084,tgtPagesOH_48,T1089,T1090,tgtPagesOH_49,T1094,T1095,
  tgtPagesOH_50,T1101,T1102,tgtPagesOH_51,T1106,T1107,tgtPagesOH_52,T1112,T1113,
  tgtPagesOH_53,T1117,T1118,tgtPagesOH_54,T1125,T1126,tgtPagesOH_55,T1130,T1131,tgtPagesOH_56,
  T1136,T1137,tgtPagesOH_57,T1141,T1142,tgtPagesOH_58,T1148,T1149,tgtPagesOH_59,
  T1153,T1154,tgtPagesOH_60,T1158,T1159,tgtPagesOH_61,T1791,T1794,T1792,T1797,T1795,
  T1800,T1798,T1803,T1801,T1806,T1804,T1809,T1807,T1812,T1810,T1815,T1813,T1818,
  T1816,T1821,T1819,T1824,T1822,T1827,T1825,T1830,T1828,T1833,T1831,T1836,T1834,
  T1839,T1837,T1842,T1840,T1845,T1843,T1848,T1846,T1851,T1849,T1854,T1852,T1857,T1855,
  T1860,T1858,T1863,T1861,T1866,T1864,T1869,T1867,T1872,T1870,T1875,T1873,T1878,
  T1876,T1881,T1879,T1884,T1882,T1887,T1885,T1890,T1888,T1893,T1891,T1896,T1894,
  T1899,T1897,T1902,T1900,T1905,T1903,T1908,T1906,T1911,T1909,T1914,T1912,T1917,T1915,
  T1920,T1918,T1923,T1921,T1926,T1924,T1929,T1927,T1932,T1930,T1935,T1933,T1938,
  T1936,T1941,T1939,T1944,T1942,T1947,T1945,T1950,T1948,T1953,T1951,T1956,T1954,
  T1959,T1957,T1962,T1960,T1965,T1963,T1968,T1966,T1971,T1969,T1974,T1972;
  wire [1:0] io_resp_bits_bht_value,T2000,T2017,T2014;
  wire io_resp_valid,io_resp_bits_taken,io_resp_bits_mask,io_resp_bits_bridx,N0,N1,N2,
  N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,
  N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,
  N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,
  N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,
  N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,
  N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,
  N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,
  N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,
  N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,
  N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,
  N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,
  N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,
  N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,
  N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,
  N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,
  N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
  N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,
  N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,
  N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,
  N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
  N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,
  N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,
  N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,
  N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,
  N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,
  N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,
  N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,
  N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,
  N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,
  N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,
  N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
  N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,
  N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,
  N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,
  N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
  N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,
  N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,
  N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,
  N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,
  N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,
  N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,
  N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,
  N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,
  N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,
  N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
  N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,
  N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,
  N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,
  N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,
  N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,
  N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,
  N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,
  N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,
  N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,
  N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,
  N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,
  N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,
  N936,N937,N938,N939,T18,T14,T15,T21,T1530,T159,T1527,T160,T161,T1162,T162,N940,
  T166,N941,T175,T176,T265,doTgtPageRepl,N942,samePage,N943,N944,T203,doPageRepl,
  doIdxPageRepl,N945,T220,T219,T222,T225,T224,T229,T228,T236,T235,T238,T241,T240,
  T245,T244,T264,T261,N946,T289,T288,T602,T601,N947,N948,N949,T801,T800,T1168,T1163,
  N950,T1165,T1174,T1169,N951,T1171,T1180,T1175,N952,T1177,T1186,T1181,N953,T1183,
  T1192,T1187,N954,T1189,T1198,T1193,N955,T1195,T1204,T1199,N956,T1201,T1210,T1205,
  N957,T1207,T1216,T1211,N958,T1213,T1222,T1217,N959,T1219,T1228,T1223,N960,T1225,
  T1234,T1229,N961,T1231,T1240,T1235,N962,T1237,T1246,T1241,N963,T1243,T1252,
  T1247,N964,T1249,T1258,T1253,N965,T1255,T1264,T1259,N966,T1261,T1270,T1265,N967,
  T1267,T1276,T1271,N968,T1273,T1282,T1277,N969,T1279,T1288,T1283,N970,T1285,T1294,
  T1289,N971,T1291,T1300,T1295,N972,T1297,T1306,T1301,N973,T1303,T1312,T1307,N974,
  T1309,T1318,T1313,N975,T1315,T1324,T1319,N976,T1321,T1330,T1325,N977,T1327,T1336,
  T1331,N978,T1333,T1342,T1337,N979,T1339,T1348,T1343,N980,T1345,T1354,T1349,N981,
  T1351,T1360,T1355,N982,T1357,T1366,T1361,N983,T1363,T1372,T1367,N984,T1369,T1378,
  T1373,N985,T1375,T1384,T1379,N986,T1381,T1390,T1385,N987,T1387,T1396,T1391,N988,
  T1393,T1402,T1397,N989,T1399,T1408,T1403,N990,T1405,T1414,T1409,N991,T1411,T1420,
  T1415,N992,T1417,T1426,T1421,N993,T1423,T1432,T1427,N994,T1429,T1438,T1433,N995,
  T1435,T1444,T1439,N996,T1441,T1450,T1445,N997,T1447,T1456,T1451,N998,T1453,T1462,
  T1457,N999,T1459,T1468,T1463,N1000,T1465,T1474,T1469,N1001,T1471,T1480,T1475,
  N1002,T1477,T1486,T1481,N1003,T1483,T1492,T1487,N1004,T1489,T1498,T1493,N1005,
  T1495,T1504,T1499,N1006,T1501,T1510,T1505,N1007,T1507,T1516,T1511,N1008,T1513,T1522,
  T1517,N1009,T1519,N1010,T1524,T2406,N1011,T2028,N1012,T1542,T1541,N1013,N1014,
  N1015,N1016,N1017,N1018,N1019,T1998,T2022,T2001,T2007,T2006,T2018,T2008,T2015,
  T2016,T2019,T2021,T2020,T2025,T2404,T2029,T2039,T2030,T2034,T2045,T2040,T2042,T2051,
  T2046,T2048,T2057,T2052,T2054,T2063,T2058,T2060,T2069,T2064,T2066,T2075,T2070,
  T2072,T2081,T2076,T2078,T2087,T2082,T2084,T2093,T2088,T2090,T2099,T2094,T2096,
  T2105,T2100,T2102,T2111,T2106,T2108,T2117,T2112,T2114,T2123,T2118,T2120,T2129,T2124,
  T2126,T2135,T2130,T2132,T2141,T2136,T2138,T2147,T2142,T2144,T2153,T2148,T2150,
  T2159,T2154,T2156,T2165,T2160,T2162,T2171,T2166,T2168,T2177,T2172,T2174,T2183,
  T2178,T2180,T2189,T2184,T2186,T2195,T2190,T2192,T2201,T2196,T2198,T2207,T2202,T2204,
  T2213,T2208,T2210,T2219,T2214,T2216,T2225,T2220,T2222,T2231,T2226,T2228,T2237,
  T2232,T2234,T2243,T2238,T2240,T2249,T2244,T2246,T2255,T2250,T2252,T2261,T2256,
  T2258,T2267,T2262,T2264,T2273,T2268,T2270,T2279,T2274,T2276,T2285,T2280,T2282,T2291,
  T2286,T2288,T2297,T2292,T2294,T2303,T2298,T2300,T2309,T2304,T2306,T2315,T2310,
  T2312,T2321,T2316,T2318,T2327,T2322,T2324,T2333,T2328,T2330,T2339,T2334,T2336,
  T2345,T2340,T2342,T2351,T2346,T2348,T2357,T2352,T2354,T2363,T2358,T2360,T2369,T2364,
  T2366,T2375,T2370,T2372,T2381,T2376,T2378,T2387,T2382,T2384,T2393,T2388,T2390,
  T2399,T2394,T2396,T2401,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,
  N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,
  N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,
  N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,
  N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,T2410,
  T2409,T2412,N1082,T2413,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,
  N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,
  N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,
  N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,
  N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,
  N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,N1198,
  N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,N1211,
  N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1238,
  N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,N1251,
  N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,N1278,
  N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,N1291,
  N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,N1318,
  N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,N1331,
  N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,N1358,
  N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,N1371,
  N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,N1398,
  N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,N1411,
  N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,N1438,
  N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,N1451,
  N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478,
  N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,
  N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,N1518,
  N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531,
  N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,N1558,
  N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571,
  N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,N1598,
  N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,N1611,
  N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638,
  N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1651,
  N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678,
  N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,N1691,
  N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718,
  N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,N1731,
  N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,N1758,
  N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1771,
  N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,
  N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,N1811,
  N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838,
  N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,N1851,
  N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878,
  N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,N1891,
  N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
  N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,N1931,
  N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958,
  N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,N1971,
  N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998,
  N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,N2011,
  N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038,
  N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,N2051,
  N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078,
  N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,N2091,
  N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118,
  N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,N2131,
  N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,
  N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,N2171,
  N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198,
  N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211,
  N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,
  N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251,
  N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278,
  N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,N2291,
  N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
  N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331,
  N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358,
  N2359,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,
  N2373,N2374,N2376,N2377,N2378,N2379,N2380,N2381,N2383,N2384,N2385,N2386,N2387,
  N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2402,
  N2403,N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,
  N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,
  N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,
  N2444,N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,
  N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,N2466,N2467,N2468,N2469,N2470,
  N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,
  N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,
  N2498,N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,
  N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,
  N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,
  N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,
  N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,
  N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,
  N2578,N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,
  N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,
  N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,
  N2618,N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,
  N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,
  N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,
  N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,
  N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,
  N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,
  N2698,N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,
  N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,
  N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,
  N2738,N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,
  N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,
  N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,
  N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,
  N2791,N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,
  N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,
  N2818,N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,
  N2831,N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,
  N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,
  N2858,N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,
  N2871,N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,
  N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,
  N2898,N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,
  N2911,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,
  N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,
  N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,
  N2951,N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,
  N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,
  N2978,N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,
  N2991,N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,
  N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,
  N3018,N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,
  N3031,N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,
  N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,
  N3058,N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,
  N3071,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,
  N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,
  N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,
  N3111,N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,
  N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,
  N3138,N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,
  N3151,N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,
  N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,
  N3178,N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,
  N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,
  N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,
  N3218,N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,
  N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,
  N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,
  N3258;
  wire [6:0] T152,T22;
  wire [0:0] T12,T2420,T2423,T2439;
  wire [61:0] T168,hits,T589,T590,T2435,T780,T782,T2438,T783,T785,T2036;
  wire [5:1] T195;
  wire [2:0] T200,T201;
  wire [26:0] T214,T232,T1976,T1788,T1980,T1977,T1984,T1981,T1988,T1985,T1992,T1989;
  wire [1:1] T2427,T2443,T2445,T2457;
  wire [3:2] T2444,T2458;
  wire [5:4] T799;
  wire [3:1] T2459;
  wire [7:4] T2460;
  wire [7:1] T2461;
  wire [15:8] T2462;
  wire [15:1] T2463;
  wire [29:16] T2464;
  wire [11:0] T1544,T1538,T1548,T1545,T1552,T1549,T1556,T1553,T1560,T1557,T1564,T1561,T1568,
  T1565,T1572,T1569,T1576,T1573,T1580,T1577,T1584,T1581,T1588,T1585,T1592,T1589,
  T1596,T1593,T1600,T1597,T1604,T1601,T1608,T1605,T1612,T1609,T1616,T1613,T1620,T1617,
  T1624,T1621,T1628,T1625,T1632,T1629,T1636,T1633,T1640,T1637,T1644,T1641,T1648,
  T1645,T1652,T1649,T1656,T1653,T1660,T1657,T1664,T1661,T1668,T1665,T1672,T1669,
  T1676,T1673,T1680,T1677,T1684,T1681,T1688,T1685,T1692,T1689,T1696,T1693,T1700,T1697,
  T1704,T1701,T1708,T1705,T1712,T1709,T1716,T1713,T1720,T1717,T1724,T1721,T1728,
  T1725,T1732,T1729,T1736,T1733,T1740,T1737,T1744,T1741,T1748,T1745,T1752,T1749,
  T1756,T1753,T1760,T1757,T1764,T1761,T1768,T1765,T1772,T1769,T1776,T1773,T1780,T1777,
  T1784,T1781;
  reg R7,isJump_61,R164,updateHit,isJump_60,isJump_59,isJump_58,isJump_57,isJump_56,
  isJump_55,isJump_54,isJump_53,isJump_52,isJump_51,isJump_50,isJump_49,isJump_48,
  isJump_47,isJump_46,isJump_45,isJump_44,isJump_43,isJump_42,isJump_41,isJump_40,
  isJump_39,isJump_38,isJump_37,isJump_36,isJump_35,isJump_34,isJump_33,isJump_32,
  isJump_31,isJump_30,isJump_29,isJump_28,isJump_27,isJump_26,isJump_25,isJump_24,
  isJump_23,isJump_22,isJump_21,isJump_20,isJump_19,isJump_18,isJump_17,isJump_16,
  isJump_15,isJump_14,isJump_13,isJump_12,isJump_11,isJump_10,isJump_9,isJump_8,
  isJump_7,isJump_6,isJump_5,isJump_4,isJump_3,isJump_2,isJump_1,isJump_0,T2027,
  useRAS_61,R2032,useRAS_60,useRAS_59,useRAS_58,useRAS_57,useRAS_56,useRAS_55,useRAS_54,
  useRAS_53,useRAS_52,useRAS_51,useRAS_50,useRAS_49,useRAS_48,useRAS_47,useRAS_46,
  useRAS_45,useRAS_44,useRAS_43,useRAS_42,useRAS_41,useRAS_40,useRAS_39,useRAS_38,
  useRAS_37,useRAS_36,useRAS_35,useRAS_34,useRAS_33,useRAS_32,useRAS_31,useRAS_30,
  useRAS_29,useRAS_28,useRAS_27,useRAS_26,useRAS_25,useRAS_24,useRAS_23,useRAS_22,
  useRAS_21,useRAS_20,useRAS_19,useRAS_18,useRAS_17,useRAS_16,useRAS_15,useRAS_14,
  useRAS_13,useRAS_12,useRAS_11,useRAS_10,useRAS_9,useRAS_8,useRAS_7,useRAS_6,
  useRAS_5,useRAS_4,useRAS_3,useRAS_2,useRAS_1,useRAS_0;
  reg [255:0] T10;
  reg [6:0] io_resp_bits_bht_history;
  reg [5:0] nextRepl,R177,pageValid;
  reg [2:0] R198,T588,T584,T580,T574,T570,T565,T561,T554,T550,T545,T541,T535,T531,T526,T522,
  T514,T510,T505,T501,T495,T491,T486,T482,T475,T471,T466,T462,T456,T452,T447,T443,
  T434,T430,T426,T420,T416,T411,T407,T400,T396,T391,T387,T381,T377,T372,T368,T360,
  T356,T351,T347,T341,T337,T332,T328,T321,T317,T312,T308,T302,T298,T293,T286,
  T1161,T1156,T1151,T1144,T1139,T1133,T1128,T1120,T1115,T1109,T1104,T1097,T1092,T1086,
  T1081,T1072,T1067,T1061,T1056,T1049,T1044,T1038,T1033,T1025,T1020,T1014,T1009,
  T1002,T997,T991,T986,T976,T971,T966,T959,T954,T948,T943,T935,T930,T924,T919,T912,
  T907,T901,T896,T887,T882,T876,T871,T864,T859,T853,T848,T840,T835,T829,T824,T817,
  T812,T806,T797;
  reg [26:0] T209,T258,T256,T254,T250,T248,T212;
  reg [11:0] T2434,T779,T777,T775,T771,T769,T766,T764,T759,T757,T754,T752,T748,T746,T743,
  T741,T735,T733,T730,T728,T724,T722,T719,T717,T712,T710,T707,T705,T701,T699,T696,
  T694,T687,T685,T683,T679,T677,T674,T672,T667,T665,T662,T660,T656,T654,T651,T649,
  T643,T641,T638,T636,T632,T630,T627,T625,T620,T618,T615,T613,T609,T607,T604,T599,
  T1539,T1546,T1550,T1554,T1558,T1562,T1566,T1570,T1574,T1578,T1582,T1586,T1590,T1594,
  T1598,T1602,T1606,T1610,T1614,T1618,T1622,T1626,T1630,T1634,T1638,T1642,T1646,
  T1650,T1654,T1658,T1662,T1666,T1670,T1674,T1678,T1682,T1686,T1690,T1694,T1698,
  T1702,T1706,T1710,T1714,T1718,T1722,T1726,T1730,T1734,T1738,T1742,T1746,T1750,T1754,
  T1758,T1762,T1766,T1770,T1774,T1778,T1782,T1785;
  reg [61:0] T2437,brIdx;
  reg [38:0] R1996,R2023;
  reg [1:0] R2010;
  assign io_resp_bits_mask = 1'b1;
  assign io_resp_bits_bht_value[1] = (N812)? T10[1] : 
                                     (N814)? T10[3] : 
                                     (N816)? T10[5] : 
                                     (N818)? T10[7] : 
                                     (N820)? T10[9] : 
                                     (N822)? T10[11] : 
                                     (N824)? T10[13] : 
                                     (N826)? T10[15] : 
                                     (N828)? T10[17] : 
                                     (N830)? T10[19] : 
                                     (N832)? T10[21] : 
                                     (N834)? T10[23] : 
                                     (N836)? T10[25] : 
                                     (N838)? T10[27] : 
                                     (N840)? T10[29] : 
                                     (N842)? T10[31] : 
                                     (N844)? T10[33] : 
                                     (N846)? T10[35] : 
                                     (N848)? T10[37] : 
                                     (N850)? T10[39] : 
                                     (N852)? T10[41] : 
                                     (N854)? T10[43] : 
                                     (N856)? T10[45] : 
                                     (N858)? T10[47] : 
                                     (N860)? T10[49] : 
                                     (N862)? T10[51] : 
                                     (N864)? T10[53] : 
                                     (N866)? T10[55] : 
                                     (N868)? T10[57] : 
                                     (N870)? T10[59] : 
                                     (N872)? T10[61] : 
                                     (N874)? T10[63] : 
                                     (N876)? T10[65] : 
                                     (N878)? T10[67] : 
                                     (N880)? T10[69] : 
                                     (N882)? T10[71] : 
                                     (N884)? T10[73] : 
                                     (N886)? T10[75] : 
                                     (N888)? T10[77] : 
                                     (N890)? T10[79] : 
                                     (N892)? T10[81] : 
                                     (N894)? T10[83] : 
                                     (N896)? T10[85] : 
                                     (N898)? T10[87] : 
                                     (N900)? T10[89] : 
                                     (N902)? T10[91] : 
                                     (N904)? T10[93] : 
                                     (N906)? T10[95] : 
                                     (N908)? T10[97] : 
                                     (N910)? T10[99] : 
                                     (N912)? T10[101] : 
                                     (N914)? T10[103] : 
                                     (N916)? T10[105] : 
                                     (N918)? T10[107] : 
                                     (N920)? T10[109] : 
                                     (N922)? T10[111] : 
                                     (N924)? T10[113] : 
                                     (N926)? T10[115] : 
                                     (N928)? T10[117] : 
                                     (N930)? T10[119] : 
                                     (N932)? T10[121] : 
                                     (N934)? T10[123] : 
                                     (N936)? T10[125] : 
                                     (N938)? T10[127] : 
                                     (N813)? T10[129] : 
                                     (N815)? T10[131] : 
                                     (N817)? T10[133] : 
                                     (N819)? T10[135] : 
                                     (N821)? T10[137] : 
                                     (N823)? T10[139] : 
                                     (N825)? T10[141] : 
                                     (N827)? T10[143] : 
                                     (N829)? T10[145] : 
                                     (N831)? T10[147] : 
                                     (N833)? T10[149] : 
                                     (N835)? T10[151] : 
                                     (N837)? T10[153] : 
                                     (N839)? T10[155] : 
                                     (N841)? T10[157] : 
                                     (N843)? T10[159] : 
                                     (N845)? T10[161] : 
                                     (N847)? T10[163] : 
                                     (N849)? T10[165] : 
                                     (N851)? T10[167] : 
                                     (N853)? T10[169] : 
                                     (N855)? T10[171] : 
                                     (N857)? T10[173] : 
                                     (N859)? T10[175] : 
                                     (N861)? T10[177] : 
                                     (N863)? T10[179] : 
                                     (N865)? T10[181] : 
                                     (N867)? T10[183] : 
                                     (N869)? T10[185] : 
                                     (N871)? T10[187] : 
                                     (N873)? T10[189] : 
                                     (N875)? T10[191] : 
                                     (N877)? T10[193] : 
                                     (N879)? T10[195] : 
                                     (N881)? T10[197] : 
                                     (N883)? T10[199] : 
                                     (N885)? T10[201] : 
                                     (N887)? T10[203] : 
                                     (N889)? T10[205] : 
                                     (N891)? T10[207] : 
                                     (N893)? T10[209] : 
                                     (N895)? T10[211] : 
                                     (N897)? T10[213] : 
                                     (N899)? T10[215] : 
                                     (N901)? T10[217] : 
                                     (N903)? T10[219] : 
                                     (N905)? T10[221] : 
                                     (N907)? T10[223] : 
                                     (N909)? T10[225] : 
                                     (N911)? T10[227] : 
                                     (N913)? T10[229] : 
                                     (N915)? T10[231] : 
                                     (N917)? T10[233] : 
                                     (N919)? T10[235] : 
                                     (N921)? T10[237] : 
                                     (N923)? T10[239] : 
                                     (N925)? T10[241] : 
                                     (N927)? T10[243] : 
                                     (N929)? T10[245] : 
                                     (N931)? T10[247] : 
                                     (N933)? T10[249] : 
                                     (N935)? T10[251] : 
                                     (N937)? T10[253] : 
                                     (N939)? T10[255] : 1'b0;
  assign io_resp_bits_bht_value[0] = (N812)? T10[0] : 
                                     (N814)? T10[2] : 
                                     (N816)? T10[4] : 
                                     (N818)? T10[6] : 
                                     (N820)? T10[8] : 
                                     (N822)? T10[10] : 
                                     (N824)? T10[12] : 
                                     (N826)? T10[14] : 
                                     (N828)? T10[16] : 
                                     (N830)? T10[18] : 
                                     (N832)? T10[20] : 
                                     (N834)? T10[22] : 
                                     (N836)? T10[24] : 
                                     (N838)? T10[26] : 
                                     (N840)? T10[28] : 
                                     (N842)? T10[30] : 
                                     (N844)? T10[32] : 
                                     (N846)? T10[34] : 
                                     (N848)? T10[36] : 
                                     (N850)? T10[38] : 
                                     (N852)? T10[40] : 
                                     (N854)? T10[42] : 
                                     (N856)? T10[44] : 
                                     (N858)? T10[46] : 
                                     (N860)? T10[48] : 
                                     (N862)? T10[50] : 
                                     (N864)? T10[52] : 
                                     (N866)? T10[54] : 
                                     (N868)? T10[56] : 
                                     (N870)? T10[58] : 
                                     (N872)? T10[60] : 
                                     (N874)? T10[62] : 
                                     (N876)? T10[64] : 
                                     (N878)? T10[66] : 
                                     (N880)? T10[68] : 
                                     (N882)? T10[70] : 
                                     (N884)? T10[72] : 
                                     (N886)? T10[74] : 
                                     (N888)? T10[76] : 
                                     (N890)? T10[78] : 
                                     (N892)? T10[80] : 
                                     (N894)? T10[82] : 
                                     (N896)? T10[84] : 
                                     (N898)? T10[86] : 
                                     (N900)? T10[88] : 
                                     (N902)? T10[90] : 
                                     (N904)? T10[92] : 
                                     (N906)? T10[94] : 
                                     (N908)? T10[96] : 
                                     (N910)? T10[98] : 
                                     (N912)? T10[100] : 
                                     (N914)? T10[102] : 
                                     (N916)? T10[104] : 
                                     (N918)? T10[106] : 
                                     (N920)? T10[108] : 
                                     (N922)? T10[110] : 
                                     (N924)? T10[112] : 
                                     (N926)? T10[114] : 
                                     (N928)? T10[116] : 
                                     (N930)? T10[118] : 
                                     (N932)? T10[120] : 
                                     (N934)? T10[122] : 
                                     (N936)? T10[124] : 
                                     (N938)? T10[126] : 
                                     (N813)? T10[128] : 
                                     (N815)? T10[130] : 
                                     (N817)? T10[132] : 
                                     (N819)? T10[134] : 
                                     (N821)? T10[136] : 
                                     (N823)? T10[138] : 
                                     (N825)? T10[140] : 
                                     (N827)? T10[142] : 
                                     (N829)? T10[144] : 
                                     (N831)? T10[146] : 
                                     (N833)? T10[148] : 
                                     (N835)? T10[150] : 
                                     (N837)? T10[152] : 
                                     (N839)? T10[154] : 
                                     (N841)? T10[156] : 
                                     (N843)? T10[158] : 
                                     (N845)? T10[160] : 
                                     (N847)? T10[162] : 
                                     (N849)? T10[164] : 
                                     (N851)? T10[166] : 
                                     (N853)? T10[168] : 
                                     (N855)? T10[170] : 
                                     (N857)? T10[172] : 
                                     (N859)? T10[174] : 
                                     (N861)? T10[176] : 
                                     (N863)? T10[178] : 
                                     (N865)? T10[180] : 
                                     (N867)? T10[182] : 
                                     (N869)? T10[184] : 
                                     (N871)? T10[186] : 
                                     (N873)? T10[188] : 
                                     (N875)? T10[190] : 
                                     (N877)? T10[192] : 
                                     (N879)? T10[194] : 
                                     (N881)? T10[196] : 
                                     (N883)? T10[198] : 
                                     (N885)? T10[200] : 
                                     (N887)? T10[202] : 
                                     (N889)? T10[204] : 
                                     (N891)? T10[206] : 
                                     (N893)? T10[208] : 
                                     (N895)? T10[210] : 
                                     (N897)? T10[212] : 
                                     (N899)? T10[214] : 
                                     (N901)? T10[216] : 
                                     (N903)? T10[218] : 
                                     (N905)? T10[220] : 
                                     (N907)? T10[222] : 
                                     (N909)? T10[224] : 
                                     (N911)? T10[226] : 
                                     (N913)? T10[228] : 
                                     (N915)? T10[230] : 
                                     (N917)? T10[232] : 
                                     (N919)? T10[234] : 
                                     (N921)? T10[236] : 
                                     (N923)? T10[238] : 
                                     (N925)? T10[240] : 
                                     (N927)? T10[242] : 
                                     (N929)? T10[244] : 
                                     (N931)? T10[246] : 
                                     (N933)? T10[248] : 
                                     (N935)? T10[250] : 
                                     (N937)? T10[252] : 
                                     (N939)? T10[254] : 1'b0;
  assign T204[0] = T212 == T209;
  assign T204[1] = T248 == T209;
  assign T204[2] = T250 == T209;
  assign T204[3] = T254 == T209;
  assign T204[4] = T256 == T209;
  assign T204[5] = T258 == T209;
  assign samePage = T209 == io_req_bits_addr[38:12];
  assign T266[0] = T212 == io_req_bits_addr[38:12];
  assign T266[1] = T248 == io_req_bits_addr[38:12];
  assign T266[2] = T250 == io_req_bits_addr[38:12];
  assign T266[3] = T254 == io_req_bits_addr[38:12];
  assign T266[4] = T256 == io_req_bits_addr[38:12];
  assign T266[5] = T258 == io_req_bits_addr[38:12];
  assign T289 = T169 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign T590[0] = T599 == io_req_bits_addr[11:0];
  assign T602 = T169 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign T590[1] = T604 == io_req_bits_addr[11:0];
  assign T590[2] = T607 == io_req_bits_addr[11:0];
  assign T590[3] = T609 == io_req_bits_addr[11:0];
  assign T590[4] = T613 == io_req_bits_addr[11:0];
  assign T590[5] = T615 == io_req_bits_addr[11:0];
  assign T590[6] = T618 == io_req_bits_addr[11:0];
  assign T590[7] = T620 == io_req_bits_addr[11:0];
  assign T590[8] = T625 == io_req_bits_addr[11:0];
  assign T590[9] = T627 == io_req_bits_addr[11:0];
  assign T590[10] = T630 == io_req_bits_addr[11:0];
  assign T590[11] = T632 == io_req_bits_addr[11:0];
  assign T590[12] = T636 == io_req_bits_addr[11:0];
  assign T590[13] = T638 == io_req_bits_addr[11:0];
  assign T590[14] = T641 == io_req_bits_addr[11:0];
  assign T590[15] = T643 == io_req_bits_addr[11:0];
  assign T590[16] = T649 == io_req_bits_addr[11:0];
  assign T590[17] = T651 == io_req_bits_addr[11:0];
  assign T590[18] = T654 == io_req_bits_addr[11:0];
  assign T590[19] = T656 == io_req_bits_addr[11:0];
  assign T590[20] = T660 == io_req_bits_addr[11:0];
  assign T590[21] = T662 == io_req_bits_addr[11:0];
  assign T590[22] = T665 == io_req_bits_addr[11:0];
  assign T590[23] = T667 == io_req_bits_addr[11:0];
  assign T590[24] = T672 == io_req_bits_addr[11:0];
  assign T590[25] = T674 == io_req_bits_addr[11:0];
  assign T590[26] = T677 == io_req_bits_addr[11:0];
  assign T590[27] = T679 == io_req_bits_addr[11:0];
  assign T590[28] = T683 == io_req_bits_addr[11:0];
  assign T590[29] = T685 == io_req_bits_addr[11:0];
  assign T590[30] = T687 == io_req_bits_addr[11:0];
  assign T590[31] = T694 == io_req_bits_addr[11:0];
  assign T590[32] = T696 == io_req_bits_addr[11:0];
  assign T590[33] = T699 == io_req_bits_addr[11:0];
  assign T590[34] = T701 == io_req_bits_addr[11:0];
  assign T590[35] = T705 == io_req_bits_addr[11:0];
  assign T590[36] = T707 == io_req_bits_addr[11:0];
  assign T590[37] = T710 == io_req_bits_addr[11:0];
  assign T590[38] = T712 == io_req_bits_addr[11:0];
  assign T590[39] = T717 == io_req_bits_addr[11:0];
  assign T590[40] = T719 == io_req_bits_addr[11:0];
  assign T590[41] = T722 == io_req_bits_addr[11:0];
  assign T590[42] = T724 == io_req_bits_addr[11:0];
  assign T590[43] = T728 == io_req_bits_addr[11:0];
  assign T590[44] = T730 == io_req_bits_addr[11:0];
  assign T590[45] = T733 == io_req_bits_addr[11:0];
  assign T590[46] = T735 == io_req_bits_addr[11:0];
  assign T590[47] = T741 == io_req_bits_addr[11:0];
  assign T590[48] = T743 == io_req_bits_addr[11:0];
  assign T590[49] = T746 == io_req_bits_addr[11:0];
  assign T590[50] = T748 == io_req_bits_addr[11:0];
  assign T590[51] = T752 == io_req_bits_addr[11:0];
  assign T590[52] = T754 == io_req_bits_addr[11:0];
  assign T590[53] = T757 == io_req_bits_addr[11:0];
  assign T590[54] = T759 == io_req_bits_addr[11:0];
  assign T590[55] = T764 == io_req_bits_addr[11:0];
  assign T590[56] = T766 == io_req_bits_addr[11:0];
  assign T590[57] = T769 == io_req_bits_addr[11:0];
  assign T590[58] = T771 == io_req_bits_addr[11:0];
  assign T590[59] = T775 == io_req_bits_addr[11:0];
  assign T590[60] = T777 == io_req_bits_addr[11:0];
  assign T590[61] = T779 == io_req_bits_addr[11:0];
  assign T801 = T169 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign T1542 = T169 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };
  assign T2000 = { 1'b0, 1'b1 } << T2001;
  assign T2410 = T169 < { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0 };

  always @(posedge clk) begin
    if(1'b1) begin
      R7 <= N1084;
    end 
  end


  always @(posedge clk) begin
    if(N1342) begin
      T10[255] <= N1344;
    end 
  end


  always @(posedge clk) begin
    if(N1342) begin
      T10[254] <= N1343;
    end 
  end


  always @(posedge clk) begin
    if(N1345) begin
      T10[253] <= N1347;
    end 
  end


  always @(posedge clk) begin
    if(N1345) begin
      T10[252] <= N1346;
    end 
  end


  always @(posedge clk) begin
    if(N1348) begin
      T10[251] <= N1350;
    end 
  end


  always @(posedge clk) begin
    if(N1348) begin
      T10[250] <= N1349;
    end 
  end


  always @(posedge clk) begin
    if(N1351) begin
      T10[249] <= N1353;
    end 
  end


  always @(posedge clk) begin
    if(N1351) begin
      T10[248] <= N1352;
    end 
  end


  always @(posedge clk) begin
    if(N1354) begin
      T10[247] <= N1356;
    end 
  end


  always @(posedge clk) begin
    if(N1354) begin
      T10[246] <= N1355;
    end 
  end


  always @(posedge clk) begin
    if(N1357) begin
      T10[245] <= N1359;
    end 
  end


  always @(posedge clk) begin
    if(N1357) begin
      T10[244] <= N1358;
    end 
  end


  always @(posedge clk) begin
    if(N1360) begin
      T10[243] <= N1362;
    end 
  end


  always @(posedge clk) begin
    if(N1360) begin
      T10[242] <= N1361;
    end 
  end


  always @(posedge clk) begin
    if(N1363) begin
      T10[241] <= N1365;
    end 
  end


  always @(posedge clk) begin
    if(N1363) begin
      T10[240] <= N1364;
    end 
  end


  always @(posedge clk) begin
    if(N1366) begin
      T10[239] <= N1368;
    end 
  end


  always @(posedge clk) begin
    if(N1366) begin
      T10[238] <= N1367;
    end 
  end


  always @(posedge clk) begin
    if(N1369) begin
      T10[237] <= N1371;
    end 
  end


  always @(posedge clk) begin
    if(N1369) begin
      T10[236] <= N1370;
    end 
  end


  always @(posedge clk) begin
    if(N1372) begin
      T10[235] <= N1374;
    end 
  end


  always @(posedge clk) begin
    if(N1372) begin
      T10[234] <= N1373;
    end 
  end


  always @(posedge clk) begin
    if(N1375) begin
      T10[233] <= N1377;
    end 
  end


  always @(posedge clk) begin
    if(N1375) begin
      T10[232] <= N1376;
    end 
  end


  always @(posedge clk) begin
    if(N1378) begin
      T10[231] <= N1380;
    end 
  end


  always @(posedge clk) begin
    if(N1378) begin
      T10[230] <= N1379;
    end 
  end


  always @(posedge clk) begin
    if(N1381) begin
      T10[229] <= N1383;
    end 
  end


  always @(posedge clk) begin
    if(N1381) begin
      T10[228] <= N1382;
    end 
  end


  always @(posedge clk) begin
    if(N1384) begin
      T10[227] <= N1386;
    end 
  end


  always @(posedge clk) begin
    if(N1384) begin
      T10[226] <= N1385;
    end 
  end


  always @(posedge clk) begin
    if(N1387) begin
      T10[225] <= N1389;
    end 
  end


  always @(posedge clk) begin
    if(N1387) begin
      T10[224] <= N1388;
    end 
  end


  always @(posedge clk) begin
    if(N1390) begin
      T10[223] <= N1392;
    end 
  end


  always @(posedge clk) begin
    if(N1390) begin
      T10[222] <= N1391;
    end 
  end


  always @(posedge clk) begin
    if(N1393) begin
      T10[221] <= N1395;
    end 
  end


  always @(posedge clk) begin
    if(N1393) begin
      T10[220] <= N1394;
    end 
  end


  always @(posedge clk) begin
    if(N1396) begin
      T10[219] <= N1398;
    end 
  end


  always @(posedge clk) begin
    if(N1396) begin
      T10[218] <= N1397;
    end 
  end


  always @(posedge clk) begin
    if(N1399) begin
      T10[217] <= N1401;
    end 
  end


  always @(posedge clk) begin
    if(N1399) begin
      T10[216] <= N1400;
    end 
  end


  always @(posedge clk) begin
    if(N1402) begin
      T10[215] <= N1404;
    end 
  end


  always @(posedge clk) begin
    if(N1402) begin
      T10[214] <= N1403;
    end 
  end


  always @(posedge clk) begin
    if(N1405) begin
      T10[213] <= N1407;
    end 
  end


  always @(posedge clk) begin
    if(N1405) begin
      T10[212] <= N1406;
    end 
  end


  always @(posedge clk) begin
    if(N1408) begin
      T10[211] <= N1410;
    end 
  end


  always @(posedge clk) begin
    if(N1408) begin
      T10[210] <= N1409;
    end 
  end


  always @(posedge clk) begin
    if(N1411) begin
      T10[209] <= N1413;
    end 
  end


  always @(posedge clk) begin
    if(N1411) begin
      T10[208] <= N1412;
    end 
  end


  always @(posedge clk) begin
    if(N1414) begin
      T10[207] <= N1416;
    end 
  end


  always @(posedge clk) begin
    if(N1414) begin
      T10[206] <= N1415;
    end 
  end


  always @(posedge clk) begin
    if(N1417) begin
      T10[205] <= N1419;
    end 
  end


  always @(posedge clk) begin
    if(N1417) begin
      T10[204] <= N1418;
    end 
  end


  always @(posedge clk) begin
    if(N1420) begin
      T10[203] <= N1422;
    end 
  end


  always @(posedge clk) begin
    if(N1420) begin
      T10[202] <= N1421;
    end 
  end


  always @(posedge clk) begin
    if(N1423) begin
      T10[201] <= N1425;
    end 
  end


  always @(posedge clk) begin
    if(N1423) begin
      T10[200] <= N1424;
    end 
  end


  always @(posedge clk) begin
    if(N1426) begin
      T10[199] <= N1428;
    end 
  end


  always @(posedge clk) begin
    if(N1426) begin
      T10[198] <= N1427;
    end 
  end


  always @(posedge clk) begin
    if(N1429) begin
      T10[197] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1429) begin
      T10[196] <= N1430;
    end 
  end


  always @(posedge clk) begin
    if(N1432) begin
      T10[195] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1432) begin
      T10[194] <= N1433;
    end 
  end


  always @(posedge clk) begin
    if(N1434) begin
      T10[193] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1434) begin
      T10[192] <= N1435;
    end 
  end


  always @(posedge clk) begin
    if(N1436) begin
      T10[191] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1436) begin
      T10[190] <= N1437;
    end 
  end


  always @(posedge clk) begin
    if(N1438) begin
      T10[189] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1438) begin
      T10[188] <= N1439;
    end 
  end


  always @(posedge clk) begin
    if(N1440) begin
      T10[187] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1440) begin
      T10[186] <= N1441;
    end 
  end


  always @(posedge clk) begin
    if(N1442) begin
      T10[185] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1442) begin
      T10[184] <= N1443;
    end 
  end


  always @(posedge clk) begin
    if(N1444) begin
      T10[183] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1444) begin
      T10[182] <= N1445;
    end 
  end


  always @(posedge clk) begin
    if(N1446) begin
      T10[181] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1446) begin
      T10[180] <= N1447;
    end 
  end


  always @(posedge clk) begin
    if(N1448) begin
      T10[179] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1448) begin
      T10[178] <= N1449;
    end 
  end


  always @(posedge clk) begin
    if(N1450) begin
      T10[177] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1450) begin
      T10[176] <= N1451;
    end 
  end


  always @(posedge clk) begin
    if(N1452) begin
      T10[175] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1452) begin
      T10[174] <= N1453;
    end 
  end


  always @(posedge clk) begin
    if(N1454) begin
      T10[173] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1454) begin
      T10[172] <= N1455;
    end 
  end


  always @(posedge clk) begin
    if(N1456) begin
      T10[171] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1456) begin
      T10[170] <= N1457;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T10[169] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1458) begin
      T10[168] <= N1459;
    end 
  end


  always @(posedge clk) begin
    if(N1460) begin
      T10[167] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1460) begin
      T10[166] <= N1461;
    end 
  end


  always @(posedge clk) begin
    if(N1462) begin
      T10[165] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1462) begin
      T10[164] <= N1463;
    end 
  end


  always @(posedge clk) begin
    if(N1464) begin
      T10[163] <= N1431;
    end 
  end


  always @(posedge clk) begin
    if(N1464) begin
      T10[162] <= N1465;
    end 
  end


  always @(posedge clk) begin
    if(N1466) begin
      T10[161] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1466) begin
      T10[160] <= N1467;
    end 
  end


  always @(posedge clk) begin
    if(N1469) begin
      T10[159] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1469) begin
      T10[158] <= N1470;
    end 
  end


  always @(posedge clk) begin
    if(N1471) begin
      T10[157] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1471) begin
      T10[156] <= N1472;
    end 
  end


  always @(posedge clk) begin
    if(N1473) begin
      T10[155] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1473) begin
      T10[154] <= N1474;
    end 
  end


  always @(posedge clk) begin
    if(N1475) begin
      T10[153] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1475) begin
      T10[152] <= N1476;
    end 
  end


  always @(posedge clk) begin
    if(N1477) begin
      T10[151] <= N1468;
    end 
  end


  always @(posedge clk) begin
    if(N1477) begin
      T10[150] <= N1478;
    end 
  end


  always @(posedge clk) begin
    if(N1479) begin
      T10[149] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1479) begin
      T10[148] <= N1480;
    end 
  end


  always @(posedge clk) begin
    if(N1482) begin
      T10[147] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1482) begin
      T10[146] <= N1483;
    end 
  end


  always @(posedge clk) begin
    if(N1484) begin
      T10[145] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1484) begin
      T10[144] <= N1485;
    end 
  end


  always @(posedge clk) begin
    if(N1486) begin
      T10[143] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1486) begin
      T10[142] <= N1487;
    end 
  end


  always @(posedge clk) begin
    if(N1488) begin
      T10[141] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1488) begin
      T10[140] <= N1489;
    end 
  end


  always @(posedge clk) begin
    if(N1490) begin
      T10[139] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1490) begin
      T10[138] <= N1491;
    end 
  end


  always @(posedge clk) begin
    if(N1492) begin
      T10[137] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1492) begin
      T10[136] <= N1493;
    end 
  end


  always @(posedge clk) begin
    if(N1494) begin
      T10[135] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1494) begin
      T10[134] <= N1495;
    end 
  end


  always @(posedge clk) begin
    if(N1496) begin
      T10[133] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1496) begin
      T10[132] <= N1497;
    end 
  end


  always @(posedge clk) begin
    if(N1498) begin
      T10[131] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1498) begin
      T10[130] <= N1499;
    end 
  end


  always @(posedge clk) begin
    if(N1500) begin
      T10[129] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1500) begin
      T10[128] <= N1501;
    end 
  end


  always @(posedge clk) begin
    if(N1502) begin
      T10[127] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1502) begin
      T10[126] <= N1503;
    end 
  end


  always @(posedge clk) begin
    if(N1504) begin
      T10[125] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1504) begin
      T10[124] <= N1505;
    end 
  end


  always @(posedge clk) begin
    if(N1506) begin
      T10[123] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1506) begin
      T10[122] <= N1507;
    end 
  end


  always @(posedge clk) begin
    if(N1508) begin
      T10[121] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1508) begin
      T10[120] <= N1509;
    end 
  end


  always @(posedge clk) begin
    if(N1510) begin
      T10[119] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1510) begin
      T10[118] <= N1511;
    end 
  end


  always @(posedge clk) begin
    if(N1512) begin
      T10[117] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1512) begin
      T10[116] <= N1513;
    end 
  end


  always @(posedge clk) begin
    if(N1514) begin
      T10[115] <= N1481;
    end 
  end


  always @(posedge clk) begin
    if(N1514) begin
      T10[114] <= N1515;
    end 
  end


  always @(posedge clk) begin
    if(N1516) begin
      T10[113] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1516) begin
      T10[112] <= N1517;
    end 
  end


  always @(posedge clk) begin
    if(N1519) begin
      T10[111] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1519) begin
      T10[110] <= N1520;
    end 
  end


  always @(posedge clk) begin
    if(N1521) begin
      T10[109] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1521) begin
      T10[108] <= N1522;
    end 
  end


  always @(posedge clk) begin
    if(N1523) begin
      T10[107] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1523) begin
      T10[106] <= N1524;
    end 
  end


  always @(posedge clk) begin
    if(N1525) begin
      T10[105] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1525) begin
      T10[104] <= N1526;
    end 
  end


  always @(posedge clk) begin
    if(N1527) begin
      T10[103] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1527) begin
      T10[102] <= N1528;
    end 
  end


  always @(posedge clk) begin
    if(N1529) begin
      T10[101] <= N1518;
    end 
  end


  always @(posedge clk) begin
    if(N1529) begin
      T10[100] <= N1530;
    end 
  end


  always @(posedge clk) begin
    if(N1531) begin
      T10[99] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1531) begin
      T10[98] <= N1532;
    end 
  end


  always @(posedge clk) begin
    if(N1534) begin
      T10[97] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1534) begin
      T10[96] <= N1535;
    end 
  end


  always @(posedge clk) begin
    if(N1536) begin
      T10[95] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1536) begin
      T10[94] <= N1537;
    end 
  end


  always @(posedge clk) begin
    if(N1538) begin
      T10[93] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1538) begin
      T10[92] <= N1539;
    end 
  end


  always @(posedge clk) begin
    if(N1540) begin
      T10[91] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1540) begin
      T10[90] <= N1541;
    end 
  end


  always @(posedge clk) begin
    if(N1542) begin
      T10[89] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1542) begin
      T10[88] <= N1543;
    end 
  end


  always @(posedge clk) begin
    if(N1544) begin
      T10[87] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1544) begin
      T10[86] <= N1545;
    end 
  end


  always @(posedge clk) begin
    if(N1546) begin
      T10[85] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1546) begin
      T10[84] <= N1547;
    end 
  end


  always @(posedge clk) begin
    if(N1548) begin
      T10[83] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1548) begin
      T10[82] <= N1549;
    end 
  end


  always @(posedge clk) begin
    if(N1550) begin
      T10[81] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1550) begin
      T10[80] <= N1551;
    end 
  end


  always @(posedge clk) begin
    if(N1552) begin
      T10[79] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1552) begin
      T10[78] <= N1553;
    end 
  end


  always @(posedge clk) begin
    if(N1554) begin
      T10[77] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1554) begin
      T10[76] <= N1555;
    end 
  end


  always @(posedge clk) begin
    if(N1556) begin
      T10[75] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1556) begin
      T10[74] <= N1557;
    end 
  end


  always @(posedge clk) begin
    if(N1558) begin
      T10[73] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1558) begin
      T10[72] <= N1559;
    end 
  end


  always @(posedge clk) begin
    if(N1560) begin
      T10[71] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1560) begin
      T10[70] <= N1561;
    end 
  end


  always @(posedge clk) begin
    if(N1562) begin
      T10[69] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1562) begin
      T10[68] <= N1563;
    end 
  end


  always @(posedge clk) begin
    if(N1564) begin
      T10[67] <= N1533;
    end 
  end


  always @(posedge clk) begin
    if(N1564) begin
      T10[66] <= N1565;
    end 
  end


  always @(posedge clk) begin
    if(N1566) begin
      T10[65] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1566) begin
      T10[64] <= N1567;
    end 
  end


  always @(posedge clk) begin
    if(N1569) begin
      T10[63] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1569) begin
      T10[62] <= N1570;
    end 
  end


  always @(posedge clk) begin
    if(N1571) begin
      T10[61] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1571) begin
      T10[60] <= N1572;
    end 
  end


  always @(posedge clk) begin
    if(N1573) begin
      T10[59] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1573) begin
      T10[58] <= N1574;
    end 
  end


  always @(posedge clk) begin
    if(N1575) begin
      T10[57] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1575) begin
      T10[56] <= N1576;
    end 
  end


  always @(posedge clk) begin
    if(N1577) begin
      T10[55] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1577) begin
      T10[54] <= N1578;
    end 
  end


  always @(posedge clk) begin
    if(N1579) begin
      T10[53] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1579) begin
      T10[52] <= N1580;
    end 
  end


  always @(posedge clk) begin
    if(N1581) begin
      T10[51] <= N1568;
    end 
  end


  always @(posedge clk) begin
    if(N1581) begin
      T10[50] <= N1582;
    end 
  end


  always @(posedge clk) begin
    if(N1583) begin
      T10[49] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1583) begin
      T10[48] <= N1584;
    end 
  end


  always @(posedge clk) begin
    if(N1586) begin
      T10[47] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1586) begin
      T10[46] <= N1587;
    end 
  end


  always @(posedge clk) begin
    if(N1588) begin
      T10[45] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1588) begin
      T10[44] <= N1589;
    end 
  end


  always @(posedge clk) begin
    if(N1590) begin
      T10[43] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1590) begin
      T10[42] <= N1591;
    end 
  end


  always @(posedge clk) begin
    if(N1592) begin
      T10[41] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1592) begin
      T10[40] <= N1593;
    end 
  end


  always @(posedge clk) begin
    if(N1594) begin
      T10[39] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1594) begin
      T10[38] <= N1595;
    end 
  end


  always @(posedge clk) begin
    if(N1596) begin
      T10[37] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1596) begin
      T10[36] <= N1597;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T10[35] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1598) begin
      T10[34] <= N1599;
    end 
  end


  always @(posedge clk) begin
    if(N1600) begin
      T10[33] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1600) begin
      T10[32] <= N1601;
    end 
  end


  always @(posedge clk) begin
    if(N1602) begin
      T10[31] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1602) begin
      T10[30] <= N1603;
    end 
  end


  always @(posedge clk) begin
    if(N1604) begin
      T10[29] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1604) begin
      T10[28] <= N1605;
    end 
  end


  always @(posedge clk) begin
    if(N1606) begin
      T10[27] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1606) begin
      T10[26] <= N1607;
    end 
  end


  always @(posedge clk) begin
    if(N1608) begin
      T10[25] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1608) begin
      T10[24] <= N1609;
    end 
  end


  always @(posedge clk) begin
    if(N1610) begin
      T10[23] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1610) begin
      T10[22] <= N1611;
    end 
  end


  always @(posedge clk) begin
    if(N1612) begin
      T10[21] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1612) begin
      T10[20] <= N1613;
    end 
  end


  always @(posedge clk) begin
    if(N1614) begin
      T10[19] <= N1585;
    end 
  end


  always @(posedge clk) begin
    if(N1614) begin
      T10[18] <= N1615;
    end 
  end


  always @(posedge clk) begin
    if(N1616) begin
      T10[17] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1616) begin
      T10[16] <= N1617;
    end 
  end


  always @(posedge clk) begin
    if(N1619) begin
      T10[15] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1619) begin
      T10[14] <= N1620;
    end 
  end


  always @(posedge clk) begin
    if(N1621) begin
      T10[13] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1621) begin
      T10[12] <= N1622;
    end 
  end


  always @(posedge clk) begin
    if(N1623) begin
      T10[11] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1623) begin
      T10[10] <= N1624;
    end 
  end


  always @(posedge clk) begin
    if(N1625) begin
      T10[9] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1625) begin
      T10[8] <= N1626;
    end 
  end


  always @(posedge clk) begin
    if(N1627) begin
      T10[7] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1627) begin
      T10[6] <= N1628;
    end 
  end


  always @(posedge clk) begin
    if(N1629) begin
      T10[5] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1629) begin
      T10[4] <= N1630;
    end 
  end


  always @(posedge clk) begin
    if(N1631) begin
      T10[3] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1631) begin
      T10[2] <= N1632;
    end 
  end


  always @(posedge clk) begin
    if(N1633) begin
      T10[1] <= N1618;
    end 
  end


  always @(posedge clk) begin
    if(N1633) begin
      T10[0] <= N1634;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[6] <= N1645;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[5] <= N1644;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[4] <= N1643;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[3] <= N1642;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[2] <= N1641;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[1] <= N1640;
    end 
  end


  always @(posedge clk) begin
    if(N1638) begin
      io_resp_bits_bht_history[0] <= N1639;
    end 
  end


  always @(posedge clk) begin
    if(T166) begin
      isJump_61 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R164 <= io_btb_update_bits_isJump;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[5] <= N1654;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[4] <= N1653;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[3] <= N1652;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[2] <= N1651;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[1] <= N1650;
    end 
  end


  always @(posedge clk) begin
    if(N1648) begin
      nextRepl[0] <= N1649;
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[5] <= io_btb_update_bits_prediction_bits_entry[5];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[4] <= io_btb_update_bits_prediction_bits_entry[4];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[3] <= io_btb_update_bits_prediction_bits_entry[3];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[2] <= io_btb_update_bits_prediction_bits_entry[2];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[1] <= io_btb_update_bits_prediction_bits_entry[1];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R177[0] <= io_btb_update_bits_prediction_bits_entry[0];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      updateHit <= io_btb_update_bits_prediction_valid;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[5] <= N1664;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[4] <= N1663;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[3] <= N1662;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[2] <= N1661;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[1] <= N1660;
    end 
  end


  always @(posedge clk) begin
    if(N1658) begin
      pageValid[0] <= N1659;
    end 
  end


  always @(posedge clk) begin
    if(N1667) begin
      R198[2] <= N1670;
    end 
  end


  always @(posedge clk) begin
    if(N1667) begin
      R198[1] <= N1669;
    end 
  end


  always @(posedge clk) begin
    if(N1667) begin
      R198[0] <= N1668;
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[26] <= io_btb_update_bits_pc[38];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[25] <= io_btb_update_bits_pc[37];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[24] <= io_btb_update_bits_pc[36];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[23] <= io_btb_update_bits_pc[35];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[22] <= io_btb_update_bits_pc[34];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[21] <= io_btb_update_bits_pc[33];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[20] <= io_btb_update_bits_pc[32];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[19] <= io_btb_update_bits_pc[31];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[18] <= io_btb_update_bits_pc[30];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[17] <= io_btb_update_bits_pc[29];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[16] <= io_btb_update_bits_pc[28];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[15] <= io_btb_update_bits_pc[27];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[14] <= io_btb_update_bits_pc[26];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[13] <= io_btb_update_bits_pc[25];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[12] <= io_btb_update_bits_pc[24];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[11] <= io_btb_update_bits_pc[23];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[10] <= io_btb_update_bits_pc[22];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[9] <= io_btb_update_bits_pc[21];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[8] <= io_btb_update_bits_pc[20];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[7] <= io_btb_update_bits_pc[19];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[6] <= io_btb_update_bits_pc[18];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[5] <= io_btb_update_bits_pc[17];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[4] <= io_btb_update_bits_pc[16];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[3] <= io_btb_update_bits_pc[15];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[2] <= io_btb_update_bits_pc[14];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[1] <= io_btb_update_bits_pc[13];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T209[0] <= io_btb_update_bits_pc[12];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[11] <= io_btb_update_bits_pc[11];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[10] <= io_btb_update_bits_pc[10];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[9] <= io_btb_update_bits_pc[9];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[8] <= io_btb_update_bits_pc[8];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[7] <= io_btb_update_bits_pc[7];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[6] <= io_btb_update_bits_pc[6];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[5] <= io_btb_update_bits_pc[5];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[4] <= io_btb_update_bits_pc[4];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[3] <= io_btb_update_bits_pc[3];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[2] <= io_btb_update_bits_pc[2];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[1] <= io_btb_update_bits_pc[1];
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      T2434[0] <= io_btb_update_bits_pc[0];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[26] <= T214[26];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[25] <= T214[25];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[24] <= T214[24];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[23] <= T214[23];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[22] <= T214[22];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[21] <= T214[21];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[20] <= T214[20];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[19] <= T214[19];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[18] <= T214[18];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[17] <= T214[17];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[16] <= T214[16];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[15] <= T214[15];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[14] <= T214[14];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[13] <= T214[13];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[12] <= T214[12];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[11] <= T214[11];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[10] <= T214[10];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[9] <= T214[9];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[8] <= T214[8];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[7] <= T214[7];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[6] <= T214[6];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[5] <= T214[5];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[4] <= T214[4];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[3] <= T214[3];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[2] <= T214[2];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[1] <= T214[1];
    end 
  end


  always @(posedge clk) begin
    if(T219) begin
      T258[0] <= T214[0];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[26] <= T232[26];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[25] <= T232[25];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[24] <= T232[24];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[23] <= T232[23];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[22] <= T232[22];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[21] <= T232[21];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[20] <= T232[20];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[19] <= T232[19];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[18] <= T232[18];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[17] <= T232[17];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[16] <= T232[16];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[15] <= T232[15];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[14] <= T232[14];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[13] <= T232[13];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[12] <= T232[12];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[11] <= T232[11];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[10] <= T232[10];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[9] <= T232[9];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[8] <= T232[8];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[7] <= T232[7];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[6] <= T232[6];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[5] <= T232[5];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[4] <= T232[4];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[3] <= T232[3];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[2] <= T232[2];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[1] <= T232[1];
    end 
  end


  always @(posedge clk) begin
    if(T235) begin
      T256[0] <= T232[0];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[26] <= T214[26];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[25] <= T214[25];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[24] <= T214[24];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[23] <= T214[23];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[22] <= T214[22];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[21] <= T214[21];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[20] <= T214[20];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[19] <= T214[19];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[18] <= T214[18];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[17] <= T214[17];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[16] <= T214[16];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[15] <= T214[15];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[14] <= T214[14];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[13] <= T214[13];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[12] <= T214[12];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[11] <= T214[11];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[10] <= T214[10];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[9] <= T214[9];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[8] <= T214[8];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[7] <= T214[7];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[6] <= T214[6];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[5] <= T214[5];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[4] <= T214[4];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[3] <= T214[3];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[2] <= T214[2];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[1] <= T214[1];
    end 
  end


  always @(posedge clk) begin
    if(T224) begin
      T254[0] <= T214[0];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[26] <= T232[26];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[25] <= T232[25];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[24] <= T232[24];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[23] <= T232[23];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[22] <= T232[22];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[21] <= T232[21];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[20] <= T232[20];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[19] <= T232[19];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[18] <= T232[18];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[17] <= T232[17];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[16] <= T232[16];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[15] <= T232[15];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[14] <= T232[14];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[13] <= T232[13];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[12] <= T232[12];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[11] <= T232[11];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[10] <= T232[10];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[9] <= T232[9];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[8] <= T232[8];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[7] <= T232[7];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[6] <= T232[6];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[5] <= T232[5];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[4] <= T232[4];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[3] <= T232[3];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[2] <= T232[2];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[1] <= T232[1];
    end 
  end


  always @(posedge clk) begin
    if(T240) begin
      T250[0] <= T232[0];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[26] <= T214[26];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[25] <= T214[25];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[24] <= T214[24];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[23] <= T214[23];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[22] <= T214[22];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[21] <= T214[21];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[20] <= T214[20];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[19] <= T214[19];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[18] <= T214[18];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[17] <= T214[17];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[16] <= T214[16];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[15] <= T214[15];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[14] <= T214[14];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[13] <= T214[13];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[12] <= T214[12];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[11] <= T214[11];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[10] <= T214[10];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[9] <= T214[9];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[8] <= T214[8];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[7] <= T214[7];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[6] <= T214[6];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[5] <= T214[5];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[4] <= T214[4];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[3] <= T214[3];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[2] <= T214[2];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[1] <= T214[1];
    end 
  end


  always @(posedge clk) begin
    if(T228) begin
      T248[0] <= T214[0];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[26] <= T232[26];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[25] <= T232[25];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[24] <= T232[24];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[23] <= T232[23];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[22] <= T232[22];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[21] <= T232[21];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[20] <= T232[20];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[19] <= T232[19];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[18] <= T232[18];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[17] <= T232[17];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[16] <= T232[16];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[15] <= T232[15];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[14] <= T232[14];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[13] <= T232[13];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[12] <= T232[12];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[11] <= T232[11];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[10] <= T232[10];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[9] <= T232[9];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[8] <= T232[8];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[7] <= T232[7];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[6] <= T232[6];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[5] <= T232[5];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[4] <= T232[4];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[3] <= T232[3];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[2] <= T232[2];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[1] <= T232[1];
    end 
  end


  always @(posedge clk) begin
    if(T244) begin
      T212[0] <= T232[0];
    end 
  end


  always @(posedge clk) begin
    if(N1795) begin
      T588[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1795) begin
      T588[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1795) begin
      T588[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1794) begin
      T584[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1794) begin
      T584[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1794) begin
      T584[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1793) begin
      T580[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1793) begin
      T580[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1793) begin
      T580[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1792) begin
      T574[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1792) begin
      T574[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1792) begin
      T574[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1791) begin
      T570[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1791) begin
      T570[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1791) begin
      T570[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1790) begin
      T565[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1790) begin
      T565[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1790) begin
      T565[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1789) begin
      T561[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1789) begin
      T561[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1789) begin
      T561[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1788) begin
      T554[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1788) begin
      T554[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1788) begin
      T554[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1787) begin
      T550[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1787) begin
      T550[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1787) begin
      T550[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1786) begin
      T545[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1786) begin
      T545[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1786) begin
      T545[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1785) begin
      T541[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1785) begin
      T541[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1785) begin
      T541[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1784) begin
      T535[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1784) begin
      T535[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1784) begin
      T535[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1783) begin
      T531[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1783) begin
      T531[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1783) begin
      T531[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1782) begin
      T526[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1782) begin
      T526[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1782) begin
      T526[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1781) begin
      T522[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1781) begin
      T522[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1781) begin
      T522[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1780) begin
      T514[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1780) begin
      T514[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1780) begin
      T514[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1779) begin
      T510[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1779) begin
      T510[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1779) begin
      T510[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1778) begin
      T505[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1778) begin
      T505[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1778) begin
      T505[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1777) begin
      T501[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1777) begin
      T501[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1777) begin
      T501[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1776) begin
      T495[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1776) begin
      T495[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1776) begin
      T495[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1775) begin
      T491[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1775) begin
      T491[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1775) begin
      T491[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1774) begin
      T486[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1774) begin
      T486[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1774) begin
      T486[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1773) begin
      T482[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1773) begin
      T482[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1773) begin
      T482[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1772) begin
      T475[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1772) begin
      T475[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1772) begin
      T475[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1771) begin
      T471[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1771) begin
      T471[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1771) begin
      T471[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1770) begin
      T466[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1770) begin
      T466[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1770) begin
      T466[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1769) begin
      T462[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1769) begin
      T462[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1769) begin
      T462[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1768) begin
      T456[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1768) begin
      T456[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1768) begin
      T456[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1767) begin
      T452[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1767) begin
      T452[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1767) begin
      T452[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1766) begin
      T447[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1766) begin
      T447[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1766) begin
      T447[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1765) begin
      T443[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1765) begin
      T443[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1765) begin
      T443[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1764) begin
      T434[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1764) begin
      T434[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1764) begin
      T434[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1763) begin
      T430[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1763) begin
      T430[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1763) begin
      T430[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1762) begin
      T426[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1762) begin
      T426[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1762) begin
      T426[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1761) begin
      T420[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1761) begin
      T420[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1761) begin
      T420[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1760) begin
      T416[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1760) begin
      T416[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1760) begin
      T416[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1759) begin
      T411[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1759) begin
      T411[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1759) begin
      T411[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1758) begin
      T407[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1758) begin
      T407[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1758) begin
      T407[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1757) begin
      T400[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1757) begin
      T400[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1757) begin
      T400[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1756) begin
      T396[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1756) begin
      T396[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1756) begin
      T396[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1755) begin
      T391[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1755) begin
      T391[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1755) begin
      T391[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1754) begin
      T387[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1754) begin
      T387[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1754) begin
      T387[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1753) begin
      T381[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1753) begin
      T381[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1753) begin
      T381[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1752) begin
      T377[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1752) begin
      T377[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1752) begin
      T377[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1751) begin
      T372[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1751) begin
      T372[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1751) begin
      T372[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1750) begin
      T368[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1750) begin
      T368[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1750) begin
      T368[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T360[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T360[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1749) begin
      T360[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1748) begin
      T356[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1748) begin
      T356[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1748) begin
      T356[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1747) begin
      T351[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1747) begin
      T351[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1747) begin
      T351[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1746) begin
      T347[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1746) begin
      T347[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1746) begin
      T347[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1745) begin
      T341[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1745) begin
      T341[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1745) begin
      T341[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1744) begin
      T337[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1744) begin
      T337[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1744) begin
      T337[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1743) begin
      T332[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1743) begin
      T332[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1743) begin
      T332[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1742) begin
      T328[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1742) begin
      T328[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1742) begin
      T328[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1741) begin
      T321[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1741) begin
      T321[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1741) begin
      T321[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1740) begin
      T317[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1740) begin
      T317[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1740) begin
      T317[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T312[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T312[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1739) begin
      T312[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1738) begin
      T308[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1738) begin
      T308[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1738) begin
      T308[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1737) begin
      T302[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1737) begin
      T302[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1737) begin
      T302[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1736) begin
      T298[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1736) begin
      T298[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1736) begin
      T298[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1735) begin
      T293[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1735) begin
      T293[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1735) begin
      T293[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1734) begin
      T286[2] <= N2328;
    end 
  end


  always @(posedge clk) begin
    if(N1734) begin
      T286[1] <= N2329;
    end 
  end


  always @(posedge clk) begin
    if(N1734) begin
      T286[0] <= T2423[0];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1920) begin
      T779[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1919) begin
      T777[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1918) begin
      T775[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1917) begin
      T771[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1916) begin
      T769[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1915) begin
      T766[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1914) begin
      T764[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1913) begin
      T759[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1912) begin
      T757[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1911) begin
      T754[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1910) begin
      T752[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1909) begin
      T748[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1908) begin
      T746[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1907) begin
      T743[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1906) begin
      T741[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1905) begin
      T735[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1904) begin
      T733[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1903) begin
      T730[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1902) begin
      T728[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1901) begin
      T724[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1900) begin
      T722[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1899) begin
      T719[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1898) begin
      T717[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1897) begin
      T712[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1896) begin
      T710[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1895) begin
      T707[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1894) begin
      T705[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1893) begin
      T701[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1892) begin
      T699[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1891) begin
      T696[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1890) begin
      T694[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1889) begin
      T687[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1888) begin
      T685[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1887) begin
      T683[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1886) begin
      T679[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1885) begin
      T677[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1884) begin
      T674[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1883) begin
      T672[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1882) begin
      T667[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1881) begin
      T665[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1880) begin
      T662[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1879) begin
      T660[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1878) begin
      T656[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1877) begin
      T654[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1876) begin
      T651[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1875) begin
      T649[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1874) begin
      T643[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1873) begin
      T641[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1872) begin
      T638[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1871) begin
      T636[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1870) begin
      T632[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1869) begin
      T630[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1868) begin
      T627[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1867) begin
      T625[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1866) begin
      T620[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1865) begin
      T618[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1864) begin
      T615[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1863) begin
      T613[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1862) begin
      T609[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1861) begin
      T607[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1860) begin
      T604[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[11] <= T2434[11];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[10] <= T2434[10];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[9] <= T2434[9];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[8] <= T2434[8];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[7] <= T2434[7];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[6] <= T2434[6];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[5] <= T2434[5];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[4] <= T2434[4];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[3] <= T2434[3];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[2] <= T2434[2];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[1] <= T2434[1];
    end 
  end


  always @(posedge clk) begin
    if(N1859) begin
      T599[0] <= T2434[0];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[61] <= T2435[61];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[60] <= T2435[60];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[59] <= T2435[59];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[58] <= T2435[58];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[57] <= T2435[57];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[56] <= T2435[56];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[55] <= T2435[55];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[54] <= T2435[54];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[53] <= T2435[53];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[52] <= T2435[52];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[51] <= T2435[51];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[50] <= T2435[50];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[49] <= T2435[49];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[48] <= T2435[48];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[47] <= T2435[47];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[46] <= T2435[46];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[45] <= T2435[45];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[44] <= T2435[44];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[43] <= T2435[43];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[42] <= T2435[42];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[41] <= T2435[41];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[40] <= T2435[40];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[39] <= T2435[39];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[38] <= T2435[38];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[37] <= T2435[37];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[36] <= T2435[36];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[35] <= T2435[35];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[34] <= T2435[34];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[33] <= T2435[33];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[32] <= T2435[32];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[31] <= T2435[31];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[30] <= T2435[30];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[29] <= T2435[29];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[28] <= T2435[28];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[27] <= T2435[27];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[26] <= T2435[26];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[25] <= T2435[25];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[24] <= T2435[24];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[23] <= T2435[23];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[22] <= T2435[22];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[21] <= T2435[21];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[20] <= T2435[20];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[19] <= T2435[19];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[18] <= T2435[18];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[17] <= T2435[17];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[16] <= T2435[16];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[15] <= T2435[15];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[14] <= T2435[14];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[13] <= T2435[13];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[12] <= T2435[12];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[11] <= T2435[11];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[10] <= T2435[10];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[9] <= T2435[9];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[8] <= T2435[8];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[7] <= T2435[7];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[6] <= T2435[6];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[5] <= T2435[5];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[4] <= T2435[4];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[3] <= T2435[3];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[2] <= T2435[2];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[1] <= T2435[1];
    end 
  end


  always @(posedge clk) begin
    if(N2327) begin
      T2437[0] <= T2435[0];
    end 
  end


  always @(posedge clk) begin
    if(N2045) begin
      T1161[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2045) begin
      T1161[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2045) begin
      T1161[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2044) begin
      T1156[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2044) begin
      T1156[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2044) begin
      T1156[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2043) begin
      T1151[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2043) begin
      T1151[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2043) begin
      T1151[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2042) begin
      T1144[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2042) begin
      T1144[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2042) begin
      T1144[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2041) begin
      T1139[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2041) begin
      T1139[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2041) begin
      T1139[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2040) begin
      T1133[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2040) begin
      T1133[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2040) begin
      T1133[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2039) begin
      T1128[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2039) begin
      T1128[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2039) begin
      T1128[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2038) begin
      T1120[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2038) begin
      T1120[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2038) begin
      T1120[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2037) begin
      T1115[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2037) begin
      T1115[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2037) begin
      T1115[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2036) begin
      T1109[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2036) begin
      T1109[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2036) begin
      T1109[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2035) begin
      T1104[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2035) begin
      T1104[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2035) begin
      T1104[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2034) begin
      T1097[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2034) begin
      T1097[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2034) begin
      T1097[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2033) begin
      T1092[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2033) begin
      T1092[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2033) begin
      T1092[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      T1086[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      T1086[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2032) begin
      T1086[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2031) begin
      T1081[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2031) begin
      T1081[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2031) begin
      T1081[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2030) begin
      T1072[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2030) begin
      T1072[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2030) begin
      T1072[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2029) begin
      T1067[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2029) begin
      T1067[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2029) begin
      T1067[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2028) begin
      T1061[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2028) begin
      T1061[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2028) begin
      T1061[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2027) begin
      T1056[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2027) begin
      T1056[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2027) begin
      T1056[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2026) begin
      T1049[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2026) begin
      T1049[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2026) begin
      T1049[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2025) begin
      T1044[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2025) begin
      T1044[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2025) begin
      T1044[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2024) begin
      T1038[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2024) begin
      T1038[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2024) begin
      T1038[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2023) begin
      T1033[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2023) begin
      T1033[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2023) begin
      T1033[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2022) begin
      T1025[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2022) begin
      T1025[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2022) begin
      T1025[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2021) begin
      T1020[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2021) begin
      T1020[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2021) begin
      T1020[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2020) begin
      T1014[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2020) begin
      T1014[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2020) begin
      T1014[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2019) begin
      T1009[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2019) begin
      T1009[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2019) begin
      T1009[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2018) begin
      T1002[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2018) begin
      T1002[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2018) begin
      T1002[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2017) begin
      T997[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2017) begin
      T997[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2017) begin
      T997[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2016) begin
      T991[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2016) begin
      T991[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2016) begin
      T991[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2015) begin
      T986[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2015) begin
      T986[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2015) begin
      T986[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2014) begin
      T976[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2014) begin
      T976[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2014) begin
      T976[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2013) begin
      T971[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2013) begin
      T971[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2013) begin
      T971[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2012) begin
      T966[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2012) begin
      T966[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2012) begin
      T966[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2011) begin
      T959[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2011) begin
      T959[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2011) begin
      T959[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2010) begin
      T954[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2010) begin
      T954[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2010) begin
      T954[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2009) begin
      T948[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2009) begin
      T948[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2009) begin
      T948[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2008) begin
      T943[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2008) begin
      T943[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2008) begin
      T943[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2007) begin
      T935[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2007) begin
      T935[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2007) begin
      T935[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2006) begin
      T930[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2006) begin
      T930[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2006) begin
      T930[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2005) begin
      T924[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2005) begin
      T924[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2005) begin
      T924[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2004) begin
      T919[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2004) begin
      T919[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2004) begin
      T919[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2003) begin
      T912[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2003) begin
      T912[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2003) begin
      T912[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2002) begin
      T907[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2002) begin
      T907[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2002) begin
      T907[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2001) begin
      T901[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2001) begin
      T901[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2001) begin
      T901[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N2000) begin
      T896[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N2000) begin
      T896[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N2000) begin
      T896[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1999) begin
      T887[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1999) begin
      T887[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1999) begin
      T887[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1998) begin
      T882[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1998) begin
      T882[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1998) begin
      T882[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1997) begin
      T876[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1997) begin
      T876[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1997) begin
      T876[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1996) begin
      T871[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1996) begin
      T871[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1996) begin
      T871[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1995) begin
      T864[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1995) begin
      T864[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1995) begin
      T864[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1994) begin
      T859[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1994) begin
      T859[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1994) begin
      T859[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1993) begin
      T853[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1993) begin
      T853[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1993) begin
      T853[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1992) begin
      T848[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1992) begin
      T848[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1992) begin
      T848[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1991) begin
      T840[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1991) begin
      T840[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1991) begin
      T840[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1990) begin
      T835[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1990) begin
      T835[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1990) begin
      T835[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1989) begin
      T829[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1989) begin
      T829[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1989) begin
      T829[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1988) begin
      T824[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1988) begin
      T824[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1988) begin
      T824[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1987) begin
      T817[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1987) begin
      T817[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1987) begin
      T817[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      T812[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      T812[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1986) begin
      T812[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1985) begin
      T806[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1985) begin
      T806[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1985) begin
      T806[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(N1984) begin
      T797[2] <= N2330;
    end 
  end


  always @(posedge clk) begin
    if(N1984) begin
      T797[1] <= N2331;
    end 
  end


  always @(posedge clk) begin
    if(N1984) begin
      T797[0] <= T2439[0];
    end 
  end


  always @(posedge clk) begin
    if(T1165) begin
      isJump_60 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1171) begin
      isJump_59 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1177) begin
      isJump_58 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1183) begin
      isJump_57 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1189) begin
      isJump_56 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1195) begin
      isJump_55 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1201) begin
      isJump_54 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1207) begin
      isJump_53 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1213) begin
      isJump_52 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1219) begin
      isJump_51 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1225) begin
      isJump_50 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1231) begin
      isJump_49 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1237) begin
      isJump_48 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1243) begin
      isJump_47 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1249) begin
      isJump_46 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1255) begin
      isJump_45 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1261) begin
      isJump_44 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1267) begin
      isJump_43 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1273) begin
      isJump_42 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1279) begin
      isJump_41 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1285) begin
      isJump_40 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1291) begin
      isJump_39 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1297) begin
      isJump_38 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1303) begin
      isJump_37 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1309) begin
      isJump_36 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1315) begin
      isJump_35 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1321) begin
      isJump_34 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1327) begin
      isJump_33 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1333) begin
      isJump_32 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1339) begin
      isJump_31 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1345) begin
      isJump_30 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1351) begin
      isJump_29 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1357) begin
      isJump_28 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1363) begin
      isJump_27 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1369) begin
      isJump_26 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1375) begin
      isJump_25 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1381) begin
      isJump_24 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1387) begin
      isJump_23 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1393) begin
      isJump_22 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1399) begin
      isJump_21 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1405) begin
      isJump_20 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1411) begin
      isJump_19 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1417) begin
      isJump_18 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1423) begin
      isJump_17 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1429) begin
      isJump_16 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1435) begin
      isJump_15 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1441) begin
      isJump_14 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1447) begin
      isJump_13 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1453) begin
      isJump_12 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1459) begin
      isJump_11 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1465) begin
      isJump_10 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1471) begin
      isJump_9 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1477) begin
      isJump_8 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1483) begin
      isJump_7 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1489) begin
      isJump_6 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1495) begin
      isJump_5 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1501) begin
      isJump_4 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1507) begin
      isJump_3 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1513) begin
      isJump_2 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1519) begin
      isJump_1 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(T1524) begin
      isJump_0 <= R164;
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2170) begin
      T1539[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2169) begin
      T1546[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2168) begin
      T1550[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2167) begin
      T1554[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2166) begin
      T1558[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2165) begin
      T1562[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2164) begin
      T1566[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2163) begin
      T1570[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2162) begin
      T1574[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2161) begin
      T1578[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2160) begin
      T1582[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2159) begin
      T1586[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2158) begin
      T1590[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2157) begin
      T1594[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2156) begin
      T1598[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2155) begin
      T1602[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2154) begin
      T1606[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2153) begin
      T1610[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2152) begin
      T1614[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2151) begin
      T1618[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2150) begin
      T1622[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2149) begin
      T1626[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2148) begin
      T1630[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2147) begin
      T1634[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2146) begin
      T1638[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2145) begin
      T1642[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2144) begin
      T1646[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2143) begin
      T1650[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2142) begin
      T1654[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2141) begin
      T1658[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2140) begin
      T1662[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2139) begin
      T1666[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2138) begin
      T1670[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2137) begin
      T1674[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2136) begin
      T1678[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2135) begin
      T1682[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2134) begin
      T1686[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2133) begin
      T1690[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2132) begin
      T1694[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2131) begin
      T1698[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2130) begin
      T1702[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2129) begin
      T1706[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2128) begin
      T1710[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2127) begin
      T1714[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2126) begin
      T1718[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2125) begin
      T1722[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2124) begin
      T1726[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2123) begin
      T1730[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2122) begin
      T1734[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2121) begin
      T1738[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2120) begin
      T1742[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2119) begin
      T1746[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2118) begin
      T1750[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2117) begin
      T1754[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2116) begin
      T1758[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2115) begin
      T1762[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2114) begin
      T1766[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2113) begin
      T1770[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2112) begin
      T1774[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2111) begin
      T1778[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2110) begin
      T1782[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[11] <= io_req_bits_addr[11];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[10] <= io_req_bits_addr[10];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[9] <= io_req_bits_addr[9];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[8] <= io_req_bits_addr[8];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[7] <= io_req_bits_addr[7];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[6] <= io_req_bits_addr[6];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[5] <= io_req_bits_addr[5];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[4] <= io_req_bits_addr[4];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[3] <= io_req_bits_addr[3];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[2] <= io_req_bits_addr[2];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[1] <= io_req_bits_addr[1];
    end 
  end


  always @(posedge clk) begin
    if(N2109) begin
      T1785[0] <= io_req_bits_addr[0];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[38] <= io_ras_update_bits_returnAddr[38];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[37] <= io_ras_update_bits_returnAddr[37];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[36] <= io_ras_update_bits_returnAddr[36];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[35] <= io_ras_update_bits_returnAddr[35];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[34] <= io_ras_update_bits_returnAddr[34];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[33] <= io_ras_update_bits_returnAddr[33];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[32] <= io_ras_update_bits_returnAddr[32];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[31] <= io_ras_update_bits_returnAddr[31];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[30] <= io_ras_update_bits_returnAddr[30];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[29] <= io_ras_update_bits_returnAddr[29];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[28] <= io_ras_update_bits_returnAddr[28];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[27] <= io_ras_update_bits_returnAddr[27];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[26] <= io_ras_update_bits_returnAddr[26];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[25] <= io_ras_update_bits_returnAddr[25];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[24] <= io_ras_update_bits_returnAddr[24];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[23] <= io_ras_update_bits_returnAddr[23];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[22] <= io_ras_update_bits_returnAddr[22];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[21] <= io_ras_update_bits_returnAddr[21];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[20] <= io_ras_update_bits_returnAddr[20];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[19] <= io_ras_update_bits_returnAddr[19];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[18] <= io_ras_update_bits_returnAddr[18];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[17] <= io_ras_update_bits_returnAddr[17];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[16] <= io_ras_update_bits_returnAddr[16];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[15] <= io_ras_update_bits_returnAddr[15];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[14] <= io_ras_update_bits_returnAddr[14];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[13] <= io_ras_update_bits_returnAddr[13];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[12] <= io_ras_update_bits_returnAddr[12];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[11] <= io_ras_update_bits_returnAddr[11];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[10] <= io_ras_update_bits_returnAddr[10];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[9] <= io_ras_update_bits_returnAddr[9];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[8] <= io_ras_update_bits_returnAddr[8];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[7] <= io_ras_update_bits_returnAddr[7];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[6] <= io_ras_update_bits_returnAddr[6];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[5] <= io_ras_update_bits_returnAddr[5];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[4] <= io_ras_update_bits_returnAddr[4];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[3] <= io_ras_update_bits_returnAddr[3];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[2] <= io_ras_update_bits_returnAddr[2];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[1] <= io_ras_update_bits_returnAddr[1];
    end 
  end


  always @(posedge clk) begin
    if(T1998) begin
      R1996[0] <= io_ras_update_bits_returnAddr[0];
    end 
  end


  always @(posedge clk) begin
    if(N2174) begin
      T2027 <= N2175;
    end 
  end


  always @(posedge clk) begin
    if(N2179) begin
      R2010[1] <= N2181;
    end 
  end


  always @(posedge clk) begin
    if(N2179) begin
      R2010[0] <= N2180;
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[38] <= io_ras_update_bits_returnAddr[38];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[37] <= io_ras_update_bits_returnAddr[37];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[36] <= io_ras_update_bits_returnAddr[36];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[35] <= io_ras_update_bits_returnAddr[35];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[34] <= io_ras_update_bits_returnAddr[34];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[33] <= io_ras_update_bits_returnAddr[33];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[32] <= io_ras_update_bits_returnAddr[32];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[31] <= io_ras_update_bits_returnAddr[31];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[30] <= io_ras_update_bits_returnAddr[30];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[29] <= io_ras_update_bits_returnAddr[29];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[28] <= io_ras_update_bits_returnAddr[28];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[27] <= io_ras_update_bits_returnAddr[27];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[26] <= io_ras_update_bits_returnAddr[26];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[25] <= io_ras_update_bits_returnAddr[25];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[24] <= io_ras_update_bits_returnAddr[24];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[23] <= io_ras_update_bits_returnAddr[23];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[22] <= io_ras_update_bits_returnAddr[22];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[21] <= io_ras_update_bits_returnAddr[21];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[20] <= io_ras_update_bits_returnAddr[20];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[19] <= io_ras_update_bits_returnAddr[19];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[18] <= io_ras_update_bits_returnAddr[18];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[17] <= io_ras_update_bits_returnAddr[17];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[16] <= io_ras_update_bits_returnAddr[16];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[15] <= io_ras_update_bits_returnAddr[15];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[14] <= io_ras_update_bits_returnAddr[14];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[13] <= io_ras_update_bits_returnAddr[13];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[12] <= io_ras_update_bits_returnAddr[12];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[11] <= io_ras_update_bits_returnAddr[11];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[10] <= io_ras_update_bits_returnAddr[10];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[9] <= io_ras_update_bits_returnAddr[9];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[8] <= io_ras_update_bits_returnAddr[8];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[7] <= io_ras_update_bits_returnAddr[7];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[6] <= io_ras_update_bits_returnAddr[6];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[5] <= io_ras_update_bits_returnAddr[5];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[4] <= io_ras_update_bits_returnAddr[4];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[3] <= io_ras_update_bits_returnAddr[3];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[2] <= io_ras_update_bits_returnAddr[2];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[1] <= io_ras_update_bits_returnAddr[1];
    end 
  end


  always @(posedge clk) begin
    if(T2025) begin
      R2023[0] <= io_ras_update_bits_returnAddr[0];
    end 
  end


  always @(posedge clk) begin
    if(T2034) begin
      useRAS_61 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(io_btb_update_valid) begin
      R2032 <= io_btb_update_bits_isReturn;
    end 
  end


  always @(posedge clk) begin
    if(T2042) begin
      useRAS_60 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2048) begin
      useRAS_59 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2054) begin
      useRAS_58 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2060) begin
      useRAS_57 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2066) begin
      useRAS_56 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2072) begin
      useRAS_55 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2078) begin
      useRAS_54 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2084) begin
      useRAS_53 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2090) begin
      useRAS_52 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2096) begin
      useRAS_51 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2102) begin
      useRAS_50 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2108) begin
      useRAS_49 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2114) begin
      useRAS_48 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2120) begin
      useRAS_47 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2126) begin
      useRAS_46 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2132) begin
      useRAS_45 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2138) begin
      useRAS_44 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2144) begin
      useRAS_43 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2150) begin
      useRAS_42 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2156) begin
      useRAS_41 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2162) begin
      useRAS_40 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2168) begin
      useRAS_39 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2174) begin
      useRAS_38 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2180) begin
      useRAS_37 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2186) begin
      useRAS_36 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2192) begin
      useRAS_35 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2198) begin
      useRAS_34 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2204) begin
      useRAS_33 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2210) begin
      useRAS_32 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2216) begin
      useRAS_31 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2222) begin
      useRAS_30 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2228) begin
      useRAS_29 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2234) begin
      useRAS_28 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2240) begin
      useRAS_27 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2246) begin
      useRAS_26 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2252) begin
      useRAS_25 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2258) begin
      useRAS_24 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2264) begin
      useRAS_23 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2270) begin
      useRAS_22 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2276) begin
      useRAS_21 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2282) begin
      useRAS_20 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2288) begin
      useRAS_19 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2294) begin
      useRAS_18 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2300) begin
      useRAS_17 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2306) begin
      useRAS_16 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2312) begin
      useRAS_15 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2318) begin
      useRAS_14 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2324) begin
      useRAS_13 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2330) begin
      useRAS_12 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2336) begin
      useRAS_11 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2342) begin
      useRAS_10 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2348) begin
      useRAS_9 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2354) begin
      useRAS_8 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2360) begin
      useRAS_7 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2366) begin
      useRAS_6 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2372) begin
      useRAS_5 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2378) begin
      useRAS_4 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2384) begin
      useRAS_3 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2390) begin
      useRAS_2 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2396) begin
      useRAS_1 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(T2401) begin
      useRAS_0 <= R2032;
    end 
  end


  always @(posedge clk) begin
    if(N2306) begin
      brIdx[61] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2305) begin
      brIdx[60] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2304) begin
      brIdx[59] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2303) begin
      brIdx[58] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2302) begin
      brIdx[57] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2301) begin
      brIdx[56] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2300) begin
      brIdx[55] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2299) begin
      brIdx[54] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2298) begin
      brIdx[53] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2297) begin
      brIdx[52] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2296) begin
      brIdx[51] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2295) begin
      brIdx[50] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2294) begin
      brIdx[49] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2293) begin
      brIdx[48] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2292) begin
      brIdx[47] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2291) begin
      brIdx[46] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2290) begin
      brIdx[45] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2289) begin
      brIdx[44] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2288) begin
      brIdx[43] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2287) begin
      brIdx[42] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2286) begin
      brIdx[41] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2285) begin
      brIdx[40] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2284) begin
      brIdx[39] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2283) begin
      brIdx[38] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2282) begin
      brIdx[37] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2281) begin
      brIdx[36] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2280) begin
      brIdx[35] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2279) begin
      brIdx[34] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2278) begin
      brIdx[33] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2277) begin
      brIdx[32] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2276) begin
      brIdx[31] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2275) begin
      brIdx[30] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2274) begin
      brIdx[29] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2273) begin
      brIdx[28] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2272) begin
      brIdx[27] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2271) begin
      brIdx[26] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2270) begin
      brIdx[25] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2269) begin
      brIdx[24] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2268) begin
      brIdx[23] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2267) begin
      brIdx[22] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2266) begin
      brIdx[21] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2265) begin
      brIdx[20] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2264) begin
      brIdx[19] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2263) begin
      brIdx[18] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2262) begin
      brIdx[17] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2261) begin
      brIdx[16] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2260) begin
      brIdx[15] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2259) begin
      brIdx[14] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2258) begin
      brIdx[13] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2257) begin
      brIdx[12] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2256) begin
      brIdx[11] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2255) begin
      brIdx[10] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2254) begin
      brIdx[9] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2253) begin
      brIdx[8] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2252) begin
      brIdx[7] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2251) begin
      brIdx[6] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2250) begin
      brIdx[5] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2249) begin
      brIdx[4] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2248) begin
      brIdx[3] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2247) begin
      brIdx[2] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2246) begin
      brIdx[1] <= 1'b0;
    end 
  end


  always @(posedge clk) begin
    if(N2245) begin
      brIdx[0] <= 1'b0;
    end 
  end

  assign N2328 = T195[5] | T2420[0];
  assign N2329 = T195[3] | T195[4];
  assign N2330 = T799[4] | T799[5];
  assign N2331 = T2444[2] | T2444[3];
  assign N2332 = hits[60] | hits[61];
  assign N2333 = hits[59] | N2332;
  assign N2334 = hits[58] | N2333;
  assign N2335 = hits[57] | N2334;
  assign N2336 = hits[56] | N2335;
  assign N2337 = hits[55] | N2336;
  assign N2338 = hits[54] | N2337;
  assign N2339 = hits[53] | N2338;
  assign N2340 = hits[52] | N2339;
  assign N2341 = hits[51] | N2340;
  assign N2342 = hits[50] | N2341;
  assign N2343 = hits[49] | N2342;
  assign N2344 = hits[48] | N2343;
  assign N2345 = hits[47] | N2344;
  assign N2346 = hits[46] | N2345;
  assign N2347 = hits[45] | N2346;
  assign N2348 = hits[44] | N2347;
  assign N2349 = hits[43] | N2348;
  assign N2350 = hits[42] | N2349;
  assign N2351 = hits[41] | N2350;
  assign N2352 = hits[40] | N2351;
  assign N2353 = hits[39] | N2352;
  assign N2354 = hits[38] | N2353;
  assign N2355 = hits[37] | N2354;
  assign N2356 = hits[36] | N2355;
  assign N2357 = hits[35] | N2356;
  assign N2358 = hits[34] | N2357;
  assign N2359 = hits[33] | N2358;
  assign io_resp_bits_entry[5] = hits[32] | N2359;
  assign N2361 = hits[30] | hits[31];
  assign N2362 = T2464[29] | N2361;
  assign N2363 = T2464[28] | N2362;
  assign N2364 = T2464[27] | N2363;
  assign N2365 = T2464[26] | N2364;
  assign N2366 = T2464[25] | N2365;
  assign N2367 = T2464[24] | N2366;
  assign N2368 = T2464[23] | N2367;
  assign N2369 = T2464[22] | N2368;
  assign N2370 = T2464[21] | N2369;
  assign N2371 = T2464[20] | N2370;
  assign N2372 = T2464[19] | N2371;
  assign N2373 = T2464[18] | N2372;
  assign N2374 = T2464[17] | N2373;
  assign io_resp_bits_entry[4] = T2464[16] | N2374;
  assign N2376 = T2462[14] | T2462[15];
  assign N2377 = T2462[13] | N2376;
  assign N2378 = T2462[12] | N2377;
  assign N2379 = T2462[11] | N2378;
  assign N2380 = T2462[10] | N2379;
  assign N2381 = T2462[9] | N2380;
  assign io_resp_bits_entry[3] = T2462[8] | N2381;
  assign N2383 = ~nextRepl[5];
  assign N2384 = ~nextRepl[4];
  assign N2385 = ~nextRepl[3];
  assign N2386 = ~nextRepl[2];
  assign N2387 = ~nextRepl[0];
  assign N2388 = N2384 | N2383;
  assign N2389 = N2385 | N2388;
  assign N2390 = N2386 | N2389;
  assign N2391 = nextRepl[1] | N2390;
  assign N2392 = N2387 | N2391;
  assign N2393 = ~N2392;
  assign N2394 = ~R198[2];
  assign N2395 = ~R198[0];
  assign N2396 = R198[1] | N2394;
  assign N2397 = N2395 | N2396;
  assign N2398 = ~N2397;
  assign T783 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T169;
  assign T168 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T169;
  assign T2036 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T169;
  assign N2399 = T2460[6] | T2460[7];
  assign N2400 = T2460[5] | N2399;
  assign io_resp_bits_entry[2] = T2460[4] | N2400;
  assign N2402 = R2010[0] | R2010[1];
  assign N2403 = ~N2402;
  assign io_resp_bits_entry[1] = T2458[2] | T2458[3];
  assign N2405 = hits[60] | hits[61];
  assign N2406 = hits[59] | N2405;
  assign N2407 = hits[58] | N2406;
  assign N2408 = hits[57] | N2407;
  assign N2409 = hits[56] | N2408;
  assign N2410 = hits[55] | N2409;
  assign N2411 = hits[54] | N2410;
  assign N2412 = hits[53] | N2411;
  assign N2413 = hits[52] | N2412;
  assign N2414 = hits[51] | N2413;
  assign N2415 = hits[50] | N2414;
  assign N2416 = hits[49] | N2415;
  assign N2417 = hits[48] | N2416;
  assign N2418 = hits[47] | N2417;
  assign N2419 = hits[46] | N2418;
  assign N2420 = hits[45] | N2419;
  assign N2421 = hits[44] | N2420;
  assign N2422 = hits[43] | N2421;
  assign N2423 = hits[42] | N2422;
  assign N2424 = hits[41] | N2423;
  assign N2425 = hits[40] | N2424;
  assign N2426 = hits[39] | N2425;
  assign N2427 = hits[38] | N2426;
  assign N2428 = hits[37] | N2427;
  assign N2429 = hits[36] | N2428;
  assign N2430 = hits[35] | N2429;
  assign N2431 = hits[34] | N2430;
  assign N2432 = hits[33] | N2431;
  assign N2433 = hits[32] | N2432;
  assign N2434 = hits[31] | N2433;
  assign N2435 = hits[30] | N2434;
  assign N2436 = hits[29] | N2435;
  assign N2437 = hits[28] | N2436;
  assign N2438 = hits[27] | N2437;
  assign N2439 = hits[26] | N2438;
  assign N2440 = hits[25] | N2439;
  assign N2441 = hits[24] | N2440;
  assign N2442 = hits[23] | N2441;
  assign N2443 = hits[22] | N2442;
  assign N2444 = hits[21] | N2443;
  assign N2445 = hits[20] | N2444;
  assign N2446 = hits[19] | N2445;
  assign N2447 = hits[18] | N2446;
  assign N2448 = hits[17] | N2447;
  assign N2449 = hits[16] | N2448;
  assign N2450 = hits[15] | N2449;
  assign N2451 = hits[14] | N2450;
  assign N2452 = hits[13] | N2451;
  assign N2453 = hits[12] | N2452;
  assign N2454 = hits[11] | N2453;
  assign N2455 = hits[10] | N2454;
  assign N2456 = hits[9] | N2455;
  assign N2457 = hits[8] | N2456;
  assign N2458 = hits[7] | N2457;
  assign N2459 = hits[6] | N2458;
  assign N2460 = hits[5] | N2459;
  assign N2461 = hits[4] | N2460;
  assign N2462 = hits[3] | N2461;
  assign N2463 = hits[2] | N2462;
  assign N2464 = hits[1] | N2463;
  assign io_resp_valid = hits[0] | N2464;
  assign N2466 = T1158[4] | T1158[5];
  assign N2467 = T1158[3] | N2466;
  assign N2468 = T1158[2] | N2467;
  assign N2469 = T1158[1] | N2468;
  assign N2470 = T1158[0] | N2469;
  assign N2471 = T1153[4] | T1153[5];
  assign N2472 = T1153[3] | N2471;
  assign N2473 = T1153[2] | N2472;
  assign N2474 = T1153[1] | N2473;
  assign N2475 = T1153[0] | N2474;
  assign N2476 = T1148[4] | T1148[5];
  assign N2477 = T1148[3] | N2476;
  assign N2478 = T1148[2] | N2477;
  assign N2479 = T1148[1] | N2478;
  assign N2480 = T1148[0] | N2479;
  assign N2481 = T1141[4] | T1141[5];
  assign N2482 = T1141[3] | N2481;
  assign N2483 = T1141[2] | N2482;
  assign N2484 = T1141[1] | N2483;
  assign N2485 = T1141[0] | N2484;
  assign N2486 = T1136[4] | T1136[5];
  assign N2487 = T1136[3] | N2486;
  assign N2488 = T1136[2] | N2487;
  assign N2489 = T1136[1] | N2488;
  assign N2490 = T1136[0] | N2489;
  assign N2491 = T1130[4] | T1130[5];
  assign N2492 = T1130[3] | N2491;
  assign N2493 = T1130[2] | N2492;
  assign N2494 = T1130[1] | N2493;
  assign N2495 = T1130[0] | N2494;
  assign N2496 = T1125[4] | T1125[5];
  assign N2497 = T1125[3] | N2496;
  assign N2498 = T1125[2] | N2497;
  assign N2499 = T1125[1] | N2498;
  assign N2500 = T1125[0] | N2499;
  assign N2501 = T1117[4] | T1117[5];
  assign N2502 = T1117[3] | N2501;
  assign N2503 = T1117[2] | N2502;
  assign N2504 = T1117[1] | N2503;
  assign N2505 = T1117[0] | N2504;
  assign N2506 = T1112[4] | T1112[5];
  assign N2507 = T1112[3] | N2506;
  assign N2508 = T1112[2] | N2507;
  assign N2509 = T1112[1] | N2508;
  assign N2510 = T1112[0] | N2509;
  assign N2511 = T1106[4] | T1106[5];
  assign N2512 = T1106[3] | N2511;
  assign N2513 = T1106[2] | N2512;
  assign N2514 = T1106[1] | N2513;
  assign N2515 = T1106[0] | N2514;
  assign N2516 = T1101[4] | T1101[5];
  assign N2517 = T1101[3] | N2516;
  assign N2518 = T1101[2] | N2517;
  assign N2519 = T1101[1] | N2518;
  assign N2520 = T1101[0] | N2519;
  assign N2521 = T1094[4] | T1094[5];
  assign N2522 = T1094[3] | N2521;
  assign N2523 = T1094[2] | N2522;
  assign N2524 = T1094[1] | N2523;
  assign N2525 = T1094[0] | N2524;
  assign N2526 = T1089[4] | T1089[5];
  assign N2527 = T1089[3] | N2526;
  assign N2528 = T1089[2] | N2527;
  assign N2529 = T1089[1] | N2528;
  assign N2530 = T1089[0] | N2529;
  assign N2531 = T1083[4] | T1083[5];
  assign N2532 = T1083[3] | N2531;
  assign N2533 = T1083[2] | N2532;
  assign N2534 = T1083[1] | N2533;
  assign N2535 = T1083[0] | N2534;
  assign N2536 = T1078[4] | T1078[5];
  assign N2537 = T1078[3] | N2536;
  assign N2538 = T1078[2] | N2537;
  assign N2539 = T1078[1] | N2538;
  assign N2540 = T1078[0] | N2539;
  assign N2541 = T1069[4] | T1069[5];
  assign N2542 = T1069[3] | N2541;
  assign N2543 = T1069[2] | N2542;
  assign N2544 = T1069[1] | N2543;
  assign N2545 = T1069[0] | N2544;
  assign N2546 = T1064[4] | T1064[5];
  assign N2547 = T1064[3] | N2546;
  assign N2548 = T1064[2] | N2547;
  assign N2549 = T1064[1] | N2548;
  assign N2550 = T1064[0] | N2549;
  assign N2551 = T1058[4] | T1058[5];
  assign N2552 = T1058[3] | N2551;
  assign N2553 = T1058[2] | N2552;
  assign N2554 = T1058[1] | N2553;
  assign N2555 = T1058[0] | N2554;
  assign N2556 = T1053[4] | T1053[5];
  assign N2557 = T1053[3] | N2556;
  assign N2558 = T1053[2] | N2557;
  assign N2559 = T1053[1] | N2558;
  assign N2560 = T1053[0] | N2559;
  assign N2561 = T1046[4] | T1046[5];
  assign N2562 = T1046[3] | N2561;
  assign N2563 = T1046[2] | N2562;
  assign N2564 = T1046[1] | N2563;
  assign N2565 = T1046[0] | N2564;
  assign N2566 = T1041[4] | T1041[5];
  assign N2567 = T1041[3] | N2566;
  assign N2568 = T1041[2] | N2567;
  assign N2569 = T1041[1] | N2568;
  assign N2570 = T1041[0] | N2569;
  assign N2571 = T1035[4] | T1035[5];
  assign N2572 = T1035[3] | N2571;
  assign N2573 = T1035[2] | N2572;
  assign N2574 = T1035[1] | N2573;
  assign N2575 = T1035[0] | N2574;
  assign N2576 = T1030[4] | T1030[5];
  assign N2577 = T1030[3] | N2576;
  assign N2578 = T1030[2] | N2577;
  assign N2579 = T1030[1] | N2578;
  assign N2580 = T1030[0] | N2579;
  assign N2581 = T1022[4] | T1022[5];
  assign N2582 = T1022[3] | N2581;
  assign N2583 = T1022[2] | N2582;
  assign N2584 = T1022[1] | N2583;
  assign N2585 = T1022[0] | N2584;
  assign N2586 = T1017[4] | T1017[5];
  assign N2587 = T1017[3] | N2586;
  assign N2588 = T1017[2] | N2587;
  assign N2589 = T1017[1] | N2588;
  assign N2590 = T1017[0] | N2589;
  assign N2591 = T1011[4] | T1011[5];
  assign N2592 = T1011[3] | N2591;
  assign N2593 = T1011[2] | N2592;
  assign N2594 = T1011[1] | N2593;
  assign N2595 = T1011[0] | N2594;
  assign N2596 = T1006[4] | T1006[5];
  assign N2597 = T1006[3] | N2596;
  assign N2598 = T1006[2] | N2597;
  assign N2599 = T1006[1] | N2598;
  assign N2600 = T1006[0] | N2599;
  assign N2601 = T999[4] | T999[5];
  assign N2602 = T999[3] | N2601;
  assign N2603 = T999[2] | N2602;
  assign N2604 = T999[1] | N2603;
  assign N2605 = T999[0] | N2604;
  assign N2606 = T994[4] | T994[5];
  assign N2607 = T994[3] | N2606;
  assign N2608 = T994[2] | N2607;
  assign N2609 = T994[1] | N2608;
  assign N2610 = T994[0] | N2609;
  assign N2611 = T988[4] | T988[5];
  assign N2612 = T988[3] | N2611;
  assign N2613 = T988[2] | N2612;
  assign N2614 = T988[1] | N2613;
  assign N2615 = T988[0] | N2614;
  assign N2616 = T983[4] | T983[5];
  assign N2617 = T983[3] | N2616;
  assign N2618 = T983[2] | N2617;
  assign N2619 = T983[1] | N2618;
  assign N2620 = T983[0] | N2619;
  assign N2621 = T973[4] | T973[5];
  assign N2622 = T973[3] | N2621;
  assign N2623 = T973[2] | N2622;
  assign N2624 = T973[1] | N2623;
  assign N2625 = T973[0] | N2624;
  assign N2626 = T968[4] | T968[5];
  assign N2627 = T968[3] | N2626;
  assign N2628 = T968[2] | N2627;
  assign N2629 = T968[1] | N2628;
  assign N2630 = T968[0] | N2629;
  assign N2631 = T963[4] | T963[5];
  assign N2632 = T963[3] | N2631;
  assign N2633 = T963[2] | N2632;
  assign N2634 = T963[1] | N2633;
  assign N2635 = T963[0] | N2634;
  assign N2636 = T956[4] | T956[5];
  assign N2637 = T956[3] | N2636;
  assign N2638 = T956[2] | N2637;
  assign N2639 = T956[1] | N2638;
  assign N2640 = T956[0] | N2639;
  assign N2641 = T951[4] | T951[5];
  assign N2642 = T951[3] | N2641;
  assign N2643 = T951[2] | N2642;
  assign N2644 = T951[1] | N2643;
  assign N2645 = T951[0] | N2644;
  assign N2646 = T945[4] | T945[5];
  assign N2647 = T945[3] | N2646;
  assign N2648 = T945[2] | N2647;
  assign N2649 = T945[1] | N2648;
  assign N2650 = T945[0] | N2649;
  assign N2651 = T940[4] | T940[5];
  assign N2652 = T940[3] | N2651;
  assign N2653 = T940[2] | N2652;
  assign N2654 = T940[1] | N2653;
  assign N2655 = T940[0] | N2654;
  assign N2656 = T932[4] | T932[5];
  assign N2657 = T932[3] | N2656;
  assign N2658 = T932[2] | N2657;
  assign N2659 = T932[1] | N2658;
  assign N2660 = T932[0] | N2659;
  assign N2661 = T927[4] | T927[5];
  assign N2662 = T927[3] | N2661;
  assign N2663 = T927[2] | N2662;
  assign N2664 = T927[1] | N2663;
  assign N2665 = T927[0] | N2664;
  assign N2666 = T921[4] | T921[5];
  assign N2667 = T921[3] | N2666;
  assign N2668 = T921[2] | N2667;
  assign N2669 = T921[1] | N2668;
  assign N2670 = T921[0] | N2669;
  assign N2671 = T916[4] | T916[5];
  assign N2672 = T916[3] | N2671;
  assign N2673 = T916[2] | N2672;
  assign N2674 = T916[1] | N2673;
  assign N2675 = T916[0] | N2674;
  assign N2676 = T909[4] | T909[5];
  assign N2677 = T909[3] | N2676;
  assign N2678 = T909[2] | N2677;
  assign N2679 = T909[1] | N2678;
  assign N2680 = T909[0] | N2679;
  assign N2681 = T904[4] | T904[5];
  assign N2682 = T904[3] | N2681;
  assign N2683 = T904[2] | N2682;
  assign N2684 = T904[1] | N2683;
  assign N2685 = T904[0] | N2684;
  assign N2686 = T898[4] | T898[5];
  assign N2687 = T898[3] | N2686;
  assign N2688 = T898[2] | N2687;
  assign N2689 = T898[1] | N2688;
  assign N2690 = T898[0] | N2689;
  assign N2691 = T893[4] | T893[5];
  assign N2692 = T893[3] | N2691;
  assign N2693 = T893[2] | N2692;
  assign N2694 = T893[1] | N2693;
  assign N2695 = T893[0] | N2694;
  assign N2696 = T884[4] | T884[5];
  assign N2697 = T884[3] | N2696;
  assign N2698 = T884[2] | N2697;
  assign N2699 = T884[1] | N2698;
  assign N2700 = T884[0] | N2699;
  assign N2701 = T879[4] | T879[5];
  assign N2702 = T879[3] | N2701;
  assign N2703 = T879[2] | N2702;
  assign N2704 = T879[1] | N2703;
  assign N2705 = T879[0] | N2704;
  assign N2706 = T873[4] | T873[5];
  assign N2707 = T873[3] | N2706;
  assign N2708 = T873[2] | N2707;
  assign N2709 = T873[1] | N2708;
  assign N2710 = T873[0] | N2709;
  assign N2711 = T868[4] | T868[5];
  assign N2712 = T868[3] | N2711;
  assign N2713 = T868[2] | N2712;
  assign N2714 = T868[1] | N2713;
  assign N2715 = T868[0] | N2714;
  assign N2716 = T861[4] | T861[5];
  assign N2717 = T861[3] | N2716;
  assign N2718 = T861[2] | N2717;
  assign N2719 = T861[1] | N2718;
  assign N2720 = T861[0] | N2719;
  assign N2721 = T856[4] | T856[5];
  assign N2722 = T856[3] | N2721;
  assign N2723 = T856[2] | N2722;
  assign N2724 = T856[1] | N2723;
  assign N2725 = T856[0] | N2724;
  assign N2726 = T850[4] | T850[5];
  assign N2727 = T850[3] | N2726;
  assign N2728 = T850[2] | N2727;
  assign N2729 = T850[1] | N2728;
  assign N2730 = T850[0] | N2729;
  assign N2731 = T845[4] | T845[5];
  assign N2732 = T845[3] | N2731;
  assign N2733 = T845[2] | N2732;
  assign N2734 = T845[1] | N2733;
  assign N2735 = T845[0] | N2734;
  assign N2736 = T837[4] | T837[5];
  assign N2737 = T837[3] | N2736;
  assign N2738 = T837[2] | N2737;
  assign N2739 = T837[1] | N2738;
  assign N2740 = T837[0] | N2739;
  assign N2741 = T832[4] | T832[5];
  assign N2742 = T832[3] | N2741;
  assign N2743 = T832[2] | N2742;
  assign N2744 = T832[1] | N2743;
  assign N2745 = T832[0] | N2744;
  assign N2746 = T826[4] | T826[5];
  assign N2747 = T826[3] | N2746;
  assign N2748 = T826[2] | N2747;
  assign N2749 = T826[1] | N2748;
  assign N2750 = T826[0] | N2749;
  assign N2751 = T821[4] | T821[5];
  assign N2752 = T821[3] | N2751;
  assign N2753 = T821[2] | N2752;
  assign N2754 = T821[1] | N2753;
  assign N2755 = T821[0] | N2754;
  assign N2756 = T814[4] | T814[5];
  assign N2757 = T814[3] | N2756;
  assign N2758 = T814[2] | N2757;
  assign N2759 = T814[1] | N2758;
  assign N2760 = T814[0] | N2759;
  assign N2761 = T809[4] | T809[5];
  assign N2762 = T809[3] | N2761;
  assign N2763 = T809[2] | N2762;
  assign N2764 = T809[1] | N2763;
  assign N2765 = T809[0] | N2764;
  assign N2766 = T803[4] | T803[5];
  assign N2767 = T803[3] | N2766;
  assign N2768 = T803[2] | N2767;
  assign N2769 = T803[1] | N2768;
  assign N2770 = T803[0] | N2769;
  assign N2771 = T794[4] | T794[5];
  assign N2772 = T794[3] | N2771;
  assign N2773 = T794[2] | N2772;
  assign N2774 = T794[1] | N2773;
  assign N2775 = T794[0] | N2774;
  assign N2776 = R2010[0] | R2010[1];
  assign N2777 = ~N2776;
  assign N2778 = T195[3] | T195[5];
  assign N2779 = T195[1] | N2778;
  assign tgtPagesOH_61 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1161;
  assign tgtPagesOH_60 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1156;
  assign tgtPagesOH_59 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1151;
  assign tgtPagesOH_58 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1144;
  assign N2780 = T586[4] | T586[5];
  assign N2781 = T586[3] | N2780;
  assign N2782 = T586[2] | N2781;
  assign N2783 = T586[1] | N2782;
  assign N2784 = T586[0] | N2783;
  assign N2785 = T262[4] | T262[5];
  assign N2786 = T262[3] | N2785;
  assign N2787 = T262[2] | N2786;
  assign N2788 = T262[1] | N2787;
  assign N2789 = T262[0] | N2788;
  assign tgtPagesOH_57 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1139;
  assign N2790 = T582[4] | T582[5];
  assign N2791 = T582[3] | N2790;
  assign N2792 = T582[2] | N2791;
  assign N2793 = T582[1] | N2792;
  assign N2794 = T582[0] | N2793;
  assign tgtPagesOH_56 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1133;
  assign N2795 = T578[4] | T578[5];
  assign N2796 = T578[3] | N2795;
  assign N2797 = T578[2] | N2796;
  assign N2798 = T578[1] | N2797;
  assign N2799 = T578[0] | N2798;
  assign idxPagesOH_61 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T588;
  assign tgtPagesOH_55 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1128;
  assign N2800 = T572[4] | T572[5];
  assign N2801 = T572[3] | N2800;
  assign N2802 = T572[2] | N2801;
  assign N2803 = T572[1] | N2802;
  assign N2804 = T572[0] | N2803;
  assign idxPagesOH_60 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T584;
  assign tgtPagesOH_54 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1120;
  assign N2805 = T568[4] | T568[5];
  assign N2806 = T568[3] | N2805;
  assign N2807 = T568[2] | N2806;
  assign N2808 = T568[1] | N2807;
  assign N2809 = T568[0] | N2808;
  assign idxPagesOH_59 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T580;
  assign idxPageRepl = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << R198;
  assign tgtPagesOH_53 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1115;
  assign N2810 = T563[4] | T563[5];
  assign N2811 = T563[3] | N2810;
  assign N2812 = T563[2] | N2811;
  assign N2813 = T563[1] | N2812;
  assign N2814 = T563[0] | N2813;
  assign idxPagesOH_58 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T574;
  assign tgtPagesOH_52 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1109;
  assign N2815 = T559[4] | T559[5];
  assign N2816 = T559[3] | N2815;
  assign N2817 = T559[2] | N2816;
  assign N2818 = T559[1] | N2817;
  assign N2819 = T559[0] | N2818;
  assign idxPagesOH_57 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T570;
  assign tgtPagesOH_51 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1104;
  assign N2820 = T552[4] | T552[5];
  assign N2821 = T552[3] | N2820;
  assign N2822 = T552[2] | N2821;
  assign N2823 = T552[1] | N2822;
  assign N2824 = T552[0] | N2823;
  assign idxPagesOH_56 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T565;
  assign N2825 = updatePageHit[4] | updatePageHit[5];
  assign N2826 = updatePageHit[3] | N2825;
  assign N2827 = updatePageHit[2] | N2826;
  assign N2828 = updatePageHit[1] | N2827;
  assign N2829 = updatePageHit[0] | N2828;
  assign tgtPagesOH_50 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1097;
  assign N2830 = T548[4] | T548[5];
  assign N2831 = T548[3] | N2830;
  assign N2832 = T548[2] | N2831;
  assign N2833 = T548[1] | N2832;
  assign N2834 = T548[0] | N2833;
  assign idxPagesOH_55 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T561;
  assign tgtPagesOH_49 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1092;
  assign N2835 = T543[4] | T543[5];
  assign N2836 = T543[3] | N2835;
  assign N2837 = T543[2] | N2836;
  assign N2838 = T543[1] | N2837;
  assign N2839 = T543[0] | N2838;
  assign idxPagesOH_54 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T554;
  assign tgtPagesOH_48 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1086;
  assign N2840 = T539[4] | T539[5];
  assign N2841 = T539[3] | N2840;
  assign N2842 = T539[2] | N2841;
  assign N2843 = T539[1] | N2842;
  assign N2844 = T539[0] | N2843;
  assign idxPagesOH_53 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T550;
  assign tgtPagesOH_47 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1081;
  assign N2845 = T533[4] | T533[5];
  assign N2846 = T533[3] | N2845;
  assign N2847 = T533[2] | N2846;
  assign N2848 = T533[1] | N2847;
  assign N2849 = T533[0] | N2848;
  assign idxPagesOH_52 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T545;
  assign tgtPagesOH_46 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1072;
  assign N2850 = T529[4] | T529[5];
  assign N2851 = T529[3] | N2850;
  assign N2852 = T529[2] | N2851;
  assign N2853 = T529[1] | N2852;
  assign N2854 = T529[0] | N2853;
  assign idxPagesOH_51 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T541;
  assign tgtPagesOH_45 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1067;
  assign N2855 = T524[4] | T524[5];
  assign N2856 = T524[3] | N2855;
  assign N2857 = T524[2] | N2856;
  assign N2858 = T524[1] | N2857;
  assign N2859 = T524[0] | N2858;
  assign idxPagesOH_50 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T535;
  assign tgtPagesOH_44 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1061;
  assign N2860 = T520[4] | T520[5];
  assign N2861 = T520[3] | N2860;
  assign N2862 = T520[2] | N2861;
  assign N2863 = T520[1] | N2862;
  assign N2864 = T520[0] | N2863;
  assign idxPagesOH_49 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T531;
  assign tgtPagesOH_43 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1056;
  assign N2865 = T512[4] | T512[5];
  assign N2866 = T512[3] | N2865;
  assign N2867 = T512[2] | N2866;
  assign N2868 = T512[1] | N2867;
  assign N2869 = T512[0] | N2868;
  assign idxPagesOH_48 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T526;
  assign tgtPagesOH_42 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1049;
  assign N2870 = T508[4] | T508[5];
  assign N2871 = T508[3] | N2870;
  assign N2872 = T508[2] | N2871;
  assign N2873 = T508[1] | N2872;
  assign N2874 = T508[0] | N2873;
  assign idxPagesOH_47 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T522;
  assign tgtPagesOH_41 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1044;
  assign N2875 = T503[4] | T503[5];
  assign N2876 = T503[3] | N2875;
  assign N2877 = T503[2] | N2876;
  assign N2878 = T503[1] | N2877;
  assign N2879 = T503[0] | N2878;
  assign idxPagesOH_46 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T514;
  assign tgtPagesOH_40 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1038;
  assign N2880 = T499[4] | T499[5];
  assign N2881 = T499[3] | N2880;
  assign N2882 = T499[2] | N2881;
  assign N2883 = T499[1] | N2882;
  assign N2884 = T499[0] | N2883;
  assign idxPagesOH_45 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T510;
  assign tgtPagesOH_39 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1033;
  assign N2885 = T493[4] | T493[5];
  assign N2886 = T493[3] | N2885;
  assign N2887 = T493[2] | N2886;
  assign N2888 = T493[1] | N2887;
  assign N2889 = T493[0] | N2888;
  assign idxPagesOH_44 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T505;
  assign tgtPagesOH_38 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1025;
  assign N2890 = T489[4] | T489[5];
  assign N2891 = T489[3] | N2890;
  assign N2892 = T489[2] | N2891;
  assign N2893 = T489[1] | N2892;
  assign N2894 = T489[0] | N2893;
  assign idxPagesOH_43 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T501;
  assign tgtPagesOH_37 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1020;
  assign N2895 = T484[4] | T484[5];
  assign N2896 = T484[3] | N2895;
  assign N2897 = T484[2] | N2896;
  assign N2898 = T484[1] | N2897;
  assign N2899 = T484[0] | N2898;
  assign idxPagesOH_42 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T495;
  assign tgtPagesOH_36 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1014;
  assign N2900 = T480[4] | T480[5];
  assign N2901 = T480[3] | N2900;
  assign N2902 = T480[2] | N2901;
  assign N2903 = T480[1] | N2902;
  assign N2904 = T480[0] | N2903;
  assign idxPagesOH_41 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T491;
  assign tgtPagesOH_35 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1009;
  assign N2905 = T473[4] | T473[5];
  assign N2906 = T473[3] | N2905;
  assign N2907 = T473[2] | N2906;
  assign N2908 = T473[1] | N2907;
  assign N2909 = T473[0] | N2908;
  assign idxPagesOH_40 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T486;
  assign tgtPagesOH_34 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T1002;
  assign N2910 = T469[4] | T469[5];
  assign N2911 = T469[3] | N2910;
  assign N2912 = T469[2] | N2911;
  assign N2913 = T469[1] | N2912;
  assign N2914 = T469[0] | N2913;
  assign idxPagesOH_39 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T482;
  assign tgtPagesOH_33 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T997;
  assign N2915 = T464[4] | T464[5];
  assign N2916 = T464[3] | N2915;
  assign N2917 = T464[2] | N2916;
  assign N2918 = T464[1] | N2917;
  assign N2919 = T464[0] | N2918;
  assign idxPagesOH_38 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T475;
  assign tgtPagesOH_32 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T991;
  assign N2920 = T460[4] | T460[5];
  assign N2921 = T460[3] | N2920;
  assign N2922 = T460[2] | N2921;
  assign N2923 = T460[1] | N2922;
  assign N2924 = T460[0] | N2923;
  assign idxPagesOH_37 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T471;
  assign tgtPagesOH_31 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T986;
  assign N2925 = T454[4] | T454[5];
  assign N2926 = T454[3] | N2925;
  assign N2927 = T454[2] | N2926;
  assign N2928 = T454[1] | N2927;
  assign N2929 = T454[0] | N2928;
  assign idxPagesOH_36 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T466;
  assign tgtPagesOH_30 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T976;
  assign N2930 = T450[4] | T450[5];
  assign N2931 = T450[3] | N2930;
  assign N2932 = T450[2] | N2931;
  assign N2933 = T450[1] | N2932;
  assign N2934 = T450[0] | N2933;
  assign idxPagesOH_35 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T462;
  assign tgtPagesOH_29 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T971;
  assign N2935 = T445[4] | T445[5];
  assign N2936 = T445[3] | N2935;
  assign N2937 = T445[2] | N2936;
  assign N2938 = T445[1] | N2937;
  assign N2939 = T445[0] | N2938;
  assign idxPagesOH_34 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T456;
  assign tgtPagesOH_28 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T966;
  assign N2940 = T441[4] | T441[5];
  assign N2941 = T441[3] | N2940;
  assign N2942 = T441[2] | N2941;
  assign N2943 = T441[1] | N2942;
  assign N2944 = T441[0] | N2943;
  assign idxPagesOH_33 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T452;
  assign tgtPagesOH_27 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T959;
  assign N2945 = T432[4] | T432[5];
  assign N2946 = T432[3] | N2945;
  assign N2947 = T432[2] | N2946;
  assign N2948 = T432[1] | N2947;
  assign N2949 = T432[0] | N2948;
  assign idxPagesOH_32 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T447;
  assign tgtPagesOH_26 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T954;
  assign N2950 = T428[4] | T428[5];
  assign N2951 = T428[3] | N2950;
  assign N2952 = T428[2] | N2951;
  assign N2953 = T428[1] | N2952;
  assign N2954 = T428[0] | N2953;
  assign idxPagesOH_31 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T443;
  assign tgtPagesOH_25 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T948;
  assign N2955 = T424[4] | T424[5];
  assign N2956 = T424[3] | N2955;
  assign N2957 = T424[2] | N2956;
  assign N2958 = T424[1] | N2957;
  assign N2959 = T424[0] | N2958;
  assign idxPagesOH_30 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T434;
  assign tgtPagesOH_24 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T943;
  assign N2960 = T418[4] | T418[5];
  assign N2961 = T418[3] | N2960;
  assign N2962 = T418[2] | N2961;
  assign N2963 = T418[1] | N2962;
  assign N2964 = T418[0] | N2963;
  assign idxPagesOH_29 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T430;
  assign tgtPagesOH_23 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T935;
  assign N2965 = T414[4] | T414[5];
  assign N2966 = T414[3] | N2965;
  assign N2967 = T414[2] | N2966;
  assign N2968 = T414[1] | N2967;
  assign N2969 = T414[0] | N2968;
  assign idxPagesOH_28 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T426;
  assign tgtPagesOH_22 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T930;
  assign N2970 = T409[4] | T409[5];
  assign N2971 = T409[3] | N2970;
  assign N2972 = T409[2] | N2971;
  assign N2973 = T409[1] | N2972;
  assign N2974 = T409[0] | N2973;
  assign idxPagesOH_27 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T420;
  assign tgtPagesOH_21 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T924;
  assign N2975 = T405[4] | T405[5];
  assign N2976 = T405[3] | N2975;
  assign N2977 = T405[2] | N2976;
  assign N2978 = T405[1] | N2977;
  assign N2979 = T405[0] | N2978;
  assign idxPagesOH_26 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T416;
  assign tgtPagesOH_20 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T919;
  assign N2980 = T398[4] | T398[5];
  assign N2981 = T398[3] | N2980;
  assign N2982 = T398[2] | N2981;
  assign N2983 = T398[1] | N2982;
  assign N2984 = T398[0] | N2983;
  assign idxPagesOH_25 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T411;
  assign tgtPagesOH_19 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T912;
  assign N2985 = T394[4] | T394[5];
  assign N2986 = T394[3] | N2985;
  assign N2987 = T394[2] | N2986;
  assign N2988 = T394[1] | N2987;
  assign N2989 = T394[0] | N2988;
  assign idxPagesOH_24 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T407;
  assign tgtPagesOH_18 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T907;
  assign N2990 = T389[4] | T389[5];
  assign N2991 = T389[3] | N2990;
  assign N2992 = T389[2] | N2991;
  assign N2993 = T389[1] | N2992;
  assign N2994 = T389[0] | N2993;
  assign idxPagesOH_23 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T400;
  assign tgtPagesOH_17 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T901;
  assign N2995 = T385[4] | T385[5];
  assign N2996 = T385[3] | N2995;
  assign N2997 = T385[2] | N2996;
  assign N2998 = T385[1] | N2997;
  assign N2999 = T385[0] | N2998;
  assign idxPagesOH_22 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T396;
  assign tgtPagesOH_16 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T896;
  assign N3000 = T379[4] | T379[5];
  assign N3001 = T379[3] | N3000;
  assign N3002 = T379[2] | N3001;
  assign N3003 = T379[1] | N3002;
  assign N3004 = T379[0] | N3003;
  assign idxPagesOH_21 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T391;
  assign tgtPagesOH_15 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T887;
  assign N3005 = T375[4] | T375[5];
  assign N3006 = T375[3] | N3005;
  assign N3007 = T375[2] | N3006;
  assign N3008 = T375[1] | N3007;
  assign N3009 = T375[0] | N3008;
  assign idxPagesOH_20 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T387;
  assign tgtPagesOH_14 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T882;
  assign N3010 = T370[4] | T370[5];
  assign N3011 = T370[3] | N3010;
  assign N3012 = T370[2] | N3011;
  assign N3013 = T370[1] | N3012;
  assign N3014 = T370[0] | N3013;
  assign idxPagesOH_19 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T381;
  assign tgtPagesOH_13 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T876;
  assign N3015 = T366[4] | T366[5];
  assign N3016 = T366[3] | N3015;
  assign N3017 = T366[2] | N3016;
  assign N3018 = T366[1] | N3017;
  assign N3019 = T366[0] | N3018;
  assign idxPagesOH_18 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T377;
  assign tgtPagesOH_12 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T871;
  assign N3020 = T358[4] | T358[5];
  assign N3021 = T358[3] | N3020;
  assign N3022 = T358[2] | N3021;
  assign N3023 = T358[1] | N3022;
  assign N3024 = T358[0] | N3023;
  assign idxPagesOH_17 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T372;
  assign tgtPagesOH_11 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T864;
  assign N3025 = T354[4] | T354[5];
  assign N3026 = T354[3] | N3025;
  assign N3027 = T354[2] | N3026;
  assign N3028 = T354[1] | N3027;
  assign N3029 = T354[0] | N3028;
  assign idxPagesOH_16 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T368;
  assign tgtPagesOH_10 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T859;
  assign N3030 = T349[4] | T349[5];
  assign N3031 = T349[3] | N3030;
  assign N3032 = T349[2] | N3031;
  assign N3033 = T349[1] | N3032;
  assign N3034 = T349[0] | N3033;
  assign idxPagesOH_15 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T360;
  assign tgtPagesOH_9 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T853;
  assign N3035 = T345[4] | T345[5];
  assign N3036 = T345[3] | N3035;
  assign N3037 = T345[2] | N3036;
  assign N3038 = T345[1] | N3037;
  assign N3039 = T345[0] | N3038;
  assign idxPagesOH_14 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T356;
  assign tgtPagesOH_8 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T848;
  assign N3040 = T339[4] | T339[5];
  assign N3041 = T339[3] | N3040;
  assign N3042 = T339[2] | N3041;
  assign N3043 = T339[1] | N3042;
  assign N3044 = T339[0] | N3043;
  assign idxPagesOH_13 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T351;
  assign tgtPagesOH_7 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T840;
  assign N3045 = T335[4] | T335[5];
  assign N3046 = T335[3] | N3045;
  assign N3047 = T335[2] | N3046;
  assign N3048 = T335[1] | N3047;
  assign N3049 = T335[0] | N3048;
  assign idxPagesOH_12 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T347;
  assign tgtPagesOH_6 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T835;
  assign N3050 = T330[4] | T330[5];
  assign N3051 = T330[3] | N3050;
  assign N3052 = T330[2] | N3051;
  assign N3053 = T330[1] | N3052;
  assign N3054 = T330[0] | N3053;
  assign idxPagesOH_11 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T341;
  assign tgtPagesOH_5 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T829;
  assign N3055 = T326[4] | T326[5];
  assign N3056 = T326[3] | N3055;
  assign N3057 = T326[2] | N3056;
  assign N3058 = T326[1] | N3057;
  assign N3059 = T326[0] | N3058;
  assign idxPagesOH_10 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T337;
  assign tgtPagesOH_4 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T824;
  assign N3060 = T319[4] | T319[5];
  assign N3061 = T319[3] | N3060;
  assign N3062 = T319[2] | N3061;
  assign N3063 = T319[1] | N3062;
  assign N3064 = T319[0] | N3063;
  assign idxPagesOH_9 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T332;
  assign tgtPagesOH_3 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T817;
  assign N3065 = T315[4] | T315[5];
  assign N3066 = T315[3] | N3065;
  assign N3067 = T315[2] | N3066;
  assign N3068 = T315[1] | N3067;
  assign N3069 = T315[0] | N3068;
  assign idxPagesOH_8 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T328;
  assign tgtPagesOH_2 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T812;
  assign N3070 = T310[4] | T310[5];
  assign N3071 = T310[3] | N3070;
  assign N3072 = T310[2] | N3071;
  assign N3073 = T310[1] | N3072;
  assign N3074 = T310[0] | N3073;
  assign idxPagesOH_7 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T321;
  assign tgtPagesOH_0 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T797;
  assign tgtPagesOH_1 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T806;
  assign N3075 = T306[4] | T306[5];
  assign N3076 = T306[3] | N3075;
  assign N3077 = T306[2] | N3076;
  assign N3078 = T306[1] | N3077;
  assign N3079 = T306[0] | N3078;
  assign idxPagesOH_6 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T317;
  assign N3080 = T300[4] | T300[5];
  assign N3081 = T300[3] | N3080;
  assign N3082 = T300[2] | N3081;
  assign N3083 = T300[1] | N3082;
  assign N3084 = T300[0] | N3083;
  assign idxPagesOH_5 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T312;
  assign N3085 = T296[4] | T296[5];
  assign N3086 = T296[3] | N3085;
  assign N3087 = T296[2] | N3086;
  assign N3088 = T296[1] | N3087;
  assign N3089 = T296[0] | N3088;
  assign idxPagesOH_4 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T308;
  assign N3090 = T189[4] | T189[5];
  assign N3091 = T189[3] | N3090;
  assign N3092 = T189[2] | N3091;
  assign N3093 = T189[1] | N3092;
  assign N3094 = T189[0] | N3093;
  assign N3095 = T291[4] | T291[5];
  assign N3096 = T291[3] | N3095;
  assign N3097 = T291[2] | N3096;
  assign N3098 = T291[1] | N3097;
  assign N3099 = T291[0] | N3098;
  assign idxPagesOH_3 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T302;
  assign idxPagesOH_2 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T298;
  assign idxPagesOH_0 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T286;
  assign idxPagesOH_1 = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << T293;
  assign T173 = nextRepl + 1'b1;
  assign T201 = R198 + 1'b1;
  assign T2001 = T2027 ^ 1'b1;
  assign T2006 = T2027 ^ 1'b1;
  assign T2014 = R2010 + 1'b1;
  assign T2017 = R2010 - 1'b1;
  assign N3100 = ~T22[6];
  assign N3101 = T22[4] & T22[5];
  assign N3102 = N0 & T22[5];
  assign N0 = ~T22[4];
  assign N3103 = T22[4] & N1;
  assign N1 = ~T22[5];
  assign N3104 = N2 & N3;
  assign N2 = ~T22[4];
  assign N3 = ~T22[5];
  assign N3105 = T22[6] & N3101;
  assign N3106 = T22[6] & N3102;
  assign N3107 = T22[6] & N3103;
  assign N3108 = T22[6] & N3104;
  assign N3109 = N3100 & N3101;
  assign N3110 = N3100 & N3102;
  assign N3111 = N3100 & N3103;
  assign N3112 = N3100 & N3104;
  assign N3113 = T22[2] & T22[3];
  assign N3114 = N4 & T22[3];
  assign N4 = ~T22[2];
  assign N3115 = T22[2] & N5;
  assign N5 = ~T22[3];
  assign N3116 = N6 & N7;
  assign N6 = ~T22[2];
  assign N7 = ~T22[3];
  assign N3117 = T22[0] & T22[1];
  assign N3118 = N8 & T22[1];
  assign N8 = ~T22[0];
  assign N3119 = T22[0] & N9;
  assign N9 = ~T22[1];
  assign N3120 = N10 & N11;
  assign N10 = ~T22[0];
  assign N11 = ~T22[1];
  assign N3121 = N3113 & N3117;
  assign N3122 = N3113 & N3118;
  assign N3123 = N3113 & N3119;
  assign N3124 = N3113 & N3120;
  assign N3125 = N3114 & N3117;
  assign N3126 = N3114 & N3118;
  assign N3127 = N3114 & N3119;
  assign N3128 = N3114 & N3120;
  assign N3129 = N3115 & N3117;
  assign N3130 = N3115 & N3118;
  assign N3131 = N3115 & N3119;
  assign N3132 = N3115 & N3120;
  assign N3133 = N3116 & N3117;
  assign N3134 = N3116 & N3118;
  assign N3135 = N3116 & N3119;
  assign N3136 = N3116 & N3120;
  assign N1213 = N3105 & N3121;
  assign N1212 = N3105 & N3122;
  assign N1211 = N3105 & N3123;
  assign N1210 = N3105 & N3124;
  assign N1209 = N3105 & N3125;
  assign N1208 = N3105 & N3126;
  assign N1207 = N3105 & N3127;
  assign N1206 = N3105 & N3128;
  assign N1205 = N3105 & N3129;
  assign N1204 = N3105 & N3130;
  assign N1203 = N3105 & N3131;
  assign N1202 = N3105 & N3132;
  assign N1201 = N3105 & N3133;
  assign N1200 = N3105 & N3134;
  assign N1199 = N3105 & N3135;
  assign N1198 = N3105 & N3136;
  assign N1197 = N3106 & N3121;
  assign N1196 = N3106 & N3122;
  assign N1195 = N3106 & N3123;
  assign N1194 = N3106 & N3124;
  assign N1193 = N3106 & N3125;
  assign N1192 = N3106 & N3126;
  assign N1191 = N3106 & N3127;
  assign N1190 = N3106 & N3128;
  assign N1189 = N3106 & N3129;
  assign N1188 = N3106 & N3130;
  assign N1187 = N3106 & N3131;
  assign N1186 = N3106 & N3132;
  assign N1185 = N3106 & N3133;
  assign N1184 = N3106 & N3134;
  assign N1183 = N3106 & N3135;
  assign N1182 = N3106 & N3136;
  assign N1181 = N3107 & N3121;
  assign N1180 = N3107 & N3122;
  assign N1179 = N3107 & N3123;
  assign N1178 = N3107 & N3124;
  assign N1177 = N3107 & N3125;
  assign N1176 = N3107 & N3126;
  assign N1175 = N3107 & N3127;
  assign N1174 = N3107 & N3128;
  assign N1173 = N3107 & N3129;
  assign N1172 = N3107 & N3130;
  assign N1171 = N3107 & N3131;
  assign N1170 = N3107 & N3132;
  assign N1169 = N3107 & N3133;
  assign N1168 = N3107 & N3134;
  assign N1167 = N3107 & N3135;
  assign N1166 = N3107 & N3136;
  assign N1165 = N3108 & N3121;
  assign N1164 = N3108 & N3122;
  assign N1163 = N3108 & N3123;
  assign N1162 = N3108 & N3124;
  assign N1161 = N3108 & N3125;
  assign N1160 = N3108 & N3126;
  assign N1159 = N3108 & N3127;
  assign N1158 = N3108 & N3128;
  assign N1157 = N3108 & N3129;
  assign N1156 = N3108 & N3130;
  assign N1155 = N3108 & N3131;
  assign N1154 = N3108 & N3132;
  assign N1153 = N3108 & N3133;
  assign N1152 = N3108 & N3134;
  assign N1151 = N3108 & N3135;
  assign N1150 = N3108 & N3136;
  assign N1149 = N3109 & N3121;
  assign N1148 = N3109 & N3122;
  assign N1147 = N3109 & N3123;
  assign N1146 = N3109 & N3124;
  assign N1145 = N3109 & N3125;
  assign N1144 = N3109 & N3126;
  assign N1143 = N3109 & N3127;
  assign N1142 = N3109 & N3128;
  assign N1141 = N3109 & N3129;
  assign N1140 = N3109 & N3130;
  assign N1139 = N3109 & N3131;
  assign N1138 = N3109 & N3132;
  assign N1137 = N3109 & N3133;
  assign N1136 = N3109 & N3134;
  assign N1135 = N3109 & N3135;
  assign N1134 = N3109 & N3136;
  assign N1133 = N3110 & N3121;
  assign N1132 = N3110 & N3122;
  assign N1131 = N3110 & N3123;
  assign N1130 = N3110 & N3124;
  assign N1129 = N3110 & N3125;
  assign N1128 = N3110 & N3126;
  assign N1127 = N3110 & N3127;
  assign N1126 = N3110 & N3128;
  assign N1125 = N3110 & N3129;
  assign N1124 = N3110 & N3130;
  assign N1123 = N3110 & N3131;
  assign N1122 = N3110 & N3132;
  assign N1121 = N3110 & N3133;
  assign N1120 = N3110 & N3134;
  assign N1119 = N3110 & N3135;
  assign N1118 = N3110 & N3136;
  assign N1117 = N3111 & N3121;
  assign N1116 = N3111 & N3122;
  assign N1115 = N3111 & N3123;
  assign N1114 = N3111 & N3124;
  assign N1113 = N3111 & N3125;
  assign N1112 = N3111 & N3126;
  assign N1111 = N3111 & N3127;
  assign N1110 = N3111 & N3128;
  assign N1109 = N3111 & N3129;
  assign N1108 = N3111 & N3130;
  assign N1107 = N3111 & N3131;
  assign N1106 = N3111 & N3132;
  assign N1105 = N3111 & N3133;
  assign N1104 = N3111 & N3134;
  assign N1103 = N3111 & N3135;
  assign N1102 = N3111 & N3136;
  assign N1101 = N3112 & N3121;
  assign N1100 = N3112 & N3122;
  assign N1099 = N3112 & N3123;
  assign N1098 = N3112 & N3124;
  assign N1097 = N3112 & N3125;
  assign N1096 = N3112 & N3126;
  assign N1095 = N3112 & N3127;
  assign N1094 = N3112 & N3128;
  assign N1093 = N3112 & N3129;
  assign N1092 = N3112 & N3130;
  assign N1091 = N3112 & N3131;
  assign N1090 = N3112 & N3132;
  assign N1089 = N3112 & N3133;
  assign N1088 = N3112 & N3134;
  assign N1087 = N3112 & N3135;
  assign N1086 = N3112 & N3136;
  assign N3137 = ~T169[5];
  assign N3138 = T169[3] & T169[4];
  assign N3139 = N12 & T169[4];
  assign N12 = ~T169[3];
  assign N3140 = T169[3] & N13;
  assign N13 = ~T169[4];
  assign N3141 = N14 & N15;
  assign N14 = ~T169[3];
  assign N15 = ~T169[4];
  assign N3142 = T169[5] & N3138;
  assign N3143 = T169[5] & N3139;
  assign N3144 = T169[5] & N3140;
  assign N3145 = T169[5] & N3141;
  assign N3146 = N3137 & N3138;
  assign N3147 = N3137 & N3139;
  assign N3148 = N3137 & N3140;
  assign N3149 = N3137 & N3141;
  assign N3150 = ~T169[2];
  assign N3151 = T169[0] & T169[1];
  assign N3152 = N16 & T169[1];
  assign N16 = ~T169[0];
  assign N3153 = T169[0] & N17;
  assign N17 = ~T169[1];
  assign N3154 = N18 & N19;
  assign N18 = ~T169[0];
  assign N19 = ~T169[1];
  assign N3155 = T169[2] & N3151;
  assign N3156 = T169[2] & N3152;
  assign N3157 = T169[2] & N3153;
  assign N3158 = T169[2] & N3154;
  assign N3159 = N3150 & N3151;
  assign N3160 = N3150 & N3152;
  assign N3161 = N3150 & N3153;
  assign N3162 = N3150 & N3154;
  assign N1733 = N3142 & N3157;
  assign N1732 = N3142 & N3158;
  assign N1731 = N3142 & N3159;
  assign N1730 = N3142 & N3160;
  assign N1729 = N3142 & N3161;
  assign N1728 = N3142 & N3162;
  assign N1727 = N3143 & N3155;
  assign N1726 = N3143 & N3156;
  assign N1725 = N3143 & N3157;
  assign N1724 = N3143 & N3158;
  assign N1723 = N3143 & N3159;
  assign N1722 = N3143 & N3160;
  assign N1721 = N3143 & N3161;
  assign N1720 = N3143 & N3162;
  assign N1719 = N3144 & N3155;
  assign N1718 = N3144 & N3156;
  assign N1717 = N3144 & N3157;
  assign N1716 = N3144 & N3158;
  assign N1715 = N3144 & N3159;
  assign N1714 = N3144 & N3160;
  assign N1713 = N3144 & N3161;
  assign N1712 = N3144 & N3162;
  assign N1711 = N3145 & N3155;
  assign N1710 = N3145 & N3156;
  assign N1709 = N3145 & N3157;
  assign N1708 = N3145 & N3158;
  assign N1707 = N3145 & N3159;
  assign N1706 = N3145 & N3160;
  assign N1705 = N3145 & N3161;
  assign N1704 = N3145 & N3162;
  assign N1703 = N3146 & N3155;
  assign N1702 = N3146 & N3156;
  assign N1701 = N3146 & N3157;
  assign N1700 = N3146 & N3158;
  assign N1699 = N3146 & N3159;
  assign N1698 = N3146 & N3160;
  assign N1697 = N3146 & N3161;
  assign N1696 = N3146 & N3162;
  assign N1695 = N3147 & N3155;
  assign N1694 = N3147 & N3156;
  assign N1693 = N3147 & N3157;
  assign N1692 = N3147 & N3158;
  assign N1691 = N3147 & N3159;
  assign N1690 = N3147 & N3160;
  assign N1689 = N3147 & N3161;
  assign N1688 = N3147 & N3162;
  assign N1687 = N3148 & N3155;
  assign N1686 = N3148 & N3156;
  assign N1685 = N3148 & N3157;
  assign N1684 = N3148 & N3158;
  assign N1683 = N3148 & N3159;
  assign N1682 = N3148 & N3160;
  assign N1681 = N3148 & N3161;
  assign N1680 = N3148 & N3162;
  assign N1679 = N3149 & N3155;
  assign N1678 = N3149 & N3156;
  assign N1677 = N3149 & N3157;
  assign N1676 = N3149 & N3158;
  assign N1675 = N3149 & N3159;
  assign N1674 = N3149 & N3160;
  assign N1673 = N3149 & N3161;
  assign N1672 = N3149 & N3162;
  assign N3163 = T169[3] & T169[4];
  assign N3164 = N20 & T169[4];
  assign N20 = ~T169[3];
  assign N3165 = T169[3] & N21;
  assign N21 = ~T169[4];
  assign N3166 = N22 & N23;
  assign N22 = ~T169[3];
  assign N23 = ~T169[4];
  assign N3167 = T169[5] & N3163;
  assign N3168 = T169[5] & N3164;
  assign N3169 = T169[5] & N3165;
  assign N3170 = T169[5] & N3166;
  assign N3171 = N3137 & N3163;
  assign N3172 = N3137 & N3164;
  assign N3173 = N3137 & N3165;
  assign N3174 = N3137 & N3166;
  assign N3175 = T169[0] & T169[1];
  assign N3176 = N24 & T169[1];
  assign N24 = ~T169[0];
  assign N3177 = T169[0] & N25;
  assign N25 = ~T169[1];
  assign N3178 = N26 & N27;
  assign N26 = ~T169[0];
  assign N27 = ~T169[1];
  assign N3179 = T169[2] & N3175;
  assign N3180 = T169[2] & N3176;
  assign N3181 = T169[2] & N3177;
  assign N3182 = T169[2] & N3178;
  assign N3183 = N3150 & N3175;
  assign N3184 = N3150 & N3176;
  assign N3185 = N3150 & N3177;
  assign N3186 = N3150 & N3178;
  assign N1858 = N3167 & N3181;
  assign N1857 = N3167 & N3182;
  assign N1856 = N3167 & N3183;
  assign N1855 = N3167 & N3184;
  assign N1854 = N3167 & N3185;
  assign N1853 = N3167 & N3186;
  assign N1852 = N3168 & N3179;
  assign N1851 = N3168 & N3180;
  assign N1850 = N3168 & N3181;
  assign N1849 = N3168 & N3182;
  assign N1848 = N3168 & N3183;
  assign N1847 = N3168 & N3184;
  assign N1846 = N3168 & N3185;
  assign N1845 = N3168 & N3186;
  assign N1844 = N3169 & N3179;
  assign N1843 = N3169 & N3180;
  assign N1842 = N3169 & N3181;
  assign N1841 = N3169 & N3182;
  assign N1840 = N3169 & N3183;
  assign N1839 = N3169 & N3184;
  assign N1838 = N3169 & N3185;
  assign N1837 = N3169 & N3186;
  assign N1836 = N3170 & N3179;
  assign N1835 = N3170 & N3180;
  assign N1834 = N3170 & N3181;
  assign N1833 = N3170 & N3182;
  assign N1832 = N3170 & N3183;
  assign N1831 = N3170 & N3184;
  assign N1830 = N3170 & N3185;
  assign N1829 = N3170 & N3186;
  assign N1828 = N3171 & N3179;
  assign N1827 = N3171 & N3180;
  assign N1826 = N3171 & N3181;
  assign N1825 = N3171 & N3182;
  assign N1824 = N3171 & N3183;
  assign N1823 = N3171 & N3184;
  assign N1822 = N3171 & N3185;
  assign N1821 = N3171 & N3186;
  assign N1820 = N3172 & N3179;
  assign N1819 = N3172 & N3180;
  assign N1818 = N3172 & N3181;
  assign N1817 = N3172 & N3182;
  assign N1816 = N3172 & N3183;
  assign N1815 = N3172 & N3184;
  assign N1814 = N3172 & N3185;
  assign N1813 = N3172 & N3186;
  assign N1812 = N3173 & N3179;
  assign N1811 = N3173 & N3180;
  assign N1810 = N3173 & N3181;
  assign N1809 = N3173 & N3182;
  assign N1808 = N3173 & N3183;
  assign N1807 = N3173 & N3184;
  assign N1806 = N3173 & N3185;
  assign N1805 = N3173 & N3186;
  assign N1804 = N3174 & N3179;
  assign N1803 = N3174 & N3180;
  assign N1802 = N3174 & N3181;
  assign N1801 = N3174 & N3182;
  assign N1800 = N3174 & N3183;
  assign N1799 = N3174 & N3184;
  assign N1798 = N3174 & N3185;
  assign N1797 = N3174 & N3186;
  assign N3187 = T169[3] & T169[4];
  assign N3188 = N28 & T169[4];
  assign N28 = ~T169[3];
  assign N3189 = T169[3] & N29;
  assign N29 = ~T169[4];
  assign N3190 = N30 & N31;
  assign N30 = ~T169[3];
  assign N31 = ~T169[4];
  assign N3191 = T169[5] & N3187;
  assign N3192 = T169[5] & N3188;
  assign N3193 = T169[5] & N3189;
  assign N3194 = T169[5] & N3190;
  assign N3195 = N3137 & N3187;
  assign N3196 = N3137 & N3188;
  assign N3197 = N3137 & N3189;
  assign N3198 = N3137 & N3190;
  assign N3199 = T169[0] & T169[1];
  assign N3200 = N32 & T169[1];
  assign N32 = ~T169[0];
  assign N3201 = T169[0] & N33;
  assign N33 = ~T169[1];
  assign N3202 = N34 & N35;
  assign N34 = ~T169[0];
  assign N35 = ~T169[1];
  assign N3203 = T169[2] & N3199;
  assign N3204 = T169[2] & N3200;
  assign N3205 = T169[2] & N3201;
  assign N3206 = T169[2] & N3202;
  assign N3207 = N3150 & N3199;
  assign N3208 = N3150 & N3200;
  assign N3209 = N3150 & N3201;
  assign N3210 = N3150 & N3202;
  assign N1983 = N3191 & N3205;
  assign N1982 = N3191 & N3206;
  assign N1981 = N3191 & N3207;
  assign N1980 = N3191 & N3208;
  assign N1979 = N3191 & N3209;
  assign N1978 = N3191 & N3210;
  assign N1977 = N3192 & N3203;
  assign N1976 = N3192 & N3204;
  assign N1975 = N3192 & N3205;
  assign N1974 = N3192 & N3206;
  assign N1973 = N3192 & N3207;
  assign N1972 = N3192 & N3208;
  assign N1971 = N3192 & N3209;
  assign N1970 = N3192 & N3210;
  assign N1969 = N3193 & N3203;
  assign N1968 = N3193 & N3204;
  assign N1967 = N3193 & N3205;
  assign N1966 = N3193 & N3206;
  assign N1965 = N3193 & N3207;
  assign N1964 = N3193 & N3208;
  assign N1963 = N3193 & N3209;
  assign N1962 = N3193 & N3210;
  assign N1961 = N3194 & N3203;
  assign N1960 = N3194 & N3204;
  assign N1959 = N3194 & N3205;
  assign N1958 = N3194 & N3206;
  assign N1957 = N3194 & N3207;
  assign N1956 = N3194 & N3208;
  assign N1955 = N3194 & N3209;
  assign N1954 = N3194 & N3210;
  assign N1953 = N3195 & N3203;
  assign N1952 = N3195 & N3204;
  assign N1951 = N3195 & N3205;
  assign N1950 = N3195 & N3206;
  assign N1949 = N3195 & N3207;
  assign N1948 = N3195 & N3208;
  assign N1947 = N3195 & N3209;
  assign N1946 = N3195 & N3210;
  assign N1945 = N3196 & N3203;
  assign N1944 = N3196 & N3204;
  assign N1943 = N3196 & N3205;
  assign N1942 = N3196 & N3206;
  assign N1941 = N3196 & N3207;
  assign N1940 = N3196 & N3208;
  assign N1939 = N3196 & N3209;
  assign N1938 = N3196 & N3210;
  assign N1937 = N3197 & N3203;
  assign N1936 = N3197 & N3204;
  assign N1935 = N3197 & N3205;
  assign N1934 = N3197 & N3206;
  assign N1933 = N3197 & N3207;
  assign N1932 = N3197 & N3208;
  assign N1931 = N3197 & N3209;
  assign N1930 = N3197 & N3210;
  assign N1929 = N3198 & N3203;
  assign N1928 = N3198 & N3204;
  assign N1927 = N3198 & N3205;
  assign N1926 = N3198 & N3206;
  assign N1925 = N3198 & N3207;
  assign N1924 = N3198 & N3208;
  assign N1923 = N3198 & N3209;
  assign N1922 = N3198 & N3210;
  assign N3211 = T169[3] & T169[4];
  assign N3212 = N36 & T169[4];
  assign N36 = ~T169[3];
  assign N3213 = T169[3] & N37;
  assign N37 = ~T169[4];
  assign N3214 = N38 & N39;
  assign N38 = ~T169[3];
  assign N39 = ~T169[4];
  assign N3215 = T169[5] & N3211;
  assign N3216 = T169[5] & N3212;
  assign N3217 = T169[5] & N3213;
  assign N3218 = T169[5] & N3214;
  assign N3219 = N3137 & N3211;
  assign N3220 = N3137 & N3212;
  assign N3221 = N3137 & N3213;
  assign N3222 = N3137 & N3214;
  assign N3223 = T169[0] & T169[1];
  assign N3224 = N40 & T169[1];
  assign N40 = ~T169[0];
  assign N3225 = T169[0] & N41;
  assign N41 = ~T169[1];
  assign N3226 = N42 & N43;
  assign N42 = ~T169[0];
  assign N43 = ~T169[1];
  assign N3227 = T169[2] & N3223;
  assign N3228 = T169[2] & N3224;
  assign N3229 = T169[2] & N3225;
  assign N3230 = T169[2] & N3226;
  assign N3231 = N3150 & N3223;
  assign N3232 = N3150 & N3224;
  assign N3233 = N3150 & N3225;
  assign N3234 = N3150 & N3226;
  assign N2108 = N3215 & N3229;
  assign N2107 = N3215 & N3230;
  assign N2106 = N3215 & N3231;
  assign N2105 = N3215 & N3232;
  assign N2104 = N3215 & N3233;
  assign N2103 = N3215 & N3234;
  assign N2102 = N3216 & N3227;
  assign N2101 = N3216 & N3228;
  assign N2100 = N3216 & N3229;
  assign N2099 = N3216 & N3230;
  assign N2098 = N3216 & N3231;
  assign N2097 = N3216 & N3232;
  assign N2096 = N3216 & N3233;
  assign N2095 = N3216 & N3234;
  assign N2094 = N3217 & N3227;
  assign N2093 = N3217 & N3228;
  assign N2092 = N3217 & N3229;
  assign N2091 = N3217 & N3230;
  assign N2090 = N3217 & N3231;
  assign N2089 = N3217 & N3232;
  assign N2088 = N3217 & N3233;
  assign N2087 = N3217 & N3234;
  assign N2086 = N3218 & N3227;
  assign N2085 = N3218 & N3228;
  assign N2084 = N3218 & N3229;
  assign N2083 = N3218 & N3230;
  assign N2082 = N3218 & N3231;
  assign N2081 = N3218 & N3232;
  assign N2080 = N3218 & N3233;
  assign N2079 = N3218 & N3234;
  assign N2078 = N3219 & N3227;
  assign N2077 = N3219 & N3228;
  assign N2076 = N3219 & N3229;
  assign N2075 = N3219 & N3230;
  assign N2074 = N3219 & N3231;
  assign N2073 = N3219 & N3232;
  assign N2072 = N3219 & N3233;
  assign N2071 = N3219 & N3234;
  assign N2070 = N3220 & N3227;
  assign N2069 = N3220 & N3228;
  assign N2068 = N3220 & N3229;
  assign N2067 = N3220 & N3230;
  assign N2066 = N3220 & N3231;
  assign N2065 = N3220 & N3232;
  assign N2064 = N3220 & N3233;
  assign N2063 = N3220 & N3234;
  assign N2062 = N3221 & N3227;
  assign N2061 = N3221 & N3228;
  assign N2060 = N3221 & N3229;
  assign N2059 = N3221 & N3230;
  assign N2058 = N3221 & N3231;
  assign N2057 = N3221 & N3232;
  assign N2056 = N3221 & N3233;
  assign N2055 = N3221 & N3234;
  assign N2054 = N3222 & N3227;
  assign N2053 = N3222 & N3228;
  assign N2052 = N3222 & N3229;
  assign N2051 = N3222 & N3230;
  assign N2050 = N3222 & N3231;
  assign N2049 = N3222 & N3232;
  assign N2048 = N3222 & N3233;
  assign N2047 = N3222 & N3234;
  assign N3235 = T169[3] & T169[4];
  assign N3236 = N44 & T169[4];
  assign N44 = ~T169[3];
  assign N3237 = T169[3] & N45;
  assign N45 = ~T169[4];
  assign N3238 = N46 & N47;
  assign N46 = ~T169[3];
  assign N47 = ~T169[4];
  assign N3239 = T169[5] & N3235;
  assign N3240 = T169[5] & N3236;
  assign N3241 = T169[5] & N3237;
  assign N3242 = T169[5] & N3238;
  assign N3243 = N3137 & N3235;
  assign N3244 = N3137 & N3236;
  assign N3245 = N3137 & N3237;
  assign N3246 = N3137 & N3238;
  assign N3247 = T169[0] & T169[1];
  assign N3248 = N48 & T169[1];
  assign N48 = ~T169[0];
  assign N3249 = T169[0] & N49;
  assign N49 = ~T169[1];
  assign N3250 = N50 & N51;
  assign N50 = ~T169[0];
  assign N51 = ~T169[1];
  assign N3251 = T169[2] & N3247;
  assign N3252 = T169[2] & N3248;
  assign N3253 = T169[2] & N3249;
  assign N3254 = T169[2] & N3250;
  assign N3255 = N3150 & N3247;
  assign N3256 = N3150 & N3248;
  assign N3257 = N3150 & N3249;
  assign N3258 = N3150 & N3250;
  assign N2244 = N3239 & N3253;
  assign N2243 = N3239 & N3254;
  assign N2242 = N3239 & N3255;
  assign N2241 = N3239 & N3256;
  assign N2240 = N3239 & N3257;
  assign N2239 = N3239 & N3258;
  assign N2238 = N3240 & N3251;
  assign N2237 = N3240 & N3252;
  assign N2236 = N3240 & N3253;
  assign N2235 = N3240 & N3254;
  assign N2234 = N3240 & N3255;
  assign N2233 = N3240 & N3256;
  assign N2232 = N3240 & N3257;
  assign N2231 = N3240 & N3258;
  assign N2230 = N3241 & N3251;
  assign N2229 = N3241 & N3252;
  assign N2228 = N3241 & N3253;
  assign N2227 = N3241 & N3254;
  assign N2226 = N3241 & N3255;
  assign N2225 = N3241 & N3256;
  assign N2224 = N3241 & N3257;
  assign N2223 = N3241 & N3258;
  assign N2222 = N3242 & N3251;
  assign N2221 = N3242 & N3252;
  assign N2220 = N3242 & N3253;
  assign N2219 = N3242 & N3254;
  assign N2218 = N3242 & N3255;
  assign N2217 = N3242 & N3256;
  assign N2216 = N3242 & N3257;
  assign N2215 = N3242 & N3258;
  assign N2214 = N3243 & N3251;
  assign N2213 = N3243 & N3252;
  assign N2212 = N3243 & N3253;
  assign N2211 = N3243 & N3254;
  assign N2210 = N3243 & N3255;
  assign N2209 = N3243 & N3256;
  assign N2208 = N3243 & N3257;
  assign N2207 = N3243 & N3258;
  assign N2206 = N3244 & N3251;
  assign N2205 = N3244 & N3252;
  assign N2204 = N3244 & N3253;
  assign N2203 = N3244 & N3254;
  assign N2202 = N3244 & N3255;
  assign N2201 = N3244 & N3256;
  assign N2200 = N3244 & N3257;
  assign N2199 = N3244 & N3258;
  assign N2198 = N3245 & N3251;
  assign N2197 = N3245 & N3252;
  assign N2196 = N3245 & N3253;
  assign N2195 = N3245 & N3254;
  assign N2194 = N3245 & N3255;
  assign N2193 = N3245 & N3256;
  assign N2192 = N3245 & N3257;
  assign N2191 = N3245 & N3258;
  assign N2190 = N3246 & N3251;
  assign N2189 = N3246 & N3252;
  assign N2188 = N3246 & N3253;
  assign N2187 = N3246 & N3254;
  assign N2186 = N3246 & N3255;
  assign N2185 = N3246 & N3256;
  assign N2184 = N3246 & N3257;
  assign N2183 = N3246 & N3258;
  assign N52 = N56 & N57;
  assign N53 = N52 & N58;
  assign N54 = N53 & N59;
  assign N55 = N54 & N60;
  assign N1020 = N55 & N61;
  assign N56 = ~io_resp_bits_entry[5];
  assign N57 = ~io_resp_bits_entry[4];
  assign N58 = ~io_resp_bits_entry[3];
  assign N59 = ~io_resp_bits_entry[2];
  assign N60 = ~io_resp_bits_entry[0];
  assign N61 = ~io_resp_bits_entry[1];
  assign N62 = io_resp_bits_entry[5] & N66;
  assign N63 = N62 & N67;
  assign N64 = N63 & N68;
  assign N65 = N64 & N69;
  assign N1021 = N65 & N70;
  assign N66 = ~io_resp_bits_entry[4];
  assign N67 = ~io_resp_bits_entry[3];
  assign N68 = ~io_resp_bits_entry[2];
  assign N69 = ~io_resp_bits_entry[0];
  assign N70 = ~io_resp_bits_entry[1];
  assign N71 = N75 & N76;
  assign N72 = N71 & N77;
  assign N73 = N72 & N78;
  assign N74 = N73 & io_resp_bits_entry[0];
  assign N1022 = N74 & N79;
  assign N75 = ~io_resp_bits_entry[5];
  assign N76 = ~io_resp_bits_entry[4];
  assign N77 = ~io_resp_bits_entry[3];
  assign N78 = ~io_resp_bits_entry[2];
  assign N79 = ~io_resp_bits_entry[1];
  assign N80 = N84 & N85;
  assign N81 = N80 & N86;
  assign N82 = N81 & N87;
  assign N83 = N82 & N88;
  assign N1024 = N83 & io_resp_bits_entry[1];
  assign N84 = ~io_resp_bits_entry[5];
  assign N85 = ~io_resp_bits_entry[4];
  assign N86 = ~io_resp_bits_entry[3];
  assign N87 = ~io_resp_bits_entry[2];
  assign N88 = ~io_resp_bits_entry[0];
  assign N89 = N93 & N94;
  assign N90 = N89 & N95;
  assign N91 = N90 & N96;
  assign N92 = N91 & io_resp_bits_entry[0];
  assign N1026 = N92 & io_resp_bits_entry[1];
  assign N93 = ~io_resp_bits_entry[5];
  assign N94 = ~io_resp_bits_entry[4];
  assign N95 = ~io_resp_bits_entry[3];
  assign N96 = ~io_resp_bits_entry[2];
  assign N97 = N101 & N102;
  assign N98 = N97 & N103;
  assign N99 = N98 & io_resp_bits_entry[2];
  assign N100 = N99 & N104;
  assign N1028 = N100 & N105;
  assign N101 = ~io_resp_bits_entry[5];
  assign N102 = ~io_resp_bits_entry[4];
  assign N103 = ~io_resp_bits_entry[3];
  assign N104 = ~io_resp_bits_entry[0];
  assign N105 = ~io_resp_bits_entry[1];
  assign N106 = N110 & N111;
  assign N107 = N106 & N112;
  assign N108 = N107 & io_resp_bits_entry[2];
  assign N109 = N108 & io_resp_bits_entry[0];
  assign N1030 = N109 & N113;
  assign N110 = ~io_resp_bits_entry[5];
  assign N111 = ~io_resp_bits_entry[4];
  assign N112 = ~io_resp_bits_entry[3];
  assign N113 = ~io_resp_bits_entry[1];
  assign N114 = N118 & N119;
  assign N115 = N114 & N120;
  assign N116 = N115 & io_resp_bits_entry[2];
  assign N117 = N116 & N121;
  assign N1032 = N117 & io_resp_bits_entry[1];
  assign N118 = ~io_resp_bits_entry[5];
  assign N119 = ~io_resp_bits_entry[4];
  assign N120 = ~io_resp_bits_entry[3];
  assign N121 = ~io_resp_bits_entry[0];
  assign N122 = N126 & N127;
  assign N123 = N122 & N128;
  assign N124 = N123 & io_resp_bits_entry[2];
  assign N125 = N124 & io_resp_bits_entry[0];
  assign N1034 = N125 & io_resp_bits_entry[1];
  assign N126 = ~io_resp_bits_entry[5];
  assign N127 = ~io_resp_bits_entry[4];
  assign N128 = ~io_resp_bits_entry[3];
  assign N129 = N133 & N134;
  assign N130 = N129 & io_resp_bits_entry[3];
  assign N131 = N130 & N135;
  assign N132 = N131 & N136;
  assign N1036 = N132 & N137;
  assign N133 = ~io_resp_bits_entry[5];
  assign N134 = ~io_resp_bits_entry[4];
  assign N135 = ~io_resp_bits_entry[2];
  assign N136 = ~io_resp_bits_entry[0];
  assign N137 = ~io_resp_bits_entry[1];
  assign N138 = N142 & N143;
  assign N139 = N138 & io_resp_bits_entry[3];
  assign N140 = N139 & N144;
  assign N141 = N140 & io_resp_bits_entry[0];
  assign N1038 = N141 & N145;
  assign N142 = ~io_resp_bits_entry[5];
  assign N143 = ~io_resp_bits_entry[4];
  assign N144 = ~io_resp_bits_entry[2];
  assign N145 = ~io_resp_bits_entry[1];
  assign N146 = N150 & N151;
  assign N147 = N146 & io_resp_bits_entry[3];
  assign N148 = N147 & N152;
  assign N149 = N148 & N153;
  assign N1040 = N149 & io_resp_bits_entry[1];
  assign N150 = ~io_resp_bits_entry[5];
  assign N151 = ~io_resp_bits_entry[4];
  assign N152 = ~io_resp_bits_entry[2];
  assign N153 = ~io_resp_bits_entry[0];
  assign N154 = N158 & N159;
  assign N155 = N154 & io_resp_bits_entry[3];
  assign N156 = N155 & N160;
  assign N157 = N156 & io_resp_bits_entry[0];
  assign N1042 = N157 & io_resp_bits_entry[1];
  assign N158 = ~io_resp_bits_entry[5];
  assign N159 = ~io_resp_bits_entry[4];
  assign N160 = ~io_resp_bits_entry[2];
  assign N161 = N165 & N166;
  assign N162 = N161 & io_resp_bits_entry[3];
  assign N163 = N162 & io_resp_bits_entry[2];
  assign N164 = N163 & N167;
  assign N1044 = N164 & N168;
  assign N165 = ~io_resp_bits_entry[5];
  assign N166 = ~io_resp_bits_entry[4];
  assign N167 = ~io_resp_bits_entry[0];
  assign N168 = ~io_resp_bits_entry[1];
  assign N169 = N173 & N174;
  assign N170 = N169 & io_resp_bits_entry[3];
  assign N171 = N170 & io_resp_bits_entry[2];
  assign N172 = N171 & io_resp_bits_entry[0];
  assign N1046 = N172 & N175;
  assign N173 = ~io_resp_bits_entry[5];
  assign N174 = ~io_resp_bits_entry[4];
  assign N175 = ~io_resp_bits_entry[1];
  assign N176 = N180 & N181;
  assign N177 = N176 & io_resp_bits_entry[3];
  assign N178 = N177 & io_resp_bits_entry[2];
  assign N179 = N178 & N182;
  assign N1048 = N179 & io_resp_bits_entry[1];
  assign N180 = ~io_resp_bits_entry[5];
  assign N181 = ~io_resp_bits_entry[4];
  assign N182 = ~io_resp_bits_entry[0];
  assign N183 = N187 & N188;
  assign N184 = N183 & io_resp_bits_entry[3];
  assign N185 = N184 & io_resp_bits_entry[2];
  assign N186 = N185 & io_resp_bits_entry[0];
  assign N1050 = N186 & io_resp_bits_entry[1];
  assign N187 = ~io_resp_bits_entry[5];
  assign N188 = ~io_resp_bits_entry[4];
  assign N189 = N193 & io_resp_bits_entry[4];
  assign N190 = N189 & N194;
  assign N191 = N190 & N195;
  assign N192 = N191 & N196;
  assign N1052 = N192 & N197;
  assign N193 = ~io_resp_bits_entry[5];
  assign N194 = ~io_resp_bits_entry[3];
  assign N195 = ~io_resp_bits_entry[2];
  assign N196 = ~io_resp_bits_entry[0];
  assign N197 = ~io_resp_bits_entry[1];
  assign N198 = N202 & io_resp_bits_entry[4];
  assign N199 = N198 & N203;
  assign N200 = N199 & N204;
  assign N201 = N200 & io_resp_bits_entry[0];
  assign N1054 = N201 & N205;
  assign N202 = ~io_resp_bits_entry[5];
  assign N203 = ~io_resp_bits_entry[3];
  assign N204 = ~io_resp_bits_entry[2];
  assign N205 = ~io_resp_bits_entry[1];
  assign N206 = N210 & io_resp_bits_entry[4];
  assign N207 = N206 & N211;
  assign N208 = N207 & N212;
  assign N209 = N208 & N213;
  assign N1056 = N209 & io_resp_bits_entry[1];
  assign N210 = ~io_resp_bits_entry[5];
  assign N211 = ~io_resp_bits_entry[3];
  assign N212 = ~io_resp_bits_entry[2];
  assign N213 = ~io_resp_bits_entry[0];
  assign N214 = N218 & io_resp_bits_entry[4];
  assign N215 = N214 & N219;
  assign N216 = N215 & N220;
  assign N217 = N216 & io_resp_bits_entry[0];
  assign N1058 = N217 & io_resp_bits_entry[1];
  assign N218 = ~io_resp_bits_entry[5];
  assign N219 = ~io_resp_bits_entry[3];
  assign N220 = ~io_resp_bits_entry[2];
  assign N221 = N225 & io_resp_bits_entry[4];
  assign N222 = N221 & N226;
  assign N223 = N222 & io_resp_bits_entry[2];
  assign N224 = N223 & N227;
  assign N1060 = N224 & N228;
  assign N225 = ~io_resp_bits_entry[5];
  assign N226 = ~io_resp_bits_entry[3];
  assign N227 = ~io_resp_bits_entry[0];
  assign N228 = ~io_resp_bits_entry[1];
  assign N229 = N233 & io_resp_bits_entry[4];
  assign N230 = N229 & N234;
  assign N231 = N230 & io_resp_bits_entry[2];
  assign N232 = N231 & io_resp_bits_entry[0];
  assign N1062 = N232 & N235;
  assign N233 = ~io_resp_bits_entry[5];
  assign N234 = ~io_resp_bits_entry[3];
  assign N235 = ~io_resp_bits_entry[1];
  assign N236 = N240 & io_resp_bits_entry[4];
  assign N237 = N236 & N241;
  assign N238 = N237 & io_resp_bits_entry[2];
  assign N239 = N238 & N242;
  assign N1064 = N239 & io_resp_bits_entry[1];
  assign N240 = ~io_resp_bits_entry[5];
  assign N241 = ~io_resp_bits_entry[3];
  assign N242 = ~io_resp_bits_entry[0];
  assign N243 = N247 & io_resp_bits_entry[4];
  assign N244 = N243 & N248;
  assign N245 = N244 & io_resp_bits_entry[2];
  assign N246 = N245 & io_resp_bits_entry[0];
  assign N1066 = N246 & io_resp_bits_entry[1];
  assign N247 = ~io_resp_bits_entry[5];
  assign N248 = ~io_resp_bits_entry[3];
  assign N249 = N253 & io_resp_bits_entry[4];
  assign N250 = N249 & io_resp_bits_entry[3];
  assign N251 = N250 & N254;
  assign N252 = N251 & N255;
  assign N1068 = N252 & N256;
  assign N253 = ~io_resp_bits_entry[5];
  assign N254 = ~io_resp_bits_entry[2];
  assign N255 = ~io_resp_bits_entry[0];
  assign N256 = ~io_resp_bits_entry[1];
  assign N257 = N261 & io_resp_bits_entry[4];
  assign N258 = N257 & io_resp_bits_entry[3];
  assign N259 = N258 & N262;
  assign N260 = N259 & io_resp_bits_entry[0];
  assign N1070 = N260 & N263;
  assign N261 = ~io_resp_bits_entry[5];
  assign N262 = ~io_resp_bits_entry[2];
  assign N263 = ~io_resp_bits_entry[1];
  assign N264 = N268 & io_resp_bits_entry[4];
  assign N265 = N264 & io_resp_bits_entry[3];
  assign N266 = N265 & N269;
  assign N267 = N266 & N270;
  assign N1072 = N267 & io_resp_bits_entry[1];
  assign N268 = ~io_resp_bits_entry[5];
  assign N269 = ~io_resp_bits_entry[2];
  assign N270 = ~io_resp_bits_entry[0];
  assign N271 = N275 & io_resp_bits_entry[4];
  assign N272 = N271 & io_resp_bits_entry[3];
  assign N273 = N272 & N276;
  assign N274 = N273 & io_resp_bits_entry[0];
  assign N1074 = N274 & io_resp_bits_entry[1];
  assign N275 = ~io_resp_bits_entry[5];
  assign N276 = ~io_resp_bits_entry[2];
  assign N277 = N281 & io_resp_bits_entry[4];
  assign N278 = N277 & io_resp_bits_entry[3];
  assign N279 = N278 & io_resp_bits_entry[2];
  assign N280 = N279 & N282;
  assign N1076 = N280 & N283;
  assign N281 = ~io_resp_bits_entry[5];
  assign N282 = ~io_resp_bits_entry[0];
  assign N283 = ~io_resp_bits_entry[1];
  assign N284 = N288 & io_resp_bits_entry[4];
  assign N285 = N284 & io_resp_bits_entry[3];
  assign N286 = N285 & io_resp_bits_entry[2];
  assign N287 = N286 & io_resp_bits_entry[0];
  assign N1078 = N287 & N289;
  assign N288 = ~io_resp_bits_entry[5];
  assign N289 = ~io_resp_bits_entry[1];
  assign N1080 = io_resp_bits_entry[4] & io_resp_bits_entry[3] & (io_resp_bits_entry[2] & N290) & io_resp_bits_entry[1];
  assign N290 = ~io_resp_bits_entry[0];
  assign N1081 = io_resp_bits_entry[4] & io_resp_bits_entry[3] & (io_resp_bits_entry[2] & io_resp_bits_entry[0]) & io_resp_bits_entry[1];
  assign N291 = io_resp_bits_entry[5] & N295;
  assign N292 = N291 & N296;
  assign N293 = N292 & N297;
  assign N294 = N293 & io_resp_bits_entry[0];
  assign N1023 = N294 & N298;
  assign N295 = ~io_resp_bits_entry[4];
  assign N296 = ~io_resp_bits_entry[3];
  assign N297 = ~io_resp_bits_entry[2];
  assign N298 = ~io_resp_bits_entry[1];
  assign N299 = io_resp_bits_entry[5] & N303;
  assign N300 = N299 & N304;
  assign N301 = N300 & N305;
  assign N302 = N301 & N306;
  assign N1025 = N302 & io_resp_bits_entry[1];
  assign N303 = ~io_resp_bits_entry[4];
  assign N304 = ~io_resp_bits_entry[3];
  assign N305 = ~io_resp_bits_entry[2];
  assign N306 = ~io_resp_bits_entry[0];
  assign N307 = io_resp_bits_entry[5] & N311;
  assign N308 = N307 & N312;
  assign N309 = N308 & N313;
  assign N310 = N309 & io_resp_bits_entry[0];
  assign N1027 = N310 & io_resp_bits_entry[1];
  assign N311 = ~io_resp_bits_entry[4];
  assign N312 = ~io_resp_bits_entry[3];
  assign N313 = ~io_resp_bits_entry[2];
  assign N314 = io_resp_bits_entry[5] & N318;
  assign N315 = N314 & N319;
  assign N316 = N315 & io_resp_bits_entry[2];
  assign N317 = N316 & N320;
  assign N1029 = N317 & N321;
  assign N318 = ~io_resp_bits_entry[4];
  assign N319 = ~io_resp_bits_entry[3];
  assign N320 = ~io_resp_bits_entry[0];
  assign N321 = ~io_resp_bits_entry[1];
  assign N322 = io_resp_bits_entry[5] & N326;
  assign N323 = N322 & N327;
  assign N324 = N323 & io_resp_bits_entry[2];
  assign N325 = N324 & io_resp_bits_entry[0];
  assign N1031 = N325 & N328;
  assign N326 = ~io_resp_bits_entry[4];
  assign N327 = ~io_resp_bits_entry[3];
  assign N328 = ~io_resp_bits_entry[1];
  assign N329 = io_resp_bits_entry[5] & N333;
  assign N330 = N329 & N334;
  assign N331 = N330 & io_resp_bits_entry[2];
  assign N332 = N331 & N335;
  assign N1033 = N332 & io_resp_bits_entry[1];
  assign N333 = ~io_resp_bits_entry[4];
  assign N334 = ~io_resp_bits_entry[3];
  assign N335 = ~io_resp_bits_entry[0];
  assign N336 = io_resp_bits_entry[5] & N340;
  assign N337 = N336 & N341;
  assign N338 = N337 & io_resp_bits_entry[2];
  assign N339 = N338 & io_resp_bits_entry[0];
  assign N1035 = N339 & io_resp_bits_entry[1];
  assign N340 = ~io_resp_bits_entry[4];
  assign N341 = ~io_resp_bits_entry[3];
  assign N342 = io_resp_bits_entry[5] & N346;
  assign N343 = N342 & io_resp_bits_entry[3];
  assign N344 = N343 & N347;
  assign N345 = N344 & N348;
  assign N1037 = N345 & N349;
  assign N346 = ~io_resp_bits_entry[4];
  assign N347 = ~io_resp_bits_entry[2];
  assign N348 = ~io_resp_bits_entry[0];
  assign N349 = ~io_resp_bits_entry[1];
  assign N350 = io_resp_bits_entry[5] & N354;
  assign N351 = N350 & io_resp_bits_entry[3];
  assign N352 = N351 & N355;
  assign N353 = N352 & io_resp_bits_entry[0];
  assign N1039 = N353 & N356;
  assign N354 = ~io_resp_bits_entry[4];
  assign N355 = ~io_resp_bits_entry[2];
  assign N356 = ~io_resp_bits_entry[1];
  assign N357 = io_resp_bits_entry[5] & N361;
  assign N358 = N357 & io_resp_bits_entry[3];
  assign N359 = N358 & N362;
  assign N360 = N359 & N363;
  assign N1041 = N360 & io_resp_bits_entry[1];
  assign N361 = ~io_resp_bits_entry[4];
  assign N362 = ~io_resp_bits_entry[2];
  assign N363 = ~io_resp_bits_entry[0];
  assign N364 = io_resp_bits_entry[5] & N368;
  assign N365 = N364 & io_resp_bits_entry[3];
  assign N366 = N365 & N369;
  assign N367 = N366 & io_resp_bits_entry[0];
  assign N1043 = N367 & io_resp_bits_entry[1];
  assign N368 = ~io_resp_bits_entry[4];
  assign N369 = ~io_resp_bits_entry[2];
  assign N370 = io_resp_bits_entry[5] & N374;
  assign N371 = N370 & io_resp_bits_entry[3];
  assign N372 = N371 & io_resp_bits_entry[2];
  assign N373 = N372 & N375;
  assign N1045 = N373 & N376;
  assign N374 = ~io_resp_bits_entry[4];
  assign N375 = ~io_resp_bits_entry[0];
  assign N376 = ~io_resp_bits_entry[1];
  assign N377 = io_resp_bits_entry[5] & N381;
  assign N378 = N377 & io_resp_bits_entry[3];
  assign N379 = N378 & io_resp_bits_entry[2];
  assign N380 = N379 & io_resp_bits_entry[0];
  assign N1047 = N380 & N382;
  assign N381 = ~io_resp_bits_entry[4];
  assign N382 = ~io_resp_bits_entry[1];
  assign N1049 = io_resp_bits_entry[5] & io_resp_bits_entry[3] & (io_resp_bits_entry[2] & N383) & io_resp_bits_entry[1];
  assign N383 = ~io_resp_bits_entry[0];
  assign N1051 = io_resp_bits_entry[5] & io_resp_bits_entry[3] & (io_resp_bits_entry[2] & io_resp_bits_entry[0]) & io_resp_bits_entry[1];
  assign N384 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N385 = N384 & N388;
  assign N386 = N385 & N389;
  assign N387 = N386 & N390;
  assign N1053 = N387 & N391;
  assign N388 = ~io_resp_bits_entry[3];
  assign N389 = ~io_resp_bits_entry[2];
  assign N390 = ~io_resp_bits_entry[0];
  assign N391 = ~io_resp_bits_entry[1];
  assign N392 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N393 = N392 & N396;
  assign N394 = N393 & N397;
  assign N395 = N394 & io_resp_bits_entry[0];
  assign N1055 = N395 & N398;
  assign N396 = ~io_resp_bits_entry[3];
  assign N397 = ~io_resp_bits_entry[2];
  assign N398 = ~io_resp_bits_entry[1];
  assign N399 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N400 = N399 & N403;
  assign N401 = N400 & N404;
  assign N402 = N401 & N405;
  assign N1057 = N402 & io_resp_bits_entry[1];
  assign N403 = ~io_resp_bits_entry[3];
  assign N404 = ~io_resp_bits_entry[2];
  assign N405 = ~io_resp_bits_entry[0];
  assign N406 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N407 = N406 & N410;
  assign N408 = N407 & N411;
  assign N409 = N408 & io_resp_bits_entry[0];
  assign N1059 = N409 & io_resp_bits_entry[1];
  assign N410 = ~io_resp_bits_entry[3];
  assign N411 = ~io_resp_bits_entry[2];
  assign N412 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N413 = N412 & N416;
  assign N414 = N413 & io_resp_bits_entry[2];
  assign N415 = N414 & N417;
  assign N1061 = N415 & N418;
  assign N416 = ~io_resp_bits_entry[3];
  assign N417 = ~io_resp_bits_entry[0];
  assign N418 = ~io_resp_bits_entry[1];
  assign N419 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N420 = N419 & N423;
  assign N421 = N420 & io_resp_bits_entry[2];
  assign N422 = N421 & io_resp_bits_entry[0];
  assign N1063 = N422 & N424;
  assign N423 = ~io_resp_bits_entry[3];
  assign N424 = ~io_resp_bits_entry[1];
  assign N1065 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[2] & N425) & io_resp_bits_entry[1];
  assign N425 = ~io_resp_bits_entry[0];
  assign N1067 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[2] & io_resp_bits_entry[0]) & io_resp_bits_entry[1];
  assign N426 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N427 = N426 & io_resp_bits_entry[3];
  assign N428 = N427 & N430;
  assign N429 = N428 & N431;
  assign N1069 = N429 & N432;
  assign N430 = ~io_resp_bits_entry[2];
  assign N431 = ~io_resp_bits_entry[0];
  assign N432 = ~io_resp_bits_entry[1];
  assign N433 = io_resp_bits_entry[5] & io_resp_bits_entry[4];
  assign N434 = N433 & io_resp_bits_entry[3];
  assign N435 = N434 & N437;
  assign N436 = N435 & io_resp_bits_entry[0];
  assign N1071 = N436 & N438;
  assign N437 = ~io_resp_bits_entry[2];
  assign N438 = ~io_resp_bits_entry[1];
  assign N1073 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[3] & N439) & io_resp_bits_entry[1];
  assign N439 = ~io_resp_bits_entry[0];
  assign N1075 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[3] & io_resp_bits_entry[0]) & io_resp_bits_entry[1];
  assign N1077 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[3] & io_resp_bits_entry[2]) & N440;
  assign N440 = ~io_resp_bits_entry[0];
  assign N1079 = io_resp_bits_entry[5] & io_resp_bits_entry[4] & (io_resp_bits_entry[3] & io_resp_bits_entry[2]) & io_resp_bits_entry[0];
  assign T162 = (N441)? isJump_61 : 
                (N442)? 1'b0 : 1'b0;
  assign N441 = hits[61];
  assign N442 = N940;
  assign T169 = (N443)? R177 : 
                (N444)? nextRepl : 1'b0;
  assign N443 = updateHit;
  assign N444 = N941;
  assign T172 = (N445)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N446)? T173 : 1'b0;
  assign N445 = N2393;
  assign N446 = N2392;
  assign tgtPageReplEn = (N447)? tgtPageRepl : 
                         (N448)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N447 = doTgtPageRepl;
  assign N448 = N942;
  assign tgtPageRepl = (N449)? { T2420[0:0], T195 } : 
                       (N450)? T193 : 1'b0;
  assign N449 = samePage;
  assign N450 = N943;
  assign { T2420[0:0], T195 } = (N451)? updatePageHit : 
                                (N452)? idxPageRepl : 1'b0;
  assign N451 = N2829;
  assign N452 = N944;
  assign T200 = (N453)? { 1'b0, 1'b0, 1'b0 } : 
                (N454)? T201 : 1'b0;
  assign N453 = N2398;
  assign N454 = N2397;
  assign T214 = (N455)? io_req_bits_addr[38:12] : 
                (N456)? T209 : 1'b0;
  assign N455 = N2779;
  assign N456 = N945;
  assign T222 = (N455)? doTgtPageRepl : 
                (N456)? doIdxPageRepl : 1'b0;
  assign T232 = (N455)? T209 : 
                (N456)? io_req_bits_addr[38:12] : 1'b0;
  assign T238 = (N455)? doIdxPageRepl : 
                (N456)? doTgtPageRepl : 1'b0;
  assign idxPageReplEn = (N457)? idxPageRepl : 
                         (N458)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N457 = doIdxPageRepl;
  assign N458 = N946;
  assign T2435 = (N459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                 (N460)? T780 : 1'b0;
  assign N459 = reset;
  assign N460 = N1083;
  assign T780 = (N461)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                (N462)? T782 : 1'b0;
  assign N461 = io_invalidate;
  assign N462 = N947;
  assign { T799, T2444, T2445[1:1] } = (N463)? pageHit[5:1] : 
                                       (N464)? tgtPageRepl[5:1] : 1'b0;
  assign N463 = N2789;
  assign N464 = N949;
  assign T1163 = (N465)? isJump_60 : 
                 (N466)? 1'b0 : 1'b0;
  assign N465 = hits[60];
  assign N466 = N950;
  assign T1169 = (N467)? isJump_59 : 
                 (N468)? 1'b0 : 1'b0;
  assign N467 = hits[59];
  assign N468 = N951;
  assign T1175 = (N469)? isJump_58 : 
                 (N470)? 1'b0 : 1'b0;
  assign N469 = hits[58];
  assign N470 = N952;
  assign T1181 = (N471)? isJump_57 : 
                 (N472)? 1'b0 : 1'b0;
  assign N471 = hits[57];
  assign N472 = N953;
  assign T1187 = (N473)? isJump_56 : 
                 (N474)? 1'b0 : 1'b0;
  assign N473 = hits[56];
  assign N474 = N954;
  assign T1193 = (N475)? isJump_55 : 
                 (N476)? 1'b0 : 1'b0;
  assign N475 = hits[55];
  assign N476 = N955;
  assign T1199 = (N477)? isJump_54 : 
                 (N478)? 1'b0 : 1'b0;
  assign N477 = hits[54];
  assign N478 = N956;
  assign T1205 = (N479)? isJump_53 : 
                 (N480)? 1'b0 : 1'b0;
  assign N479 = hits[53];
  assign N480 = N957;
  assign T1211 = (N481)? isJump_52 : 
                 (N482)? 1'b0 : 1'b0;
  assign N481 = hits[52];
  assign N482 = N958;
  assign T1217 = (N483)? isJump_51 : 
                 (N484)? 1'b0 : 1'b0;
  assign N483 = hits[51];
  assign N484 = N959;
  assign T1223 = (N485)? isJump_50 : 
                 (N486)? 1'b0 : 1'b0;
  assign N485 = hits[50];
  assign N486 = N960;
  assign T1229 = (N487)? isJump_49 : 
                 (N488)? 1'b0 : 1'b0;
  assign N487 = hits[49];
  assign N488 = N961;
  assign T1235 = (N489)? isJump_48 : 
                 (N490)? 1'b0 : 1'b0;
  assign N489 = hits[48];
  assign N490 = N962;
  assign T1241 = (N491)? isJump_47 : 
                 (N492)? 1'b0 : 1'b0;
  assign N491 = hits[47];
  assign N492 = N963;
  assign T1247 = (N493)? isJump_46 : 
                 (N494)? 1'b0 : 1'b0;
  assign N493 = hits[46];
  assign N494 = N964;
  assign T1253 = (N495)? isJump_45 : 
                 (N496)? 1'b0 : 1'b0;
  assign N495 = hits[45];
  assign N496 = N965;
  assign T1259 = (N497)? isJump_44 : 
                 (N498)? 1'b0 : 1'b0;
  assign N497 = hits[44];
  assign N498 = N966;
  assign T1265 = (N499)? isJump_43 : 
                 (N500)? 1'b0 : 1'b0;
  assign N499 = hits[43];
  assign N500 = N967;
  assign T1271 = (N501)? isJump_42 : 
                 (N502)? 1'b0 : 1'b0;
  assign N501 = hits[42];
  assign N502 = N968;
  assign T1277 = (N503)? isJump_41 : 
                 (N504)? 1'b0 : 1'b0;
  assign N503 = hits[41];
  assign N504 = N969;
  assign T1283 = (N505)? isJump_40 : 
                 (N506)? 1'b0 : 1'b0;
  assign N505 = hits[40];
  assign N506 = N970;
  assign T1289 = (N507)? isJump_39 : 
                 (N508)? 1'b0 : 1'b0;
  assign N507 = hits[39];
  assign N508 = N971;
  assign T1295 = (N509)? isJump_38 : 
                 (N510)? 1'b0 : 1'b0;
  assign N509 = hits[38];
  assign N510 = N972;
  assign T1301 = (N511)? isJump_37 : 
                 (N512)? 1'b0 : 1'b0;
  assign N511 = hits[37];
  assign N512 = N973;
  assign T1307 = (N513)? isJump_36 : 
                 (N514)? 1'b0 : 1'b0;
  assign N513 = hits[36];
  assign N514 = N974;
  assign T1313 = (N515)? isJump_35 : 
                 (N516)? 1'b0 : 1'b0;
  assign N515 = hits[35];
  assign N516 = N975;
  assign T1319 = (N517)? isJump_34 : 
                 (N518)? 1'b0 : 1'b0;
  assign N517 = hits[34];
  assign N518 = N976;
  assign T1325 = (N519)? isJump_33 : 
                 (N520)? 1'b0 : 1'b0;
  assign N519 = hits[33];
  assign N520 = N977;
  assign T1331 = (N521)? isJump_32 : 
                 (N522)? 1'b0 : 1'b0;
  assign N521 = hits[32];
  assign N522 = N978;
  assign T1337 = (N523)? isJump_31 : 
                 (N524)? 1'b0 : 1'b0;
  assign N523 = hits[31];
  assign N524 = N979;
  assign T1343 = (N525)? isJump_30 : 
                 (N526)? 1'b0 : 1'b0;
  assign N525 = hits[30];
  assign N526 = N980;
  assign T1349 = (N527)? isJump_29 : 
                 (N528)? 1'b0 : 1'b0;
  assign N527 = hits[29];
  assign N528 = N981;
  assign T1355 = (N529)? isJump_28 : 
                 (N530)? 1'b0 : 1'b0;
  assign N529 = hits[28];
  assign N530 = N982;
  assign T1361 = (N531)? isJump_27 : 
                 (N532)? 1'b0 : 1'b0;
  assign N531 = hits[27];
  assign N532 = N983;
  assign T1367 = (N533)? isJump_26 : 
                 (N534)? 1'b0 : 1'b0;
  assign N533 = hits[26];
  assign N534 = N984;
  assign T1373 = (N535)? isJump_25 : 
                 (N536)? 1'b0 : 1'b0;
  assign N535 = hits[25];
  assign N536 = N985;
  assign T1379 = (N537)? isJump_24 : 
                 (N538)? 1'b0 : 1'b0;
  assign N537 = hits[24];
  assign N538 = N986;
  assign T1385 = (N539)? isJump_23 : 
                 (N540)? 1'b0 : 1'b0;
  assign N539 = hits[23];
  assign N540 = N987;
  assign T1391 = (N541)? isJump_22 : 
                 (N542)? 1'b0 : 1'b0;
  assign N541 = hits[22];
  assign N542 = N988;
  assign T1397 = (N543)? isJump_21 : 
                 (N544)? 1'b0 : 1'b0;
  assign N543 = hits[21];
  assign N544 = N989;
  assign T1403 = (N545)? isJump_20 : 
                 (N546)? 1'b0 : 1'b0;
  assign N545 = hits[20];
  assign N546 = N990;
  assign T1409 = (N547)? isJump_19 : 
                 (N548)? 1'b0 : 1'b0;
  assign N547 = hits[19];
  assign N548 = N991;
  assign T1415 = (N549)? isJump_18 : 
                 (N550)? 1'b0 : 1'b0;
  assign N549 = hits[18];
  assign N550 = N992;
  assign T1421 = (N551)? isJump_17 : 
                 (N552)? 1'b0 : 1'b0;
  assign N551 = hits[17];
  assign N552 = N993;
  assign T1427 = (N553)? isJump_16 : 
                 (N554)? 1'b0 : 1'b0;
  assign N553 = hits[16];
  assign N554 = N994;
  assign T1433 = (N555)? isJump_15 : 
                 (N556)? 1'b0 : 1'b0;
  assign N555 = hits[15];
  assign N556 = N995;
  assign T1439 = (N557)? isJump_14 : 
                 (N558)? 1'b0 : 1'b0;
  assign N557 = hits[14];
  assign N558 = N996;
  assign T1445 = (N559)? isJump_13 : 
                 (N560)? 1'b0 : 1'b0;
  assign N559 = hits[13];
  assign N560 = N997;
  assign T1451 = (N561)? isJump_12 : 
                 (N562)? 1'b0 : 1'b0;
  assign N561 = hits[12];
  assign N562 = N998;
  assign T1457 = (N563)? isJump_11 : 
                 (N564)? 1'b0 : 1'b0;
  assign N563 = hits[11];
  assign N564 = N999;
  assign T1463 = (N565)? isJump_10 : 
                 (N566)? 1'b0 : 1'b0;
  assign N565 = hits[10];
  assign N566 = N1000;
  assign T1469 = (N567)? isJump_9 : 
                 (N568)? 1'b0 : 1'b0;
  assign N567 = hits[9];
  assign N568 = N1001;
  assign T1475 = (N569)? isJump_8 : 
                 (N570)? 1'b0 : 1'b0;
  assign N569 = hits[8];
  assign N570 = N1002;
  assign T1481 = (N571)? isJump_7 : 
                 (N572)? 1'b0 : 1'b0;
  assign N571 = hits[7];
  assign N572 = N1003;
  assign T1487 = (N573)? isJump_6 : 
                 (N574)? 1'b0 : 1'b0;
  assign N573 = hits[6];
  assign N574 = N1004;
  assign T1493 = (N575)? isJump_5 : 
                 (N576)? 1'b0 : 1'b0;
  assign N575 = hits[5];
  assign N576 = N1005;
  assign T1499 = (N577)? isJump_4 : 
                 (N578)? 1'b0 : 1'b0;
  assign N577 = hits[4];
  assign N578 = N1006;
  assign T1505 = (N579)? isJump_3 : 
                 (N580)? 1'b0 : 1'b0;
  assign N579 = hits[3];
  assign N580 = N1007;
  assign T1511 = (N581)? isJump_2 : 
                 (N582)? 1'b0 : 1'b0;
  assign N581 = hits[2];
  assign N582 = N1008;
  assign T1517 = (N583)? isJump_1 : 
                 (N584)? 1'b0 : 1'b0;
  assign N583 = hits[1];
  assign N584 = N1009;
  assign T1522 = (N585)? isJump_0 : 
                 (N586)? 1'b0 : 1'b0;
  assign N585 = hits[0];
  assign N586 = N1010;
  assign io_resp_bits_target = (N587)? io_ras_update_bits_returnAddr : 
                               (N588)? T1535 : 1'b0;
  assign N587 = T2406;
  assign N588 = N1011;
  assign T1535 = (N589)? T1995 : 
                 (N590)? T1536 : 1'b0;
  assign N589 = T2028;
  assign N590 = N1012;
  assign T1538 = (N441)? T1539 : 
                 (N442)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1545 = (N465)? T1546 : 
                 (N466)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1549 = (N467)? T1550 : 
                 (N468)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1553 = (N469)? T1554 : 
                 (N470)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1557 = (N471)? T1558 : 
                 (N472)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1561 = (N473)? T1562 : 
                 (N474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1565 = (N475)? T1566 : 
                 (N476)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1569 = (N477)? T1570 : 
                 (N478)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1573 = (N479)? T1574 : 
                 (N480)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1577 = (N481)? T1578 : 
                 (N482)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1581 = (N483)? T1582 : 
                 (N484)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1585 = (N485)? T1586 : 
                 (N486)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1589 = (N487)? T1590 : 
                 (N488)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1593 = (N489)? T1594 : 
                 (N490)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1597 = (N491)? T1598 : 
                 (N492)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1601 = (N493)? T1602 : 
                 (N494)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1605 = (N495)? T1606 : 
                 (N496)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1609 = (N497)? T1610 : 
                 (N498)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1613 = (N499)? T1614 : 
                 (N500)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1617 = (N501)? T1618 : 
                 (N502)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1621 = (N503)? T1622 : 
                 (N504)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1625 = (N505)? T1626 : 
                 (N506)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1629 = (N507)? T1630 : 
                 (N508)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1633 = (N509)? T1634 : 
                 (N510)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1637 = (N511)? T1638 : 
                 (N512)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1641 = (N513)? T1642 : 
                 (N514)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1645 = (N515)? T1646 : 
                 (N516)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1649 = (N517)? T1650 : 
                 (N518)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1653 = (N519)? T1654 : 
                 (N520)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1657 = (N521)? T1658 : 
                 (N522)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1661 = (N523)? T1662 : 
                 (N524)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1665 = (N525)? T1666 : 
                 (N526)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1669 = (N527)? T1670 : 
                 (N528)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1673 = (N529)? T1674 : 
                 (N530)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1677 = (N531)? T1678 : 
                 (N532)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1681 = (N533)? T1682 : 
                 (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1685 = (N535)? T1686 : 
                 (N536)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1689 = (N537)? T1690 : 
                 (N538)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1693 = (N539)? T1694 : 
                 (N540)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1697 = (N541)? T1698 : 
                 (N542)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1701 = (N543)? T1702 : 
                 (N544)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1705 = (N545)? T1706 : 
                 (N546)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1709 = (N547)? T1710 : 
                 (N548)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1713 = (N549)? T1714 : 
                 (N550)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1717 = (N551)? T1718 : 
                 (N552)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1721 = (N553)? T1722 : 
                 (N554)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1725 = (N555)? T1726 : 
                 (N556)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1729 = (N557)? T1730 : 
                 (N558)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1733 = (N559)? T1734 : 
                 (N560)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1737 = (N561)? T1738 : 
                 (N562)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1741 = (N563)? T1742 : 
                 (N564)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1745 = (N565)? T1746 : 
                 (N566)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1749 = (N567)? T1750 : 
                 (N568)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1753 = (N569)? T1754 : 
                 (N570)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1757 = (N571)? T1758 : 
                 (N572)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1761 = (N573)? T1762 : 
                 (N574)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1765 = (N575)? T1766 : 
                 (N576)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1769 = (N577)? T1770 : 
                 (N578)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1773 = (N579)? T1774 : 
                 (N580)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1777 = (N581)? T1778 : 
                 (N582)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1781 = (N583)? T1782 : 
                 (N584)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1784 = (N585)? T1785 : 
                 (N586)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1788 = (N591)? T258 : 
                 (N592)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N591 = T1791[5];
  assign N592 = N1013;
  assign T1792 = (N441)? tgtPagesOH_61 : 
                 (N442)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1795 = (N465)? tgtPagesOH_60 : 
                 (N466)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1798 = (N467)? tgtPagesOH_59 : 
                 (N468)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1801 = (N469)? tgtPagesOH_58 : 
                 (N470)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1804 = (N471)? tgtPagesOH_57 : 
                 (N472)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1807 = (N473)? tgtPagesOH_56 : 
                 (N474)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1810 = (N475)? tgtPagesOH_55 : 
                 (N476)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1813 = (N477)? tgtPagesOH_54 : 
                 (N478)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1816 = (N479)? tgtPagesOH_53 : 
                 (N480)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1819 = (N481)? tgtPagesOH_52 : 
                 (N482)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1822 = (N483)? tgtPagesOH_51 : 
                 (N484)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1825 = (N485)? tgtPagesOH_50 : 
                 (N486)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1828 = (N487)? tgtPagesOH_49 : 
                 (N488)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1831 = (N489)? tgtPagesOH_48 : 
                 (N490)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1834 = (N491)? tgtPagesOH_47 : 
                 (N492)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1837 = (N493)? tgtPagesOH_46 : 
                 (N494)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1840 = (N495)? tgtPagesOH_45 : 
                 (N496)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1843 = (N497)? tgtPagesOH_44 : 
                 (N498)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1846 = (N499)? tgtPagesOH_43 : 
                 (N500)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1849 = (N501)? tgtPagesOH_42 : 
                 (N502)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1852 = (N503)? tgtPagesOH_41 : 
                 (N504)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1855 = (N505)? tgtPagesOH_40 : 
                 (N506)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1858 = (N507)? tgtPagesOH_39 : 
                 (N508)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1861 = (N509)? tgtPagesOH_38 : 
                 (N510)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1864 = (N511)? tgtPagesOH_37 : 
                 (N512)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1867 = (N513)? tgtPagesOH_36 : 
                 (N514)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1870 = (N515)? tgtPagesOH_35 : 
                 (N516)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1873 = (N517)? tgtPagesOH_34 : 
                 (N518)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1876 = (N519)? tgtPagesOH_33 : 
                 (N520)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1879 = (N521)? tgtPagesOH_32 : 
                 (N522)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1882 = (N523)? tgtPagesOH_31 : 
                 (N524)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1885 = (N525)? tgtPagesOH_30 : 
                 (N526)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1888 = (N527)? tgtPagesOH_29 : 
                 (N528)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1891 = (N529)? tgtPagesOH_28 : 
                 (N530)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1894 = (N531)? tgtPagesOH_27 : 
                 (N532)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1897 = (N533)? tgtPagesOH_26 : 
                 (N534)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1900 = (N535)? tgtPagesOH_25 : 
                 (N536)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1903 = (N537)? tgtPagesOH_24 : 
                 (N538)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1906 = (N539)? tgtPagesOH_23 : 
                 (N540)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1909 = (N541)? tgtPagesOH_22 : 
                 (N542)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1912 = (N543)? tgtPagesOH_21 : 
                 (N544)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1915 = (N545)? tgtPagesOH_20 : 
                 (N546)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1918 = (N547)? tgtPagesOH_19 : 
                 (N548)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1921 = (N549)? tgtPagesOH_18 : 
                 (N550)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1924 = (N551)? tgtPagesOH_17 : 
                 (N552)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1927 = (N553)? tgtPagesOH_16 : 
                 (N554)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1930 = (N555)? tgtPagesOH_15 : 
                 (N556)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1933 = (N557)? tgtPagesOH_14 : 
                 (N558)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1936 = (N559)? tgtPagesOH_13 : 
                 (N560)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1939 = (N561)? tgtPagesOH_12 : 
                 (N562)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1942 = (N563)? tgtPagesOH_11 : 
                 (N564)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1945 = (N565)? tgtPagesOH_10 : 
                 (N566)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1948 = (N567)? tgtPagesOH_9 : 
                 (N568)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1951 = (N569)? tgtPagesOH_8 : 
                 (N570)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1954 = (N571)? tgtPagesOH_7 : 
                 (N572)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1957 = (N573)? tgtPagesOH_6 : 
                 (N574)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1960 = (N575)? tgtPagesOH_5 : 
                 (N576)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1963 = (N577)? tgtPagesOH_4 : 
                 (N578)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1966 = (N579)? tgtPagesOH_3 : 
                 (N580)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1969 = (N581)? tgtPagesOH_2 : 
                 (N582)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1972 = (N583)? tgtPagesOH_1 : 
                 (N584)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1974 = (N585)? tgtPagesOH_0 : 
                 (N586)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign T1977 = (N593)? T256 : 
                 (N594)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N593 = T1791[4];
  assign N594 = N1014;
  assign T1981 = (N595)? T254 : 
                 (N596)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N595 = T1791[3];
  assign N596 = N1015;
  assign T1985 = (N597)? T250 : 
                 (N598)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N597 = T1791[2];
  assign N598 = N1016;
  assign T1989 = (N599)? T248 : 
                 (N600)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N599 = T1791[1];
  assign N600 = N1017;
  assign T1992 = (N601)? T212 : 
                 (N602)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N601 = T1791[0];
  assign N602 = N1018;
  assign T1995 = (N603)? R2023 : 
                 (N604)? R1996 : 1'b0;
  assign N603 = T2027;
  assign N604 = N1019;
  assign T2030 = (N441)? useRAS_61 : 
                 (N442)? 1'b0 : 1'b0;
  assign T2040 = (N465)? useRAS_60 : 
                 (N466)? 1'b0 : 1'b0;
  assign T2046 = (N467)? useRAS_59 : 
                 (N468)? 1'b0 : 1'b0;
  assign T2052 = (N469)? useRAS_58 : 
                 (N470)? 1'b0 : 1'b0;
  assign T2058 = (N471)? useRAS_57 : 
                 (N472)? 1'b0 : 1'b0;
  assign T2064 = (N473)? useRAS_56 : 
                 (N474)? 1'b0 : 1'b0;
  assign T2070 = (N475)? useRAS_55 : 
                 (N476)? 1'b0 : 1'b0;
  assign T2076 = (N477)? useRAS_54 : 
                 (N478)? 1'b0 : 1'b0;
  assign T2082 = (N479)? useRAS_53 : 
                 (N480)? 1'b0 : 1'b0;
  assign T2088 = (N481)? useRAS_52 : 
                 (N482)? 1'b0 : 1'b0;
  assign T2094 = (N483)? useRAS_51 : 
                 (N484)? 1'b0 : 1'b0;
  assign T2100 = (N485)? useRAS_50 : 
                 (N486)? 1'b0 : 1'b0;
  assign T2106 = (N487)? useRAS_49 : 
                 (N488)? 1'b0 : 1'b0;
  assign T2112 = (N489)? useRAS_48 : 
                 (N490)? 1'b0 : 1'b0;
  assign T2118 = (N491)? useRAS_47 : 
                 (N492)? 1'b0 : 1'b0;
  assign T2124 = (N493)? useRAS_46 : 
                 (N494)? 1'b0 : 1'b0;
  assign T2130 = (N495)? useRAS_45 : 
                 (N496)? 1'b0 : 1'b0;
  assign T2136 = (N497)? useRAS_44 : 
                 (N498)? 1'b0 : 1'b0;
  assign T2142 = (N499)? useRAS_43 : 
                 (N500)? 1'b0 : 1'b0;
  assign T2148 = (N501)? useRAS_42 : 
                 (N502)? 1'b0 : 1'b0;
  assign T2154 = (N503)? useRAS_41 : 
                 (N504)? 1'b0 : 1'b0;
  assign T2160 = (N505)? useRAS_40 : 
                 (N506)? 1'b0 : 1'b0;
  assign T2166 = (N507)? useRAS_39 : 
                 (N508)? 1'b0 : 1'b0;
  assign T2172 = (N509)? useRAS_38 : 
                 (N510)? 1'b0 : 1'b0;
  assign T2178 = (N511)? useRAS_37 : 
                 (N512)? 1'b0 : 1'b0;
  assign T2184 = (N513)? useRAS_36 : 
                 (N514)? 1'b0 : 1'b0;
  assign T2190 = (N515)? useRAS_35 : 
                 (N516)? 1'b0 : 1'b0;
  assign T2196 = (N517)? useRAS_34 : 
                 (N518)? 1'b0 : 1'b0;
  assign T2202 = (N519)? useRAS_33 : 
                 (N520)? 1'b0 : 1'b0;
  assign T2208 = (N521)? useRAS_32 : 
                 (N522)? 1'b0 : 1'b0;
  assign T2214 = (N523)? useRAS_31 : 
                 (N524)? 1'b0 : 1'b0;
  assign T2220 = (N525)? useRAS_30 : 
                 (N526)? 1'b0 : 1'b0;
  assign T2226 = (N527)? useRAS_29 : 
                 (N528)? 1'b0 : 1'b0;
  assign T2232 = (N529)? useRAS_28 : 
                 (N530)? 1'b0 : 1'b0;
  assign T2238 = (N531)? useRAS_27 : 
                 (N532)? 1'b0 : 1'b0;
  assign T2244 = (N533)? useRAS_26 : 
                 (N534)? 1'b0 : 1'b0;
  assign T2250 = (N535)? useRAS_25 : 
                 (N536)? 1'b0 : 1'b0;
  assign T2256 = (N537)? useRAS_24 : 
                 (N538)? 1'b0 : 1'b0;
  assign T2262 = (N539)? useRAS_23 : 
                 (N540)? 1'b0 : 1'b0;
  assign T2268 = (N541)? useRAS_22 : 
                 (N542)? 1'b0 : 1'b0;
  assign T2274 = (N543)? useRAS_21 : 
                 (N544)? 1'b0 : 1'b0;
  assign T2280 = (N545)? useRAS_20 : 
                 (N546)? 1'b0 : 1'b0;
  assign T2286 = (N547)? useRAS_19 : 
                 (N548)? 1'b0 : 1'b0;
  assign T2292 = (N549)? useRAS_18 : 
                 (N550)? 1'b0 : 1'b0;
  assign T2298 = (N551)? useRAS_17 : 
                 (N552)? 1'b0 : 1'b0;
  assign T2304 = (N553)? useRAS_16 : 
                 (N554)? 1'b0 : 1'b0;
  assign T2310 = (N555)? useRAS_15 : 
                 (N556)? 1'b0 : 1'b0;
  assign T2316 = (N557)? useRAS_14 : 
                 (N558)? 1'b0 : 1'b0;
  assign T2322 = (N559)? useRAS_13 : 
                 (N560)? 1'b0 : 1'b0;
  assign T2328 = (N561)? useRAS_12 : 
                 (N562)? 1'b0 : 1'b0;
  assign T2334 = (N563)? useRAS_11 : 
                 (N564)? 1'b0 : 1'b0;
  assign T2340 = (N565)? useRAS_10 : 
                 (N566)? 1'b0 : 1'b0;
  assign T2346 = (N567)? useRAS_9 : 
                 (N568)? 1'b0 : 1'b0;
  assign T2352 = (N569)? useRAS_8 : 
                 (N570)? 1'b0 : 1'b0;
  assign T2358 = (N571)? useRAS_7 : 
                 (N572)? 1'b0 : 1'b0;
  assign T2364 = (N573)? useRAS_6 : 
                 (N574)? 1'b0 : 1'b0;
  assign T2370 = (N575)? useRAS_5 : 
                 (N576)? 1'b0 : 1'b0;
  assign T2376 = (N577)? useRAS_4 : 
                 (N578)? 1'b0 : 1'b0;
  assign T2382 = (N579)? useRAS_3 : 
                 (N580)? 1'b0 : 1'b0;
  assign T2388 = (N581)? useRAS_2 : 
                 (N582)? 1'b0 : 1'b0;
  assign T2394 = (N583)? useRAS_1 : 
                 (N584)? 1'b0 : 1'b0;
  assign T2399 = (N585)? useRAS_0 : 
                 (N586)? 1'b0 : 1'b0;
  assign io_resp_bits_taken = (N605)? 1'b0 : 
                              (N606)? io_resp_valid : 1'b0;
  assign N605 = T2412;
  assign N606 = N1082;
  assign N1084 = (N459)? 1'b0 : 
                 (N460)? io_btb_update_valid : 1'b0;
  assign { N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214 } = (N607)? { N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N608)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N607 = T21;
  assign N608 = N1085;
  assign N1342 = (N459)? 1'b1 : 
                 (N460)? N1341 : 1'b0;
  assign { N1344, N1343 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1345 = (N459)? 1'b1 : 
                 (N460)? N1340 : 1'b0;
  assign { N1347, N1346 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1348 = (N459)? 1'b1 : 
                 (N460)? N1339 : 1'b0;
  assign { N1350, N1349 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1351 = (N459)? 1'b1 : 
                 (N460)? N1338 : 1'b0;
  assign { N1353, N1352 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1354 = (N459)? 1'b1 : 
                 (N460)? N1337 : 1'b0;
  assign { N1356, N1355 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1357 = (N459)? 1'b1 : 
                 (N460)? N1336 : 1'b0;
  assign { N1359, N1358 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1360 = (N459)? 1'b1 : 
                 (N460)? N1335 : 1'b0;
  assign { N1362, N1361 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1363 = (N459)? 1'b1 : 
                 (N460)? N1334 : 1'b0;
  assign { N1365, N1364 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1366 = (N459)? 1'b1 : 
                 (N460)? N1333 : 1'b0;
  assign { N1368, N1367 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1369 = (N459)? 1'b1 : 
                 (N460)? N1332 : 1'b0;
  assign { N1371, N1370 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1372 = (N459)? 1'b1 : 
                 (N460)? N1331 : 1'b0;
  assign { N1374, N1373 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1375 = (N459)? 1'b1 : 
                 (N460)? N1330 : 1'b0;
  assign { N1377, N1376 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1378 = (N459)? 1'b1 : 
                 (N460)? N1329 : 1'b0;
  assign { N1380, N1379 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1381 = (N459)? 1'b1 : 
                 (N460)? N1328 : 1'b0;
  assign { N1383, N1382 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1384 = (N459)? 1'b1 : 
                 (N460)? N1327 : 1'b0;
  assign { N1386, N1385 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1387 = (N459)? 1'b1 : 
                 (N460)? N1326 : 1'b0;
  assign { N1389, N1388 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1390 = (N459)? 1'b1 : 
                 (N460)? N1325 : 1'b0;
  assign { N1392, N1391 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1393 = (N459)? 1'b1 : 
                 (N460)? N1324 : 1'b0;
  assign { N1395, N1394 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1396 = (N459)? 1'b1 : 
                 (N460)? N1323 : 1'b0;
  assign { N1398, N1397 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1399 = (N459)? 1'b1 : 
                 (N460)? N1322 : 1'b0;
  assign { N1401, N1400 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1402 = (N459)? 1'b1 : 
                 (N460)? N1321 : 1'b0;
  assign { N1404, N1403 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1405 = (N459)? 1'b1 : 
                 (N460)? N1320 : 1'b0;
  assign { N1407, N1406 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1408 = (N459)? 1'b1 : 
                 (N460)? N1319 : 1'b0;
  assign { N1410, N1409 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1411 = (N459)? 1'b1 : 
                 (N460)? N1318 : 1'b0;
  assign { N1413, N1412 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1414 = (N459)? 1'b1 : 
                 (N460)? N1317 : 1'b0;
  assign { N1416, N1415 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1417 = (N459)? 1'b1 : 
                 (N460)? N1316 : 1'b0;
  assign { N1419, N1418 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1420 = (N459)? 1'b1 : 
                 (N460)? N1315 : 1'b0;
  assign { N1422, N1421 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1423 = (N459)? 1'b1 : 
                 (N460)? N1314 : 1'b0;
  assign { N1425, N1424 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1426 = (N459)? 1'b1 : 
                 (N460)? N1313 : 1'b0;
  assign { N1428, N1427 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1429 = (N459)? 1'b1 : 
                 (N460)? N1312 : 1'b0;
  assign { N1431, N1430 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1432 = (N459)? 1'b1 : 
                 (N460)? N1311 : 1'b0;
  assign N1433 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1434 = (N459)? 1'b1 : 
                 (N460)? N1310 : 1'b0;
  assign N1435 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1436 = (N459)? 1'b1 : 
                 (N460)? N1309 : 1'b0;
  assign N1437 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1438 = (N459)? 1'b1 : 
                 (N460)? N1308 : 1'b0;
  assign N1439 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1440 = (N459)? 1'b1 : 
                 (N460)? N1307 : 1'b0;
  assign N1441 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1442 = (N459)? 1'b1 : 
                 (N460)? N1306 : 1'b0;
  assign N1443 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1444 = (N459)? 1'b1 : 
                 (N460)? N1305 : 1'b0;
  assign N1445 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1446 = (N459)? 1'b1 : 
                 (N460)? N1304 : 1'b0;
  assign N1447 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1448 = (N459)? 1'b1 : 
                 (N460)? N1303 : 1'b0;
  assign N1449 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1450 = (N459)? 1'b1 : 
                 (N460)? N1302 : 1'b0;
  assign N1451 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1452 = (N459)? 1'b1 : 
                 (N460)? N1301 : 1'b0;
  assign N1453 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1454 = (N459)? 1'b1 : 
                 (N460)? N1300 : 1'b0;
  assign N1455 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1456 = (N459)? 1'b1 : 
                 (N460)? N1299 : 1'b0;
  assign N1457 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1458 = (N459)? 1'b1 : 
                 (N460)? N1298 : 1'b0;
  assign N1459 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1460 = (N459)? 1'b1 : 
                 (N460)? N1297 : 1'b0;
  assign N1461 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1462 = (N459)? 1'b1 : 
                 (N460)? N1296 : 1'b0;
  assign N1463 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1464 = (N459)? 1'b1 : 
                 (N460)? N1295 : 1'b0;
  assign N1465 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1466 = (N459)? 1'b1 : 
                 (N460)? N1294 : 1'b0;
  assign { N1468, N1467 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1469 = (N459)? 1'b1 : 
                 (N460)? N1293 : 1'b0;
  assign N1470 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1471 = (N459)? 1'b1 : 
                 (N460)? N1292 : 1'b0;
  assign N1472 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1473 = (N459)? 1'b1 : 
                 (N460)? N1291 : 1'b0;
  assign N1474 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1475 = (N459)? 1'b1 : 
                 (N460)? N1290 : 1'b0;
  assign N1476 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1477 = (N459)? 1'b1 : 
                 (N460)? N1289 : 1'b0;
  assign N1478 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1479 = (N459)? 1'b1 : 
                 (N460)? N1288 : 1'b0;
  assign { N1481, N1480 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1482 = (N459)? 1'b1 : 
                 (N460)? N1287 : 1'b0;
  assign N1483 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1484 = (N459)? 1'b1 : 
                 (N460)? N1286 : 1'b0;
  assign N1485 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1486 = (N459)? 1'b1 : 
                 (N460)? N1285 : 1'b0;
  assign N1487 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1488 = (N459)? 1'b1 : 
                 (N460)? N1284 : 1'b0;
  assign N1489 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1490 = (N459)? 1'b1 : 
                 (N460)? N1283 : 1'b0;
  assign N1491 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1492 = (N459)? 1'b1 : 
                 (N460)? N1282 : 1'b0;
  assign N1493 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1494 = (N459)? 1'b1 : 
                 (N460)? N1281 : 1'b0;
  assign N1495 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1496 = (N459)? 1'b1 : 
                 (N460)? N1280 : 1'b0;
  assign N1497 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1498 = (N459)? 1'b1 : 
                 (N460)? N1279 : 1'b0;
  assign N1499 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1500 = (N459)? 1'b1 : 
                 (N460)? N1278 : 1'b0;
  assign N1501 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1502 = (N459)? 1'b1 : 
                 (N460)? N1277 : 1'b0;
  assign N1503 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1504 = (N459)? 1'b1 : 
                 (N460)? N1276 : 1'b0;
  assign N1505 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1506 = (N459)? 1'b1 : 
                 (N460)? N1275 : 1'b0;
  assign N1507 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1508 = (N459)? 1'b1 : 
                 (N460)? N1274 : 1'b0;
  assign N1509 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1510 = (N459)? 1'b1 : 
                 (N460)? N1273 : 1'b0;
  assign N1511 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1512 = (N459)? 1'b1 : 
                 (N460)? N1272 : 1'b0;
  assign N1513 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1514 = (N459)? 1'b1 : 
                 (N460)? N1271 : 1'b0;
  assign N1515 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1516 = (N459)? 1'b1 : 
                 (N460)? N1270 : 1'b0;
  assign { N1518, N1517 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1519 = (N459)? 1'b1 : 
                 (N460)? N1269 : 1'b0;
  assign N1520 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1521 = (N459)? 1'b1 : 
                 (N460)? N1268 : 1'b0;
  assign N1522 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1523 = (N459)? 1'b1 : 
                 (N460)? N1267 : 1'b0;
  assign N1524 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1525 = (N459)? 1'b1 : 
                 (N460)? N1266 : 1'b0;
  assign N1526 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1527 = (N459)? 1'b1 : 
                 (N460)? N1265 : 1'b0;
  assign N1528 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1529 = (N459)? 1'b1 : 
                 (N460)? N1264 : 1'b0;
  assign N1530 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1531 = (N459)? 1'b1 : 
                 (N460)? N1263 : 1'b0;
  assign { N1533, N1532 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1534 = (N459)? 1'b1 : 
                 (N460)? N1262 : 1'b0;
  assign N1535 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1536 = (N459)? 1'b1 : 
                 (N460)? N1261 : 1'b0;
  assign N1537 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1538 = (N459)? 1'b1 : 
                 (N460)? N1260 : 1'b0;
  assign N1539 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1540 = (N459)? 1'b1 : 
                 (N460)? N1259 : 1'b0;
  assign N1541 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1542 = (N459)? 1'b1 : 
                 (N460)? N1258 : 1'b0;
  assign N1543 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1544 = (N459)? 1'b1 : 
                 (N460)? N1257 : 1'b0;
  assign N1545 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1546 = (N459)? 1'b1 : 
                 (N460)? N1256 : 1'b0;
  assign N1547 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1548 = (N459)? 1'b1 : 
                 (N460)? N1255 : 1'b0;
  assign N1549 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1550 = (N459)? 1'b1 : 
                 (N460)? N1254 : 1'b0;
  assign N1551 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1552 = (N459)? 1'b1 : 
                 (N460)? N1253 : 1'b0;
  assign N1553 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1554 = (N459)? 1'b1 : 
                 (N460)? N1252 : 1'b0;
  assign N1555 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1556 = (N459)? 1'b1 : 
                 (N460)? N1251 : 1'b0;
  assign N1557 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1558 = (N459)? 1'b1 : 
                 (N460)? N1250 : 1'b0;
  assign N1559 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1560 = (N459)? 1'b1 : 
                 (N460)? N1249 : 1'b0;
  assign N1561 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1562 = (N459)? 1'b1 : 
                 (N460)? N1248 : 1'b0;
  assign N1563 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1564 = (N459)? 1'b1 : 
                 (N460)? N1247 : 1'b0;
  assign N1565 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1566 = (N459)? 1'b1 : 
                 (N460)? N1246 : 1'b0;
  assign { N1568, N1567 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1569 = (N459)? 1'b1 : 
                 (N460)? N1245 : 1'b0;
  assign N1570 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1571 = (N459)? 1'b1 : 
                 (N460)? N1244 : 1'b0;
  assign N1572 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1573 = (N459)? 1'b1 : 
                 (N460)? N1243 : 1'b0;
  assign N1574 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1575 = (N459)? 1'b1 : 
                 (N460)? N1242 : 1'b0;
  assign N1576 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1577 = (N459)? 1'b1 : 
                 (N460)? N1241 : 1'b0;
  assign N1578 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1579 = (N459)? 1'b1 : 
                 (N460)? N1240 : 1'b0;
  assign N1580 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1581 = (N459)? 1'b1 : 
                 (N460)? N1239 : 1'b0;
  assign N1582 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1583 = (N459)? 1'b1 : 
                 (N460)? N1238 : 1'b0;
  assign { N1585, N1584 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1586 = (N459)? 1'b1 : 
                 (N460)? N1237 : 1'b0;
  assign N1587 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1588 = (N459)? 1'b1 : 
                 (N460)? N1236 : 1'b0;
  assign N1589 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1590 = (N459)? 1'b1 : 
                 (N460)? N1235 : 1'b0;
  assign N1591 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1592 = (N459)? 1'b1 : 
                 (N460)? N1234 : 1'b0;
  assign N1593 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1594 = (N459)? 1'b1 : 
                 (N460)? N1233 : 1'b0;
  assign N1595 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1596 = (N459)? 1'b1 : 
                 (N460)? N1232 : 1'b0;
  assign N1597 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1598 = (N459)? 1'b1 : 
                 (N460)? N1231 : 1'b0;
  assign N1599 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1600 = (N459)? 1'b1 : 
                 (N460)? N1230 : 1'b0;
  assign N1601 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1602 = (N459)? 1'b1 : 
                 (N460)? N1229 : 1'b0;
  assign N1603 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1604 = (N459)? 1'b1 : 
                 (N460)? N1228 : 1'b0;
  assign N1605 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1606 = (N459)? 1'b1 : 
                 (N460)? N1227 : 1'b0;
  assign N1607 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1608 = (N459)? 1'b1 : 
                 (N460)? N1226 : 1'b0;
  assign N1609 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1610 = (N459)? 1'b1 : 
                 (N460)? N1225 : 1'b0;
  assign N1611 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1612 = (N459)? 1'b1 : 
                 (N460)? N1224 : 1'b0;
  assign N1613 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1614 = (N459)? 1'b1 : 
                 (N460)? N1223 : 1'b0;
  assign N1615 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1616 = (N459)? 1'b1 : 
                 (N460)? N1222 : 1'b0;
  assign { N1618, N1617 } = (N459)? { 1'b0, 1'b0 } : 
                            (N460)? { io_bht_update_bits_taken, T12[0:0] } : 1'b0;
  assign N1619 = (N459)? 1'b1 : 
                 (N460)? N1221 : 1'b0;
  assign N1620 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1621 = (N459)? 1'b1 : 
                 (N460)? N1220 : 1'b0;
  assign N1622 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1623 = (N459)? 1'b1 : 
                 (N460)? N1219 : 1'b0;
  assign N1624 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1625 = (N459)? 1'b1 : 
                 (N460)? N1218 : 1'b0;
  assign N1626 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1627 = (N459)? 1'b1 : 
                 (N460)? N1217 : 1'b0;
  assign N1628 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1629 = (N459)? 1'b1 : 
                 (N460)? N1216 : 1'b0;
  assign N1630 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1631 = (N459)? 1'b1 : 
                 (N460)? N1215 : 1'b0;
  assign N1632 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1633 = (N459)? 1'b1 : 
                 (N460)? N1214 : 1'b0;
  assign N1634 = (N459)? 1'b0 : 
                 (N460)? T12[0] : 1'b0;
  assign N1638 = (N459)? 1'b1 : 
                 (N2307)? 1'b1 : 
                 (N2310)? 1'b1 : 
                 (N1637)? 1'b0 : 1'b0;
  assign { N1645, N1644, N1643, N1642, N1641, N1640, N1639 } = (N459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                               (N2307)? { io_bht_update_bits_taken, io_bht_update_bits_prediction_bits_bht_history[6:1] } : 
                                                               (N2310)? { io_resp_bits_bht_value[0:0], io_resp_bits_bht_history[6:1] } : 1'b0;
  assign N1648 = (N459)? 1'b1 : 
                 (N2312)? 1'b1 : 
                 (N1647)? 1'b0 : 1'b0;
  assign { N1654, N1653, N1652, N1651, N1650, N1649 } = (N459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2312)? T172 : 1'b0;
  assign N1658 = (N459)? 1'b1 : 
                 (N2313)? 1'b1 : 
                 (N2316)? 1'b1 : 
                 (N1657)? 1'b0 : 1'b0;
  assign { N1664, N1663, N1662, N1661, N1660, N1659 } = (N459)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2313)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                        (N2316)? T192 : 1'b0;
  assign N1667 = (N459)? 1'b1 : 
                 (N2317)? 1'b1 : 
                 (N1666)? 1'b0 : 1'b0;
  assign { N1670, N1669, N1668 } = (N459)? { 1'b0, 1'b0, 1'b0 } : 
                                   (N2317)? T200 : 1'b0;
  assign { N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734 } = (N609)? { N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N610)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N609 = T288;
  assign N610 = N1671;
  assign { N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859 } = (N611)? { N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N612)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N611 = T601;
  assign N612 = N1796;
  assign { N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984 } = (N613)? { N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N614)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N613 = T800;
  assign N614 = N1921;
  assign { N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109 } = (N615)? { N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N616)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N615 = T1541;
  assign N616 = N2046;
  assign N2174 = (N459)? 1'b1 : 
                 (N2318)? 1'b1 : 
                 (N2321)? 1'b1 : 
                 (N2173)? 1'b0 : 1'b0;
  assign N2175 = (N459)? 1'b0 : 
                 (N2318)? T2006 : 
                 (N2321)? T2001 : 1'b0;
  assign N2179 = (N459)? 1'b1 : 
                 (N2313)? 1'b1 : 
                 (N2322)? 1'b1 : 
                 (N2324)? 1'b1 : 
                 (N2178)? 1'b0 : 1'b0;
  assign { N2181, N2180 } = (N459)? { 1'b0, 1'b0 } : 
                            (N2313)? { 1'b0, 1'b0 } : 
                            (N2322)? T2017 : 
                            (N2324)? T2014 : 1'b0;
  assign { N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245 } = (N617)? { N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N618)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N617 = T2409;
  assign N618 = N2182;
  assign io_resp_bits_bridx = (N619)? brIdx[0] : 
                              (N620)? brIdx[1] : 
                              (N621)? brIdx[2] : 
                              (N622)? brIdx[3] : 
                              (N623)? brIdx[4] : 
                              (N624)? brIdx[5] : 
                              (N625)? brIdx[6] : 
                              (N626)? brIdx[7] : 
                              (N627)? brIdx[8] : 
                              (N628)? brIdx[9] : 
                              (N629)? brIdx[10] : 
                              (N630)? brIdx[11] : 
                              (N631)? brIdx[12] : 
                              (N632)? brIdx[13] : 
                              (N633)? brIdx[14] : 
                              (N634)? brIdx[15] : 
                              (N635)? brIdx[16] : 
                              (N636)? brIdx[17] : 
                              (N637)? brIdx[18] : 
                              (N638)? brIdx[19] : 
                              (N639)? brIdx[20] : 
                              (N640)? brIdx[21] : 
                              (N641)? brIdx[22] : 
                              (N642)? brIdx[23] : 
                              (N643)? brIdx[24] : 
                              (N644)? brIdx[25] : 
                              (N645)? brIdx[26] : 
                              (N646)? brIdx[27] : 
                              (N647)? brIdx[28] : 
                              (N648)? brIdx[29] : 
                              (N649)? brIdx[30] : 
                              (N650)? brIdx[31] : 
                              (N651)? brIdx[32] : 
                              (N652)? brIdx[33] : 
                              (N653)? brIdx[34] : 
                              (N654)? brIdx[35] : 
                              (N655)? brIdx[36] : 
                              (N656)? brIdx[37] : 
                              (N657)? brIdx[38] : 
                              (N658)? brIdx[39] : 
                              (N659)? brIdx[40] : 
                              (N660)? brIdx[41] : 
                              (N661)? brIdx[42] : 
                              (N662)? brIdx[43] : 
                              (N663)? brIdx[44] : 
                              (N664)? brIdx[45] : 
                              (N665)? brIdx[46] : 
                              (N666)? brIdx[47] : 
                              (N667)? brIdx[48] : 
                              (N668)? brIdx[49] : 
                              (N669)? brIdx[50] : 
                              (N670)? brIdx[51] : 
                              (N671)? brIdx[52] : 
                              (N672)? brIdx[53] : 
                              (N673)? brIdx[54] : 
                              (N674)? brIdx[55] : 
                              (N675)? brIdx[56] : 
                              (N676)? brIdx[57] : 
                              (N677)? brIdx[58] : 
                              (N678)? brIdx[59] : 
                              (N679)? brIdx[60] : 
                              (N680)? brIdx[61] : 1'b0;
  assign N619 = N1020;
  assign N620 = N1022;
  assign N621 = N1024;
  assign N622 = N1026;
  assign N623 = N1028;
  assign N624 = N1030;
  assign N625 = N1032;
  assign N626 = N1034;
  assign N627 = N1036;
  assign N628 = N1038;
  assign N629 = N1040;
  assign N630 = N1042;
  assign N631 = N1044;
  assign N632 = N1046;
  assign N633 = N1048;
  assign N634 = N1050;
  assign N635 = N1052;
  assign N636 = N1054;
  assign N637 = N1056;
  assign N638 = N1058;
  assign N639 = N1060;
  assign N640 = N1062;
  assign N641 = N1064;
  assign N642 = N1066;
  assign N643 = N1068;
  assign N644 = N1070;
  assign N645 = N1072;
  assign N646 = N1074;
  assign N647 = N1076;
  assign N648 = N1078;
  assign N649 = N1080;
  assign N650 = N1081;
  assign N651 = N1021;
  assign N652 = N1023;
  assign N653 = N1025;
  assign N654 = N1027;
  assign N655 = N1029;
  assign N656 = N1031;
  assign N657 = N1033;
  assign N658 = N1035;
  assign N659 = N1037;
  assign N660 = N1039;
  assign N661 = N1041;
  assign N662 = N1043;
  assign N663 = N1045;
  assign N664 = N1047;
  assign N665 = N1049;
  assign N666 = N1051;
  assign N667 = N1053;
  assign N668 = N1055;
  assign N669 = N1057;
  assign N670 = N1059;
  assign N671 = N1061;
  assign N672 = N1063;
  assign N673 = N1065;
  assign N674 = N1067;
  assign N675 = N1069;
  assign N676 = N1071;
  assign N677 = N1073;
  assign N678 = N1075;
  assign N679 = N1077;
  assign N680 = N1079;
  assign N681 = ~T152[0];
  assign N682 = ~T152[1];
  assign N683 = N681 & N682;
  assign N684 = N681 & T152[1];
  assign N685 = T152[0] & N682;
  assign N686 = T152[0] & T152[1];
  assign N687 = ~T152[2];
  assign N688 = N683 & N687;
  assign N689 = N683 & T152[2];
  assign N690 = N685 & N687;
  assign N691 = N685 & T152[2];
  assign N692 = N684 & N687;
  assign N693 = N684 & T152[2];
  assign N694 = N686 & N687;
  assign N695 = N686 & T152[2];
  assign N696 = ~T152[3];
  assign N697 = N688 & N696;
  assign N698 = N688 & T152[3];
  assign N699 = N690 & N696;
  assign N700 = N690 & T152[3];
  assign N701 = N692 & N696;
  assign N702 = N692 & T152[3];
  assign N703 = N694 & N696;
  assign N704 = N694 & T152[3];
  assign N705 = N689 & N696;
  assign N706 = N689 & T152[3];
  assign N707 = N691 & N696;
  assign N708 = N691 & T152[3];
  assign N709 = N693 & N696;
  assign N710 = N693 & T152[3];
  assign N711 = N695 & N696;
  assign N712 = N695 & T152[3];
  assign N713 = ~T152[4];
  assign N714 = N697 & N713;
  assign N715 = N697 & T152[4];
  assign N716 = N699 & N713;
  assign N717 = N699 & T152[4];
  assign N718 = N701 & N713;
  assign N719 = N701 & T152[4];
  assign N720 = N703 & N713;
  assign N721 = N703 & T152[4];
  assign N722 = N705 & N713;
  assign N723 = N705 & T152[4];
  assign N724 = N707 & N713;
  assign N725 = N707 & T152[4];
  assign N726 = N709 & N713;
  assign N727 = N709 & T152[4];
  assign N728 = N711 & N713;
  assign N729 = N711 & T152[4];
  assign N730 = N698 & N713;
  assign N731 = N698 & T152[4];
  assign N732 = N700 & N713;
  assign N733 = N700 & T152[4];
  assign N734 = N702 & N713;
  assign N735 = N702 & T152[4];
  assign N736 = N704 & N713;
  assign N737 = N704 & T152[4];
  assign N738 = N706 & N713;
  assign N739 = N706 & T152[4];
  assign N740 = N708 & N713;
  assign N741 = N708 & T152[4];
  assign N742 = N710 & N713;
  assign N743 = N710 & T152[4];
  assign N744 = N712 & N713;
  assign N745 = N712 & T152[4];
  assign N746 = ~T152[5];
  assign N747 = N714 & N746;
  assign N748 = N714 & T152[5];
  assign N749 = N716 & N746;
  assign N750 = N716 & T152[5];
  assign N751 = N718 & N746;
  assign N752 = N718 & T152[5];
  assign N753 = N720 & N746;
  assign N754 = N720 & T152[5];
  assign N755 = N722 & N746;
  assign N756 = N722 & T152[5];
  assign N757 = N724 & N746;
  assign N758 = N724 & T152[5];
  assign N759 = N726 & N746;
  assign N760 = N726 & T152[5];
  assign N761 = N728 & N746;
  assign N762 = N728 & T152[5];
  assign N763 = N730 & N746;
  assign N764 = N730 & T152[5];
  assign N765 = N732 & N746;
  assign N766 = N732 & T152[5];
  assign N767 = N734 & N746;
  assign N768 = N734 & T152[5];
  assign N769 = N736 & N746;
  assign N770 = N736 & T152[5];
  assign N771 = N738 & N746;
  assign N772 = N738 & T152[5];
  assign N773 = N740 & N746;
  assign N774 = N740 & T152[5];
  assign N775 = N742 & N746;
  assign N776 = N742 & T152[5];
  assign N777 = N744 & N746;
  assign N778 = N744 & T152[5];
  assign N779 = N715 & N746;
  assign N780 = N715 & T152[5];
  assign N781 = N717 & N746;
  assign N782 = N717 & T152[5];
  assign N783 = N719 & N746;
  assign N784 = N719 & T152[5];
  assign N785 = N721 & N746;
  assign N786 = N721 & T152[5];
  assign N787 = N723 & N746;
  assign N788 = N723 & T152[5];
  assign N789 = N725 & N746;
  assign N790 = N725 & T152[5];
  assign N791 = N727 & N746;
  assign N792 = N727 & T152[5];
  assign N793 = N729 & N746;
  assign N794 = N729 & T152[5];
  assign N795 = N731 & N746;
  assign N796 = N731 & T152[5];
  assign N797 = N733 & N746;
  assign N798 = N733 & T152[5];
  assign N799 = N735 & N746;
  assign N800 = N735 & T152[5];
  assign N801 = N737 & N746;
  assign N802 = N737 & T152[5];
  assign N803 = N739 & N746;
  assign N804 = N739 & T152[5];
  assign N805 = N741 & N746;
  assign N806 = N741 & T152[5];
  assign N807 = N743 & N746;
  assign N808 = N743 & T152[5];
  assign N809 = N745 & N746;
  assign N810 = N745 & T152[5];
  assign N811 = ~T152[6];
  assign N812 = N747 & N811;
  assign N813 = N747 & T152[6];
  assign N814 = N749 & N811;
  assign N815 = N749 & T152[6];
  assign N816 = N751 & N811;
  assign N817 = N751 & T152[6];
  assign N818 = N753 & N811;
  assign N819 = N753 & T152[6];
  assign N820 = N755 & N811;
  assign N821 = N755 & T152[6];
  assign N822 = N757 & N811;
  assign N823 = N757 & T152[6];
  assign N824 = N759 & N811;
  assign N825 = N759 & T152[6];
  assign N826 = N761 & N811;
  assign N827 = N761 & T152[6];
  assign N828 = N763 & N811;
  assign N829 = N763 & T152[6];
  assign N830 = N765 & N811;
  assign N831 = N765 & T152[6];
  assign N832 = N767 & N811;
  assign N833 = N767 & T152[6];
  assign N834 = N769 & N811;
  assign N835 = N769 & T152[6];
  assign N836 = N771 & N811;
  assign N837 = N771 & T152[6];
  assign N838 = N773 & N811;
  assign N839 = N773 & T152[6];
  assign N840 = N775 & N811;
  assign N841 = N775 & T152[6];
  assign N842 = N777 & N811;
  assign N843 = N777 & T152[6];
  assign N844 = N779 & N811;
  assign N845 = N779 & T152[6];
  assign N846 = N781 & N811;
  assign N847 = N781 & T152[6];
  assign N848 = N783 & N811;
  assign N849 = N783 & T152[6];
  assign N850 = N785 & N811;
  assign N851 = N785 & T152[6];
  assign N852 = N787 & N811;
  assign N853 = N787 & T152[6];
  assign N854 = N789 & N811;
  assign N855 = N789 & T152[6];
  assign N856 = N791 & N811;
  assign N857 = N791 & T152[6];
  assign N858 = N793 & N811;
  assign N859 = N793 & T152[6];
  assign N860 = N795 & N811;
  assign N861 = N795 & T152[6];
  assign N862 = N797 & N811;
  assign N863 = N797 & T152[6];
  assign N864 = N799 & N811;
  assign N865 = N799 & T152[6];
  assign N866 = N801 & N811;
  assign N867 = N801 & T152[6];
  assign N868 = N803 & N811;
  assign N869 = N803 & T152[6];
  assign N870 = N805 & N811;
  assign N871 = N805 & T152[6];
  assign N872 = N807 & N811;
  assign N873 = N807 & T152[6];
  assign N874 = N809 & N811;
  assign N875 = N809 & T152[6];
  assign N876 = N748 & N811;
  assign N877 = N748 & T152[6];
  assign N878 = N750 & N811;
  assign N879 = N750 & T152[6];
  assign N880 = N752 & N811;
  assign N881 = N752 & T152[6];
  assign N882 = N754 & N811;
  assign N883 = N754 & T152[6];
  assign N884 = N756 & N811;
  assign N885 = N756 & T152[6];
  assign N886 = N758 & N811;
  assign N887 = N758 & T152[6];
  assign N888 = N760 & N811;
  assign N889 = N760 & T152[6];
  assign N890 = N762 & N811;
  assign N891 = N762 & T152[6];
  assign N892 = N764 & N811;
  assign N893 = N764 & T152[6];
  assign N894 = N766 & N811;
  assign N895 = N766 & T152[6];
  assign N896 = N768 & N811;
  assign N897 = N768 & T152[6];
  assign N898 = N770 & N811;
  assign N899 = N770 & T152[6];
  assign N900 = N772 & N811;
  assign N901 = N772 & T152[6];
  assign N902 = N774 & N811;
  assign N903 = N774 & T152[6];
  assign N904 = N776 & N811;
  assign N905 = N776 & T152[6];
  assign N906 = N778 & N811;
  assign N907 = N778 & T152[6];
  assign N908 = N780 & N811;
  assign N909 = N780 & T152[6];
  assign N910 = N782 & N811;
  assign N911 = N782 & T152[6];
  assign N912 = N784 & N811;
  assign N913 = N784 & T152[6];
  assign N914 = N786 & N811;
  assign N915 = N786 & T152[6];
  assign N916 = N788 & N811;
  assign N917 = N788 & T152[6];
  assign N918 = N790 & N811;
  assign N919 = N790 & T152[6];
  assign N920 = N792 & N811;
  assign N921 = N792 & T152[6];
  assign N922 = N794 & N811;
  assign N923 = N794 & T152[6];
  assign N924 = N796 & N811;
  assign N925 = N796 & T152[6];
  assign N926 = N798 & N811;
  assign N927 = N798 & T152[6];
  assign N928 = N800 & N811;
  assign N929 = N800 & T152[6];
  assign N930 = N802 & N811;
  assign N931 = N802 & T152[6];
  assign N932 = N804 & N811;
  assign N933 = N804 & T152[6];
  assign N934 = N806 & N811;
  assign N935 = N806 & T152[6];
  assign N936 = N808 & N811;
  assign N937 = N808 & T152[6];
  assign N938 = N810 & N811;
  assign N939 = N810 & T152[6];
  assign T12[0] = T18 | T14;
  assign T14 = T15 & io_bht_update_bits_taken;
  assign T15 = io_bht_update_bits_prediction_bits_bht_value[1] | io_bht_update_bits_prediction_bits_bht_value[0];
  assign T18 = io_bht_update_bits_prediction_bits_bht_value[1] & io_bht_update_bits_prediction_bits_bht_value[0];
  assign T21 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T22[6] = io_bht_update_bits_pc[8] ^ io_bht_update_bits_prediction_bits_bht_history[6];
  assign T22[5] = io_bht_update_bits_pc[7] ^ io_bht_update_bits_prediction_bits_bht_history[5];
  assign T22[4] = io_bht_update_bits_pc[6] ^ io_bht_update_bits_prediction_bits_bht_history[4];
  assign T22[3] = io_bht_update_bits_pc[5] ^ io_bht_update_bits_prediction_bits_bht_history[3];
  assign T22[2] = io_bht_update_bits_pc[4] ^ io_bht_update_bits_prediction_bits_bht_history[2];
  assign T22[1] = io_bht_update_bits_pc[3] ^ io_bht_update_bits_prediction_bits_bht_history[1];
  assign T22[0] = io_bht_update_bits_pc[2] ^ io_bht_update_bits_prediction_bits_bht_history[0];
  assign T152[6] = io_req_bits_addr[8] ^ io_resp_bits_bht_history[6];
  assign T152[5] = io_req_bits_addr[7] ^ io_resp_bits_bht_history[5];
  assign T152[4] = io_req_bits_addr[6] ^ io_resp_bits_bht_history[4];
  assign T152[3] = io_req_bits_addr[5] ^ io_resp_bits_bht_history[3];
  assign T152[2] = io_req_bits_addr[4] ^ io_resp_bits_bht_history[2];
  assign T152[1] = io_req_bits_addr[3] ^ io_resp_bits_bht_history[1];
  assign T152[0] = io_req_bits_addr[2] ^ io_resp_bits_bht_history[0];
  assign T159 = T1527 & T160;
  assign T160 = ~T161;
  assign T161 = T1162 | T162;
  assign N940 = ~hits[61];
  assign T166 = R7 & T168[61];
  assign N941 = ~updateHit;
  assign T175 = R7 & T176;
  assign T176 = ~updateHit;
  assign hits[61] = T589[61] & N2784;
  assign hits[60] = T589[60] & N2794;
  assign hits[59] = T589[59] & N2799;
  assign hits[58] = T589[58] & N2804;
  assign hits[57] = T589[57] & N2809;
  assign hits[56] = T589[56] & N2814;
  assign hits[55] = T589[55] & N2819;
  assign hits[54] = T589[54] & N2824;
  assign hits[53] = T589[53] & N2834;
  assign hits[52] = T589[52] & N2839;
  assign hits[51] = T589[51] & N2844;
  assign hits[50] = T589[50] & N2849;
  assign hits[49] = T589[49] & N2854;
  assign hits[48] = T589[48] & N2859;
  assign hits[47] = T589[47] & N2864;
  assign hits[46] = T589[46] & N2869;
  assign hits[45] = T589[45] & N2874;
  assign hits[44] = T589[44] & N2879;
  assign hits[43] = T589[43] & N2884;
  assign hits[42] = T589[42] & N2889;
  assign hits[41] = T589[41] & N2894;
  assign hits[40] = T589[40] & N2899;
  assign hits[39] = T589[39] & N2904;
  assign hits[38] = T589[38] & N2909;
  assign hits[37] = T589[37] & N2914;
  assign hits[36] = T589[36] & N2919;
  assign hits[35] = T589[35] & N2924;
  assign hits[34] = T589[34] & N2929;
  assign hits[33] = T589[33] & N2934;
  assign hits[32] = T589[32] & N2939;
  assign hits[31] = T589[31] & N2944;
  assign hits[30] = T589[30] & N2949;
  assign hits[29] = T589[29] & N2954;
  assign hits[28] = T589[28] & N2959;
  assign hits[27] = T589[27] & N2964;
  assign hits[26] = T589[26] & N2969;
  assign hits[25] = T589[25] & N2974;
  assign hits[24] = T589[24] & N2979;
  assign hits[23] = T589[23] & N2984;
  assign hits[22] = T589[22] & N2989;
  assign hits[21] = T589[21] & N2994;
  assign hits[20] = T589[20] & N2999;
  assign hits[19] = T589[19] & N3004;
  assign hits[18] = T589[18] & N3009;
  assign hits[17] = T589[17] & N3014;
  assign hits[16] = T589[16] & N3019;
  assign hits[15] = T589[15] & N3024;
  assign hits[14] = T589[14] & N3029;
  assign hits[13] = T589[13] & N3034;
  assign hits[12] = T589[12] & N3039;
  assign hits[11] = T589[11] & N3044;
  assign hits[10] = T589[10] & N3049;
  assign hits[9] = T589[9] & N3054;
  assign hits[8] = T589[8] & N3059;
  assign hits[7] = T589[7] & N3064;
  assign hits[6] = T589[6] & N3069;
  assign hits[5] = T589[5] & N3074;
  assign hits[4] = T589[4] & N3079;
  assign hits[3] = T589[3] & N3084;
  assign hits[2] = T589[2] & N3089;
  assign hits[1] = T589[1] & N3099;
  assign hits[0] = T589[0] & N3094;
  assign T189[5] = idxPagesOH_0[5] & pageHit[5];
  assign T189[4] = idxPagesOH_0[4] & pageHit[4];
  assign T189[3] = idxPagesOH_0[3] & pageHit[3];
  assign T189[2] = idxPagesOH_0[2] & pageHit[2];
  assign T189[1] = idxPagesOH_0[1] & pageHit[1];
  assign T189[0] = idxPagesOH_0[0] & pageHit[0];
  assign pageHit[5] = T266[5] & pageValid[5];
  assign pageHit[4] = T266[4] & pageValid[4];
  assign pageHit[3] = T266[3] & pageValid[3];
  assign pageHit[2] = T266[2] & pageValid[2];
  assign pageHit[1] = T266[1] & pageValid[1];
  assign pageHit[0] = T266[0] & pageValid[0];
  assign T192[5] = pageValid[5] | pageReplEn[5];
  assign T192[4] = pageValid[4] | pageReplEn[4];
  assign T192[3] = pageValid[3] | pageReplEn[3];
  assign T192[2] = pageValid[2] | pageReplEn[2];
  assign T192[1] = pageValid[1] | pageReplEn[1];
  assign T192[0] = pageValid[0] | pageReplEn[0];
  assign pageReplEn[5] = idxPageReplEn[5] | tgtPageReplEn[5];
  assign pageReplEn[4] = idxPageReplEn[4] | tgtPageReplEn[4];
  assign pageReplEn[3] = idxPageReplEn[3] | tgtPageReplEn[3];
  assign pageReplEn[2] = idxPageReplEn[2] | tgtPageReplEn[2];
  assign pageReplEn[1] = idxPageReplEn[1] | tgtPageReplEn[1];
  assign pageReplEn[0] = idxPageReplEn[0] | tgtPageReplEn[0];
  assign N942 = ~doTgtPageRepl;
  assign N943 = ~samePage;
  assign T193[5] = T195[5] | 1'b0;
  assign T193[4] = T195[4] | 1'b0;
  assign T193[3] = T195[3] | 1'b0;
  assign T193[2] = T195[2] | 1'b0;
  assign T193[1] = T195[1] | 1'b0;
  assign T193[0] = 1'b0 | T2420[0];
  assign N944 = ~N2829;
  assign T203 = R7 & doPageRepl;
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign doIdxPageRepl = ~N2829;
  assign updatePageHit[5] = T204[5] & pageValid[5];
  assign updatePageHit[4] = T204[4] & pageValid[4];
  assign updatePageHit[3] = T204[3] & pageValid[3];
  assign updatePageHit[2] = T204[2] & pageValid[2];
  assign updatePageHit[1] = T204[1] & pageValid[1];
  assign updatePageHit[0] = T204[0] & pageValid[0];
  assign N945 = ~N2779;
  assign T219 = R7 & T220;
  assign T220 = T222 & pageReplEn[5];
  assign T224 = R7 & T225;
  assign T225 = T222 & pageReplEn[3];
  assign T228 = R7 & T229;
  assign T229 = T222 & pageReplEn[1];
  assign T235 = R7 & T236;
  assign T236 = T238 & pageReplEn[4];
  assign T240 = R7 & T241;
  assign T241 = T238 & pageReplEn[2];
  assign T244 = R7 & T245;
  assign T245 = T238 & pageReplEn[0];
  assign doTgtPageRepl = T264 & T261;
  assign T261 = ~N2789;
  assign T262[5] = pageHit[5] & T263[5];
  assign T262[4] = pageHit[4] & T263[4];
  assign T262[3] = pageHit[3] & T263[3];
  assign T262[2] = pageHit[2] & T263[2];
  assign T262[1] = pageHit[1] & T263[1];
  assign T262[0] = pageHit[0] & T263[0];
  assign T263[5] = ~idxPageReplEn[5];
  assign T263[4] = ~idxPageReplEn[4];
  assign T263[3] = ~idxPageReplEn[3];
  assign T263[2] = ~idxPageReplEn[2];
  assign T263[1] = ~idxPageReplEn[1];
  assign T263[0] = ~idxPageReplEn[0];
  assign T264 = ~samePage;
  assign N946 = ~doIdxPageRepl;
  assign T265 = R7 & doPageRepl;
  assign T2423[0] = T195[4] | T2427[1];
  assign T2427[1] = T2420[0] | T195[2];
  assign T288 = R7 & T289;
  assign T291[5] = idxPagesOH_1[5] & pageHit[5];
  assign T291[4] = idxPagesOH_1[4] & pageHit[4];
  assign T291[3] = idxPagesOH_1[3] & pageHit[3];
  assign T291[2] = idxPagesOH_1[2] & pageHit[2];
  assign T291[1] = idxPagesOH_1[1] & pageHit[1];
  assign T291[0] = idxPagesOH_1[0] & pageHit[0];
  assign T296[5] = idxPagesOH_2[5] & pageHit[5];
  assign T296[4] = idxPagesOH_2[4] & pageHit[4];
  assign T296[3] = idxPagesOH_2[3] & pageHit[3];
  assign T296[2] = idxPagesOH_2[2] & pageHit[2];
  assign T296[1] = idxPagesOH_2[1] & pageHit[1];
  assign T296[0] = idxPagesOH_2[0] & pageHit[0];
  assign T300[5] = idxPagesOH_3[5] & pageHit[5];
  assign T300[4] = idxPagesOH_3[4] & pageHit[4];
  assign T300[3] = idxPagesOH_3[3] & pageHit[3];
  assign T300[2] = idxPagesOH_3[2] & pageHit[2];
  assign T300[1] = idxPagesOH_3[1] & pageHit[1];
  assign T300[0] = idxPagesOH_3[0] & pageHit[0];
  assign T306[5] = idxPagesOH_4[5] & pageHit[5];
  assign T306[4] = idxPagesOH_4[4] & pageHit[4];
  assign T306[3] = idxPagesOH_4[3] & pageHit[3];
  assign T306[2] = idxPagesOH_4[2] & pageHit[2];
  assign T306[1] = idxPagesOH_4[1] & pageHit[1];
  assign T306[0] = idxPagesOH_4[0] & pageHit[0];
  assign T310[5] = idxPagesOH_5[5] & pageHit[5];
  assign T310[4] = idxPagesOH_5[4] & pageHit[4];
  assign T310[3] = idxPagesOH_5[3] & pageHit[3];
  assign T310[2] = idxPagesOH_5[2] & pageHit[2];
  assign T310[1] = idxPagesOH_5[1] & pageHit[1];
  assign T310[0] = idxPagesOH_5[0] & pageHit[0];
  assign T315[5] = idxPagesOH_6[5] & pageHit[5];
  assign T315[4] = idxPagesOH_6[4] & pageHit[4];
  assign T315[3] = idxPagesOH_6[3] & pageHit[3];
  assign T315[2] = idxPagesOH_6[2] & pageHit[2];
  assign T315[1] = idxPagesOH_6[1] & pageHit[1];
  assign T315[0] = idxPagesOH_6[0] & pageHit[0];
  assign T319[5] = idxPagesOH_7[5] & pageHit[5];
  assign T319[4] = idxPagesOH_7[4] & pageHit[4];
  assign T319[3] = idxPagesOH_7[3] & pageHit[3];
  assign T319[2] = idxPagesOH_7[2] & pageHit[2];
  assign T319[1] = idxPagesOH_7[1] & pageHit[1];
  assign T319[0] = idxPagesOH_7[0] & pageHit[0];
  assign T326[5] = idxPagesOH_8[5] & pageHit[5];
  assign T326[4] = idxPagesOH_8[4] & pageHit[4];
  assign T326[3] = idxPagesOH_8[3] & pageHit[3];
  assign T326[2] = idxPagesOH_8[2] & pageHit[2];
  assign T326[1] = idxPagesOH_8[1] & pageHit[1];
  assign T326[0] = idxPagesOH_8[0] & pageHit[0];
  assign T330[5] = idxPagesOH_9[5] & pageHit[5];
  assign T330[4] = idxPagesOH_9[4] & pageHit[4];
  assign T330[3] = idxPagesOH_9[3] & pageHit[3];
  assign T330[2] = idxPagesOH_9[2] & pageHit[2];
  assign T330[1] = idxPagesOH_9[1] & pageHit[1];
  assign T330[0] = idxPagesOH_9[0] & pageHit[0];
  assign T335[5] = idxPagesOH_10[5] & pageHit[5];
  assign T335[4] = idxPagesOH_10[4] & pageHit[4];
  assign T335[3] = idxPagesOH_10[3] & pageHit[3];
  assign T335[2] = idxPagesOH_10[2] & pageHit[2];
  assign T335[1] = idxPagesOH_10[1] & pageHit[1];
  assign T335[0] = idxPagesOH_10[0] & pageHit[0];
  assign T339[5] = idxPagesOH_11[5] & pageHit[5];
  assign T339[4] = idxPagesOH_11[4] & pageHit[4];
  assign T339[3] = idxPagesOH_11[3] & pageHit[3];
  assign T339[2] = idxPagesOH_11[2] & pageHit[2];
  assign T339[1] = idxPagesOH_11[1] & pageHit[1];
  assign T339[0] = idxPagesOH_11[0] & pageHit[0];
  assign T345[5] = idxPagesOH_12[5] & pageHit[5];
  assign T345[4] = idxPagesOH_12[4] & pageHit[4];
  assign T345[3] = idxPagesOH_12[3] & pageHit[3];
  assign T345[2] = idxPagesOH_12[2] & pageHit[2];
  assign T345[1] = idxPagesOH_12[1] & pageHit[1];
  assign T345[0] = idxPagesOH_12[0] & pageHit[0];
  assign T349[5] = idxPagesOH_13[5] & pageHit[5];
  assign T349[4] = idxPagesOH_13[4] & pageHit[4];
  assign T349[3] = idxPagesOH_13[3] & pageHit[3];
  assign T349[2] = idxPagesOH_13[2] & pageHit[2];
  assign T349[1] = idxPagesOH_13[1] & pageHit[1];
  assign T349[0] = idxPagesOH_13[0] & pageHit[0];
  assign T354[5] = idxPagesOH_14[5] & pageHit[5];
  assign T354[4] = idxPagesOH_14[4] & pageHit[4];
  assign T354[3] = idxPagesOH_14[3] & pageHit[3];
  assign T354[2] = idxPagesOH_14[2] & pageHit[2];
  assign T354[1] = idxPagesOH_14[1] & pageHit[1];
  assign T354[0] = idxPagesOH_14[0] & pageHit[0];
  assign T358[5] = idxPagesOH_15[5] & pageHit[5];
  assign T358[4] = idxPagesOH_15[4] & pageHit[4];
  assign T358[3] = idxPagesOH_15[3] & pageHit[3];
  assign T358[2] = idxPagesOH_15[2] & pageHit[2];
  assign T358[1] = idxPagesOH_15[1] & pageHit[1];
  assign T358[0] = idxPagesOH_15[0] & pageHit[0];
  assign T366[5] = idxPagesOH_16[5] & pageHit[5];
  assign T366[4] = idxPagesOH_16[4] & pageHit[4];
  assign T366[3] = idxPagesOH_16[3] & pageHit[3];
  assign T366[2] = idxPagesOH_16[2] & pageHit[2];
  assign T366[1] = idxPagesOH_16[1] & pageHit[1];
  assign T366[0] = idxPagesOH_16[0] & pageHit[0];
  assign T370[5] = idxPagesOH_17[5] & pageHit[5];
  assign T370[4] = idxPagesOH_17[4] & pageHit[4];
  assign T370[3] = idxPagesOH_17[3] & pageHit[3];
  assign T370[2] = idxPagesOH_17[2] & pageHit[2];
  assign T370[1] = idxPagesOH_17[1] & pageHit[1];
  assign T370[0] = idxPagesOH_17[0] & pageHit[0];
  assign T375[5] = idxPagesOH_18[5] & pageHit[5];
  assign T375[4] = idxPagesOH_18[4] & pageHit[4];
  assign T375[3] = idxPagesOH_18[3] & pageHit[3];
  assign T375[2] = idxPagesOH_18[2] & pageHit[2];
  assign T375[1] = idxPagesOH_18[1] & pageHit[1];
  assign T375[0] = idxPagesOH_18[0] & pageHit[0];
  assign T379[5] = idxPagesOH_19[5] & pageHit[5];
  assign T379[4] = idxPagesOH_19[4] & pageHit[4];
  assign T379[3] = idxPagesOH_19[3] & pageHit[3];
  assign T379[2] = idxPagesOH_19[2] & pageHit[2];
  assign T379[1] = idxPagesOH_19[1] & pageHit[1];
  assign T379[0] = idxPagesOH_19[0] & pageHit[0];
  assign T385[5] = idxPagesOH_20[5] & pageHit[5];
  assign T385[4] = idxPagesOH_20[4] & pageHit[4];
  assign T385[3] = idxPagesOH_20[3] & pageHit[3];
  assign T385[2] = idxPagesOH_20[2] & pageHit[2];
  assign T385[1] = idxPagesOH_20[1] & pageHit[1];
  assign T385[0] = idxPagesOH_20[0] & pageHit[0];
  assign T389[5] = idxPagesOH_21[5] & pageHit[5];
  assign T389[4] = idxPagesOH_21[4] & pageHit[4];
  assign T389[3] = idxPagesOH_21[3] & pageHit[3];
  assign T389[2] = idxPagesOH_21[2] & pageHit[2];
  assign T389[1] = idxPagesOH_21[1] & pageHit[1];
  assign T389[0] = idxPagesOH_21[0] & pageHit[0];
  assign T394[5] = idxPagesOH_22[5] & pageHit[5];
  assign T394[4] = idxPagesOH_22[4] & pageHit[4];
  assign T394[3] = idxPagesOH_22[3] & pageHit[3];
  assign T394[2] = idxPagesOH_22[2] & pageHit[2];
  assign T394[1] = idxPagesOH_22[1] & pageHit[1];
  assign T394[0] = idxPagesOH_22[0] & pageHit[0];
  assign T398[5] = idxPagesOH_23[5] & pageHit[5];
  assign T398[4] = idxPagesOH_23[4] & pageHit[4];
  assign T398[3] = idxPagesOH_23[3] & pageHit[3];
  assign T398[2] = idxPagesOH_23[2] & pageHit[2];
  assign T398[1] = idxPagesOH_23[1] & pageHit[1];
  assign T398[0] = idxPagesOH_23[0] & pageHit[0];
  assign T405[5] = idxPagesOH_24[5] & pageHit[5];
  assign T405[4] = idxPagesOH_24[4] & pageHit[4];
  assign T405[3] = idxPagesOH_24[3] & pageHit[3];
  assign T405[2] = idxPagesOH_24[2] & pageHit[2];
  assign T405[1] = idxPagesOH_24[1] & pageHit[1];
  assign T405[0] = idxPagesOH_24[0] & pageHit[0];
  assign T409[5] = idxPagesOH_25[5] & pageHit[5];
  assign T409[4] = idxPagesOH_25[4] & pageHit[4];
  assign T409[3] = idxPagesOH_25[3] & pageHit[3];
  assign T409[2] = idxPagesOH_25[2] & pageHit[2];
  assign T409[1] = idxPagesOH_25[1] & pageHit[1];
  assign T409[0] = idxPagesOH_25[0] & pageHit[0];
  assign T414[5] = idxPagesOH_26[5] & pageHit[5];
  assign T414[4] = idxPagesOH_26[4] & pageHit[4];
  assign T414[3] = idxPagesOH_26[3] & pageHit[3];
  assign T414[2] = idxPagesOH_26[2] & pageHit[2];
  assign T414[1] = idxPagesOH_26[1] & pageHit[1];
  assign T414[0] = idxPagesOH_26[0] & pageHit[0];
  assign T418[5] = idxPagesOH_27[5] & pageHit[5];
  assign T418[4] = idxPagesOH_27[4] & pageHit[4];
  assign T418[3] = idxPagesOH_27[3] & pageHit[3];
  assign T418[2] = idxPagesOH_27[2] & pageHit[2];
  assign T418[1] = idxPagesOH_27[1] & pageHit[1];
  assign T418[0] = idxPagesOH_27[0] & pageHit[0];
  assign T424[5] = idxPagesOH_28[5] & pageHit[5];
  assign T424[4] = idxPagesOH_28[4] & pageHit[4];
  assign T424[3] = idxPagesOH_28[3] & pageHit[3];
  assign T424[2] = idxPagesOH_28[2] & pageHit[2];
  assign T424[1] = idxPagesOH_28[1] & pageHit[1];
  assign T424[0] = idxPagesOH_28[0] & pageHit[0];
  assign T428[5] = idxPagesOH_29[5] & pageHit[5];
  assign T428[4] = idxPagesOH_29[4] & pageHit[4];
  assign T428[3] = idxPagesOH_29[3] & pageHit[3];
  assign T428[2] = idxPagesOH_29[2] & pageHit[2];
  assign T428[1] = idxPagesOH_29[1] & pageHit[1];
  assign T428[0] = idxPagesOH_29[0] & pageHit[0];
  assign T432[5] = idxPagesOH_30[5] & pageHit[5];
  assign T432[4] = idxPagesOH_30[4] & pageHit[4];
  assign T432[3] = idxPagesOH_30[3] & pageHit[3];
  assign T432[2] = idxPagesOH_30[2] & pageHit[2];
  assign T432[1] = idxPagesOH_30[1] & pageHit[1];
  assign T432[0] = idxPagesOH_30[0] & pageHit[0];
  assign T441[5] = idxPagesOH_31[5] & pageHit[5];
  assign T441[4] = idxPagesOH_31[4] & pageHit[4];
  assign T441[3] = idxPagesOH_31[3] & pageHit[3];
  assign T441[2] = idxPagesOH_31[2] & pageHit[2];
  assign T441[1] = idxPagesOH_31[1] & pageHit[1];
  assign T441[0] = idxPagesOH_31[0] & pageHit[0];
  assign T445[5] = idxPagesOH_32[5] & pageHit[5];
  assign T445[4] = idxPagesOH_32[4] & pageHit[4];
  assign T445[3] = idxPagesOH_32[3] & pageHit[3];
  assign T445[2] = idxPagesOH_32[2] & pageHit[2];
  assign T445[1] = idxPagesOH_32[1] & pageHit[1];
  assign T445[0] = idxPagesOH_32[0] & pageHit[0];
  assign T450[5] = idxPagesOH_33[5] & pageHit[5];
  assign T450[4] = idxPagesOH_33[4] & pageHit[4];
  assign T450[3] = idxPagesOH_33[3] & pageHit[3];
  assign T450[2] = idxPagesOH_33[2] & pageHit[2];
  assign T450[1] = idxPagesOH_33[1] & pageHit[1];
  assign T450[0] = idxPagesOH_33[0] & pageHit[0];
  assign T454[5] = idxPagesOH_34[5] & pageHit[5];
  assign T454[4] = idxPagesOH_34[4] & pageHit[4];
  assign T454[3] = idxPagesOH_34[3] & pageHit[3];
  assign T454[2] = idxPagesOH_34[2] & pageHit[2];
  assign T454[1] = idxPagesOH_34[1] & pageHit[1];
  assign T454[0] = idxPagesOH_34[0] & pageHit[0];
  assign T460[5] = idxPagesOH_35[5] & pageHit[5];
  assign T460[4] = idxPagesOH_35[4] & pageHit[4];
  assign T460[3] = idxPagesOH_35[3] & pageHit[3];
  assign T460[2] = idxPagesOH_35[2] & pageHit[2];
  assign T460[1] = idxPagesOH_35[1] & pageHit[1];
  assign T460[0] = idxPagesOH_35[0] & pageHit[0];
  assign T464[5] = idxPagesOH_36[5] & pageHit[5];
  assign T464[4] = idxPagesOH_36[4] & pageHit[4];
  assign T464[3] = idxPagesOH_36[3] & pageHit[3];
  assign T464[2] = idxPagesOH_36[2] & pageHit[2];
  assign T464[1] = idxPagesOH_36[1] & pageHit[1];
  assign T464[0] = idxPagesOH_36[0] & pageHit[0];
  assign T469[5] = idxPagesOH_37[5] & pageHit[5];
  assign T469[4] = idxPagesOH_37[4] & pageHit[4];
  assign T469[3] = idxPagesOH_37[3] & pageHit[3];
  assign T469[2] = idxPagesOH_37[2] & pageHit[2];
  assign T469[1] = idxPagesOH_37[1] & pageHit[1];
  assign T469[0] = idxPagesOH_37[0] & pageHit[0];
  assign T473[5] = idxPagesOH_38[5] & pageHit[5];
  assign T473[4] = idxPagesOH_38[4] & pageHit[4];
  assign T473[3] = idxPagesOH_38[3] & pageHit[3];
  assign T473[2] = idxPagesOH_38[2] & pageHit[2];
  assign T473[1] = idxPagesOH_38[1] & pageHit[1];
  assign T473[0] = idxPagesOH_38[0] & pageHit[0];
  assign T480[5] = idxPagesOH_39[5] & pageHit[5];
  assign T480[4] = idxPagesOH_39[4] & pageHit[4];
  assign T480[3] = idxPagesOH_39[3] & pageHit[3];
  assign T480[2] = idxPagesOH_39[2] & pageHit[2];
  assign T480[1] = idxPagesOH_39[1] & pageHit[1];
  assign T480[0] = idxPagesOH_39[0] & pageHit[0];
  assign T484[5] = idxPagesOH_40[5] & pageHit[5];
  assign T484[4] = idxPagesOH_40[4] & pageHit[4];
  assign T484[3] = idxPagesOH_40[3] & pageHit[3];
  assign T484[2] = idxPagesOH_40[2] & pageHit[2];
  assign T484[1] = idxPagesOH_40[1] & pageHit[1];
  assign T484[0] = idxPagesOH_40[0] & pageHit[0];
  assign T489[5] = idxPagesOH_41[5] & pageHit[5];
  assign T489[4] = idxPagesOH_41[4] & pageHit[4];
  assign T489[3] = idxPagesOH_41[3] & pageHit[3];
  assign T489[2] = idxPagesOH_41[2] & pageHit[2];
  assign T489[1] = idxPagesOH_41[1] & pageHit[1];
  assign T489[0] = idxPagesOH_41[0] & pageHit[0];
  assign T493[5] = idxPagesOH_42[5] & pageHit[5];
  assign T493[4] = idxPagesOH_42[4] & pageHit[4];
  assign T493[3] = idxPagesOH_42[3] & pageHit[3];
  assign T493[2] = idxPagesOH_42[2] & pageHit[2];
  assign T493[1] = idxPagesOH_42[1] & pageHit[1];
  assign T493[0] = idxPagesOH_42[0] & pageHit[0];
  assign T499[5] = idxPagesOH_43[5] & pageHit[5];
  assign T499[4] = idxPagesOH_43[4] & pageHit[4];
  assign T499[3] = idxPagesOH_43[3] & pageHit[3];
  assign T499[2] = idxPagesOH_43[2] & pageHit[2];
  assign T499[1] = idxPagesOH_43[1] & pageHit[1];
  assign T499[0] = idxPagesOH_43[0] & pageHit[0];
  assign T503[5] = idxPagesOH_44[5] & pageHit[5];
  assign T503[4] = idxPagesOH_44[4] & pageHit[4];
  assign T503[3] = idxPagesOH_44[3] & pageHit[3];
  assign T503[2] = idxPagesOH_44[2] & pageHit[2];
  assign T503[1] = idxPagesOH_44[1] & pageHit[1];
  assign T503[0] = idxPagesOH_44[0] & pageHit[0];
  assign T508[5] = idxPagesOH_45[5] & pageHit[5];
  assign T508[4] = idxPagesOH_45[4] & pageHit[4];
  assign T508[3] = idxPagesOH_45[3] & pageHit[3];
  assign T508[2] = idxPagesOH_45[2] & pageHit[2];
  assign T508[1] = idxPagesOH_45[1] & pageHit[1];
  assign T508[0] = idxPagesOH_45[0] & pageHit[0];
  assign T512[5] = idxPagesOH_46[5] & pageHit[5];
  assign T512[4] = idxPagesOH_46[4] & pageHit[4];
  assign T512[3] = idxPagesOH_46[3] & pageHit[3];
  assign T512[2] = idxPagesOH_46[2] & pageHit[2];
  assign T512[1] = idxPagesOH_46[1] & pageHit[1];
  assign T512[0] = idxPagesOH_46[0] & pageHit[0];
  assign T520[5] = idxPagesOH_47[5] & pageHit[5];
  assign T520[4] = idxPagesOH_47[4] & pageHit[4];
  assign T520[3] = idxPagesOH_47[3] & pageHit[3];
  assign T520[2] = idxPagesOH_47[2] & pageHit[2];
  assign T520[1] = idxPagesOH_47[1] & pageHit[1];
  assign T520[0] = idxPagesOH_47[0] & pageHit[0];
  assign T524[5] = idxPagesOH_48[5] & pageHit[5];
  assign T524[4] = idxPagesOH_48[4] & pageHit[4];
  assign T524[3] = idxPagesOH_48[3] & pageHit[3];
  assign T524[2] = idxPagesOH_48[2] & pageHit[2];
  assign T524[1] = idxPagesOH_48[1] & pageHit[1];
  assign T524[0] = idxPagesOH_48[0] & pageHit[0];
  assign T529[5] = idxPagesOH_49[5] & pageHit[5];
  assign T529[4] = idxPagesOH_49[4] & pageHit[4];
  assign T529[3] = idxPagesOH_49[3] & pageHit[3];
  assign T529[2] = idxPagesOH_49[2] & pageHit[2];
  assign T529[1] = idxPagesOH_49[1] & pageHit[1];
  assign T529[0] = idxPagesOH_49[0] & pageHit[0];
  assign T533[5] = idxPagesOH_50[5] & pageHit[5];
  assign T533[4] = idxPagesOH_50[4] & pageHit[4];
  assign T533[3] = idxPagesOH_50[3] & pageHit[3];
  assign T533[2] = idxPagesOH_50[2] & pageHit[2];
  assign T533[1] = idxPagesOH_50[1] & pageHit[1];
  assign T533[0] = idxPagesOH_50[0] & pageHit[0];
  assign T539[5] = idxPagesOH_51[5] & pageHit[5];
  assign T539[4] = idxPagesOH_51[4] & pageHit[4];
  assign T539[3] = idxPagesOH_51[3] & pageHit[3];
  assign T539[2] = idxPagesOH_51[2] & pageHit[2];
  assign T539[1] = idxPagesOH_51[1] & pageHit[1];
  assign T539[0] = idxPagesOH_51[0] & pageHit[0];
  assign T543[5] = idxPagesOH_52[5] & pageHit[5];
  assign T543[4] = idxPagesOH_52[4] & pageHit[4];
  assign T543[3] = idxPagesOH_52[3] & pageHit[3];
  assign T543[2] = idxPagesOH_52[2] & pageHit[2];
  assign T543[1] = idxPagesOH_52[1] & pageHit[1];
  assign T543[0] = idxPagesOH_52[0] & pageHit[0];
  assign T548[5] = idxPagesOH_53[5] & pageHit[5];
  assign T548[4] = idxPagesOH_53[4] & pageHit[4];
  assign T548[3] = idxPagesOH_53[3] & pageHit[3];
  assign T548[2] = idxPagesOH_53[2] & pageHit[2];
  assign T548[1] = idxPagesOH_53[1] & pageHit[1];
  assign T548[0] = idxPagesOH_53[0] & pageHit[0];
  assign T552[5] = idxPagesOH_54[5] & pageHit[5];
  assign T552[4] = idxPagesOH_54[4] & pageHit[4];
  assign T552[3] = idxPagesOH_54[3] & pageHit[3];
  assign T552[2] = idxPagesOH_54[2] & pageHit[2];
  assign T552[1] = idxPagesOH_54[1] & pageHit[1];
  assign T552[0] = idxPagesOH_54[0] & pageHit[0];
  assign T559[5] = idxPagesOH_55[5] & pageHit[5];
  assign T559[4] = idxPagesOH_55[4] & pageHit[4];
  assign T559[3] = idxPagesOH_55[3] & pageHit[3];
  assign T559[2] = idxPagesOH_55[2] & pageHit[2];
  assign T559[1] = idxPagesOH_55[1] & pageHit[1];
  assign T559[0] = idxPagesOH_55[0] & pageHit[0];
  assign T563[5] = idxPagesOH_56[5] & pageHit[5];
  assign T563[4] = idxPagesOH_56[4] & pageHit[4];
  assign T563[3] = idxPagesOH_56[3] & pageHit[3];
  assign T563[2] = idxPagesOH_56[2] & pageHit[2];
  assign T563[1] = idxPagesOH_56[1] & pageHit[1];
  assign T563[0] = idxPagesOH_56[0] & pageHit[0];
  assign T568[5] = idxPagesOH_57[5] & pageHit[5];
  assign T568[4] = idxPagesOH_57[4] & pageHit[4];
  assign T568[3] = idxPagesOH_57[3] & pageHit[3];
  assign T568[2] = idxPagesOH_57[2] & pageHit[2];
  assign T568[1] = idxPagesOH_57[1] & pageHit[1];
  assign T568[0] = idxPagesOH_57[0] & pageHit[0];
  assign T572[5] = idxPagesOH_58[5] & pageHit[5];
  assign T572[4] = idxPagesOH_58[4] & pageHit[4];
  assign T572[3] = idxPagesOH_58[3] & pageHit[3];
  assign T572[2] = idxPagesOH_58[2] & pageHit[2];
  assign T572[1] = idxPagesOH_58[1] & pageHit[1];
  assign T572[0] = idxPagesOH_58[0] & pageHit[0];
  assign T578[5] = idxPagesOH_59[5] & pageHit[5];
  assign T578[4] = idxPagesOH_59[4] & pageHit[4];
  assign T578[3] = idxPagesOH_59[3] & pageHit[3];
  assign T578[2] = idxPagesOH_59[2] & pageHit[2];
  assign T578[1] = idxPagesOH_59[1] & pageHit[1];
  assign T578[0] = idxPagesOH_59[0] & pageHit[0];
  assign T582[5] = idxPagesOH_60[5] & pageHit[5];
  assign T582[4] = idxPagesOH_60[4] & pageHit[4];
  assign T582[3] = idxPagesOH_60[3] & pageHit[3];
  assign T582[2] = idxPagesOH_60[2] & pageHit[2];
  assign T582[1] = idxPagesOH_60[1] & pageHit[1];
  assign T582[0] = idxPagesOH_60[0] & pageHit[0];
  assign T586[5] = idxPagesOH_61[5] & pageHit[5];
  assign T586[4] = idxPagesOH_61[4] & pageHit[4];
  assign T586[3] = idxPagesOH_61[3] & pageHit[3];
  assign T586[2] = idxPagesOH_61[2] & pageHit[2];
  assign T586[1] = idxPagesOH_61[1] & pageHit[1];
  assign T586[0] = idxPagesOH_61[0] & pageHit[0];
  assign T589[61] = T2437[61] & T590[61];
  assign T589[60] = T2437[60] & T590[60];
  assign T589[59] = T2437[59] & T590[59];
  assign T589[58] = T2437[58] & T590[58];
  assign T589[57] = T2437[57] & T590[57];
  assign T589[56] = T2437[56] & T590[56];
  assign T589[55] = T2437[55] & T590[55];
  assign T589[54] = T2437[54] & T590[54];
  assign T589[53] = T2437[53] & T590[53];
  assign T589[52] = T2437[52] & T590[52];
  assign T589[51] = T2437[51] & T590[51];
  assign T589[50] = T2437[50] & T590[50];
  assign T589[49] = T2437[49] & T590[49];
  assign T589[48] = T2437[48] & T590[48];
  assign T589[47] = T2437[47] & T590[47];
  assign T589[46] = T2437[46] & T590[46];
  assign T589[45] = T2437[45] & T590[45];
  assign T589[44] = T2437[44] & T590[44];
  assign T589[43] = T2437[43] & T590[43];
  assign T589[42] = T2437[42] & T590[42];
  assign T589[41] = T2437[41] & T590[41];
  assign T589[40] = T2437[40] & T590[40];
  assign T589[39] = T2437[39] & T590[39];
  assign T589[38] = T2437[38] & T590[38];
  assign T589[37] = T2437[37] & T590[37];
  assign T589[36] = T2437[36] & T590[36];
  assign T589[35] = T2437[35] & T590[35];
  assign T589[34] = T2437[34] & T590[34];
  assign T589[33] = T2437[33] & T590[33];
  assign T589[32] = T2437[32] & T590[32];
  assign T589[31] = T2437[31] & T590[31];
  assign T589[30] = T2437[30] & T590[30];
  assign T589[29] = T2437[29] & T590[29];
  assign T589[28] = T2437[28] & T590[28];
  assign T589[27] = T2437[27] & T590[27];
  assign T589[26] = T2437[26] & T590[26];
  assign T589[25] = T2437[25] & T590[25];
  assign T589[24] = T2437[24] & T590[24];
  assign T589[23] = T2437[23] & T590[23];
  assign T589[22] = T2437[22] & T590[22];
  assign T589[21] = T2437[21] & T590[21];
  assign T589[20] = T2437[20] & T590[20];
  assign T589[19] = T2437[19] & T590[19];
  assign T589[18] = T2437[18] & T590[18];
  assign T589[17] = T2437[17] & T590[17];
  assign T589[16] = T2437[16] & T590[16];
  assign T589[15] = T2437[15] & T590[15];
  assign T589[14] = T2437[14] & T590[14];
  assign T589[13] = T2437[13] & T590[13];
  assign T589[12] = T2437[12] & T590[12];
  assign T589[11] = T2437[11] & T590[11];
  assign T589[10] = T2437[10] & T590[10];
  assign T589[9] = T2437[9] & T590[9];
  assign T589[8] = T2437[8] & T590[8];
  assign T589[7] = T2437[7] & T590[7];
  assign T589[6] = T2437[6] & T590[6];
  assign T589[5] = T2437[5] & T590[5];
  assign T589[4] = T2437[4] & T590[4];
  assign T589[3] = T2437[3] & T590[3];
  assign T589[2] = T2437[2] & T590[2];
  assign T589[1] = T2437[1] & T590[1];
  assign T589[0] = T2437[0] & T590[0];
  assign T601 = R7 & T602;
  assign N947 = ~io_invalidate;
  assign N948 = ~R7;
  assign T782[61] = T2438[61] | T783[61];
  assign T782[60] = T2438[60] | T783[60];
  assign T782[59] = T2438[59] | T783[59];
  assign T782[58] = T2438[58] | T783[58];
  assign T782[57] = T2438[57] | T783[57];
  assign T782[56] = T2438[56] | T783[56];
  assign T782[55] = T2438[55] | T783[55];
  assign T782[54] = T2438[54] | T783[54];
  assign T782[53] = T2438[53] | T783[53];
  assign T782[52] = T2438[52] | T783[52];
  assign T782[51] = T2438[51] | T783[51];
  assign T782[50] = T2438[50] | T783[50];
  assign T782[49] = T2438[49] | T783[49];
  assign T782[48] = T2438[48] | T783[48];
  assign T782[47] = T2438[47] | T783[47];
  assign T782[46] = T2438[46] | T783[46];
  assign T782[45] = T2438[45] | T783[45];
  assign T782[44] = T2438[44] | T783[44];
  assign T782[43] = T2438[43] | T783[43];
  assign T782[42] = T2438[42] | T783[42];
  assign T782[41] = T2438[41] | T783[41];
  assign T782[40] = T2438[40] | T783[40];
  assign T782[39] = T2438[39] | T783[39];
  assign T782[38] = T2438[38] | T783[38];
  assign T782[37] = T2438[37] | T783[37];
  assign T782[36] = T2438[36] | T783[36];
  assign T782[35] = T2438[35] | T783[35];
  assign T782[34] = T2438[34] | T783[34];
  assign T782[33] = T2438[33] | T783[33];
  assign T782[32] = T2438[32] | T783[32];
  assign T782[31] = T2438[31] | T783[31];
  assign T782[30] = T2438[30] | T783[30];
  assign T782[29] = T2438[29] | T783[29];
  assign T782[28] = T2438[28] | T783[28];
  assign T782[27] = T2438[27] | T783[27];
  assign T782[26] = T2438[26] | T783[26];
  assign T782[25] = T2438[25] | T783[25];
  assign T782[24] = T2438[24] | T783[24];
  assign T782[23] = T2438[23] | T783[23];
  assign T782[22] = T2438[22] | T783[22];
  assign T782[21] = T2438[21] | T783[21];
  assign T782[20] = T2438[20] | T783[20];
  assign T782[19] = T2438[19] | T783[19];
  assign T782[18] = T2438[18] | T783[18];
  assign T782[17] = T2438[17] | T783[17];
  assign T782[16] = T2438[16] | T783[16];
  assign T782[15] = T2438[15] | T783[15];
  assign T782[14] = T2438[14] | T783[14];
  assign T782[13] = T2438[13] | T783[13];
  assign T782[12] = T2438[12] | T783[12];
  assign T782[11] = T2438[11] | T783[11];
  assign T782[10] = T2438[10] | T783[10];
  assign T782[9] = T2438[9] | T783[9];
  assign T782[8] = T2438[8] | T783[8];
  assign T782[7] = T2438[7] | T783[7];
  assign T782[6] = T2438[6] | T783[6];
  assign T782[5] = T2438[5] | T783[5];
  assign T782[4] = T2438[4] | T783[4];
  assign T782[3] = T2438[3] | T783[3];
  assign T782[2] = T2438[2] | T783[2];
  assign T782[1] = T2438[1] | T783[1];
  assign T782[0] = T2438[0] | T783[0];
  assign T2438[61] = T2437[61] & T785[61];
  assign T2438[60] = T2437[60] & T785[60];
  assign T2438[59] = T2437[59] & T785[59];
  assign T2438[58] = T2437[58] & T785[58];
  assign T2438[57] = T2437[57] & T785[57];
  assign T2438[56] = T2437[56] & T785[56];
  assign T2438[55] = T2437[55] & T785[55];
  assign T2438[54] = T2437[54] & T785[54];
  assign T2438[53] = T2437[53] & T785[53];
  assign T2438[52] = T2437[52] & T785[52];
  assign T2438[51] = T2437[51] & T785[51];
  assign T2438[50] = T2437[50] & T785[50];
  assign T2438[49] = T2437[49] & T785[49];
  assign T2438[48] = T2437[48] & T785[48];
  assign T2438[47] = T2437[47] & T785[47];
  assign T2438[46] = T2437[46] & T785[46];
  assign T2438[45] = T2437[45] & T785[45];
  assign T2438[44] = T2437[44] & T785[44];
  assign T2438[43] = T2437[43] & T785[43];
  assign T2438[42] = T2437[42] & T785[42];
  assign T2438[41] = T2437[41] & T785[41];
  assign T2438[40] = T2437[40] & T785[40];
  assign T2438[39] = T2437[39] & T785[39];
  assign T2438[38] = T2437[38] & T785[38];
  assign T2438[37] = T2437[37] & T785[37];
  assign T2438[36] = T2437[36] & T785[36];
  assign T2438[35] = T2437[35] & T785[35];
  assign T2438[34] = T2437[34] & T785[34];
  assign T2438[33] = T2437[33] & T785[33];
  assign T2438[32] = T2437[32] & T785[32];
  assign T2438[31] = T2437[31] & T785[31];
  assign T2438[30] = T2437[30] & T785[30];
  assign T2438[29] = T2437[29] & T785[29];
  assign T2438[28] = T2437[28] & T785[28];
  assign T2438[27] = T2437[27] & T785[27];
  assign T2438[26] = T2437[26] & T785[26];
  assign T2438[25] = T2437[25] & T785[25];
  assign T2438[24] = T2437[24] & T785[24];
  assign T2438[23] = T2437[23] & T785[23];
  assign T2438[22] = T2437[22] & T785[22];
  assign T2438[21] = T2437[21] & T785[21];
  assign T2438[20] = T2437[20] & T785[20];
  assign T2438[19] = T2437[19] & T785[19];
  assign T2438[18] = T2437[18] & T785[18];
  assign T2438[17] = T2437[17] & T785[17];
  assign T2438[16] = T2437[16] & T785[16];
  assign T2438[15] = T2437[15] & T785[15];
  assign T2438[14] = T2437[14] & T785[14];
  assign T2438[13] = T2437[13] & T785[13];
  assign T2438[12] = T2437[12] & T785[12];
  assign T2438[11] = T2437[11] & T785[11];
  assign T2438[10] = T2437[10] & T785[10];
  assign T2438[9] = T2437[9] & T785[9];
  assign T2438[8] = T2437[8] & T785[8];
  assign T2438[7] = T2437[7] & T785[7];
  assign T2438[6] = T2437[6] & T785[6];
  assign T2438[5] = T2437[5] & T785[5];
  assign T2438[4] = T2437[4] & T785[4];
  assign T2438[3] = T2437[3] & T785[3];
  assign T2438[2] = T2437[2] & T785[2];
  assign T2438[1] = T2437[1] & T785[1];
  assign T2438[0] = T2437[0] & T785[0];
  assign T785[61] = ~N2470;
  assign T785[60] = ~N2475;
  assign T785[59] = ~N2480;
  assign T785[58] = ~N2485;
  assign T785[57] = ~N2490;
  assign T785[56] = ~N2495;
  assign T785[55] = ~N2500;
  assign T785[54] = ~N2505;
  assign T785[53] = ~N2510;
  assign T785[52] = ~N2515;
  assign T785[51] = ~N2520;
  assign T785[50] = ~N2525;
  assign T785[49] = ~N2530;
  assign T785[48] = ~N2535;
  assign T785[47] = ~N2540;
  assign T785[46] = ~N2545;
  assign T785[45] = ~N2550;
  assign T785[44] = ~N2555;
  assign T785[43] = ~N2560;
  assign T785[42] = ~N2565;
  assign T785[41] = ~N2570;
  assign T785[40] = ~N2575;
  assign T785[39] = ~N2580;
  assign T785[38] = ~N2585;
  assign T785[37] = ~N2590;
  assign T785[36] = ~N2595;
  assign T785[35] = ~N2600;
  assign T785[34] = ~N2605;
  assign T785[33] = ~N2610;
  assign T785[32] = ~N2615;
  assign T785[31] = ~N2620;
  assign T785[30] = ~N2625;
  assign T785[29] = ~N2630;
  assign T785[28] = ~N2635;
  assign T785[27] = ~N2640;
  assign T785[26] = ~N2645;
  assign T785[25] = ~N2650;
  assign T785[24] = ~N2655;
  assign T785[23] = ~N2660;
  assign T785[22] = ~N2665;
  assign T785[21] = ~N2670;
  assign T785[20] = ~N2675;
  assign T785[19] = ~N2680;
  assign T785[18] = ~N2685;
  assign T785[17] = ~N2690;
  assign T785[16] = ~N2695;
  assign T785[15] = ~N2700;
  assign T785[14] = ~N2705;
  assign T785[13] = ~N2710;
  assign T785[12] = ~N2715;
  assign T785[11] = ~N2720;
  assign T785[10] = ~N2725;
  assign T785[9] = ~N2730;
  assign T785[8] = ~N2735;
  assign T785[7] = ~N2740;
  assign T785[6] = ~N2745;
  assign T785[5] = ~N2750;
  assign T785[4] = ~N2755;
  assign T785[3] = ~N2760;
  assign T785[2] = ~N2765;
  assign T785[1] = ~N2770;
  assign T785[0] = ~N2775;
  assign T794[5] = pageReplEn[5] & T795[5];
  assign T794[4] = pageReplEn[4] & T795[4];
  assign T794[3] = pageReplEn[3] & T795[3];
  assign T794[2] = pageReplEn[2] & T795[2];
  assign T794[1] = pageReplEn[1] & T795[1];
  assign T794[0] = pageReplEn[0] & T795[0];
  assign T795[5] = idxPagesOH_0[5] | tgtPagesOH_0[5];
  assign T795[4] = idxPagesOH_0[4] | tgtPagesOH_0[4];
  assign T795[3] = idxPagesOH_0[3] | tgtPagesOH_0[3];
  assign T795[2] = idxPagesOH_0[2] | tgtPagesOH_0[2];
  assign T795[1] = idxPagesOH_0[1] | tgtPagesOH_0[1];
  assign T795[0] = idxPagesOH_0[0] | tgtPagesOH_0[0];
  assign T2439[0] = T2444[3] | T2443[1];
  assign T2443[1] = T799[5] | T2445[1];
  assign N949 = ~N2789;
  assign T800 = R7 & T801;
  assign T803[5] = pageReplEn[5] & T804[5];
  assign T803[4] = pageReplEn[4] & T804[4];
  assign T803[3] = pageReplEn[3] & T804[3];
  assign T803[2] = pageReplEn[2] & T804[2];
  assign T803[1] = pageReplEn[1] & T804[1];
  assign T803[0] = pageReplEn[0] & T804[0];
  assign T804[5] = idxPagesOH_1[5] | tgtPagesOH_1[5];
  assign T804[4] = idxPagesOH_1[4] | tgtPagesOH_1[4];
  assign T804[3] = idxPagesOH_1[3] | tgtPagesOH_1[3];
  assign T804[2] = idxPagesOH_1[2] | tgtPagesOH_1[2];
  assign T804[1] = idxPagesOH_1[1] | tgtPagesOH_1[1];
  assign T804[0] = idxPagesOH_1[0] | tgtPagesOH_1[0];
  assign T809[5] = pageReplEn[5] & T810[5];
  assign T809[4] = pageReplEn[4] & T810[4];
  assign T809[3] = pageReplEn[3] & T810[3];
  assign T809[2] = pageReplEn[2] & T810[2];
  assign T809[1] = pageReplEn[1] & T810[1];
  assign T809[0] = pageReplEn[0] & T810[0];
  assign T810[5] = idxPagesOH_2[5] | tgtPagesOH_2[5];
  assign T810[4] = idxPagesOH_2[4] | tgtPagesOH_2[4];
  assign T810[3] = idxPagesOH_2[3] | tgtPagesOH_2[3];
  assign T810[2] = idxPagesOH_2[2] | tgtPagesOH_2[2];
  assign T810[1] = idxPagesOH_2[1] | tgtPagesOH_2[1];
  assign T810[0] = idxPagesOH_2[0] | tgtPagesOH_2[0];
  assign T814[5] = pageReplEn[5] & T815[5];
  assign T814[4] = pageReplEn[4] & T815[4];
  assign T814[3] = pageReplEn[3] & T815[3];
  assign T814[2] = pageReplEn[2] & T815[2];
  assign T814[1] = pageReplEn[1] & T815[1];
  assign T814[0] = pageReplEn[0] & T815[0];
  assign T815[5] = idxPagesOH_3[5] | tgtPagesOH_3[5];
  assign T815[4] = idxPagesOH_3[4] | tgtPagesOH_3[4];
  assign T815[3] = idxPagesOH_3[3] | tgtPagesOH_3[3];
  assign T815[2] = idxPagesOH_3[2] | tgtPagesOH_3[2];
  assign T815[1] = idxPagesOH_3[1] | tgtPagesOH_3[1];
  assign T815[0] = idxPagesOH_3[0] | tgtPagesOH_3[0];
  assign T821[5] = pageReplEn[5] & T822[5];
  assign T821[4] = pageReplEn[4] & T822[4];
  assign T821[3] = pageReplEn[3] & T822[3];
  assign T821[2] = pageReplEn[2] & T822[2];
  assign T821[1] = pageReplEn[1] & T822[1];
  assign T821[0] = pageReplEn[0] & T822[0];
  assign T822[5] = idxPagesOH_4[5] | tgtPagesOH_4[5];
  assign T822[4] = idxPagesOH_4[4] | tgtPagesOH_4[4];
  assign T822[3] = idxPagesOH_4[3] | tgtPagesOH_4[3];
  assign T822[2] = idxPagesOH_4[2] | tgtPagesOH_4[2];
  assign T822[1] = idxPagesOH_4[1] | tgtPagesOH_4[1];
  assign T822[0] = idxPagesOH_4[0] | tgtPagesOH_4[0];
  assign T826[5] = pageReplEn[5] & T827[5];
  assign T826[4] = pageReplEn[4] & T827[4];
  assign T826[3] = pageReplEn[3] & T827[3];
  assign T826[2] = pageReplEn[2] & T827[2];
  assign T826[1] = pageReplEn[1] & T827[1];
  assign T826[0] = pageReplEn[0] & T827[0];
  assign T827[5] = idxPagesOH_5[5] | tgtPagesOH_5[5];
  assign T827[4] = idxPagesOH_5[4] | tgtPagesOH_5[4];
  assign T827[3] = idxPagesOH_5[3] | tgtPagesOH_5[3];
  assign T827[2] = idxPagesOH_5[2] | tgtPagesOH_5[2];
  assign T827[1] = idxPagesOH_5[1] | tgtPagesOH_5[1];
  assign T827[0] = idxPagesOH_5[0] | tgtPagesOH_5[0];
  assign T832[5] = pageReplEn[5] & T833[5];
  assign T832[4] = pageReplEn[4] & T833[4];
  assign T832[3] = pageReplEn[3] & T833[3];
  assign T832[2] = pageReplEn[2] & T833[2];
  assign T832[1] = pageReplEn[1] & T833[1];
  assign T832[0] = pageReplEn[0] & T833[0];
  assign T833[5] = idxPagesOH_6[5] | tgtPagesOH_6[5];
  assign T833[4] = idxPagesOH_6[4] | tgtPagesOH_6[4];
  assign T833[3] = idxPagesOH_6[3] | tgtPagesOH_6[3];
  assign T833[2] = idxPagesOH_6[2] | tgtPagesOH_6[2];
  assign T833[1] = idxPagesOH_6[1] | tgtPagesOH_6[1];
  assign T833[0] = idxPagesOH_6[0] | tgtPagesOH_6[0];
  assign T837[5] = pageReplEn[5] & T838[5];
  assign T837[4] = pageReplEn[4] & T838[4];
  assign T837[3] = pageReplEn[3] & T838[3];
  assign T837[2] = pageReplEn[2] & T838[2];
  assign T837[1] = pageReplEn[1] & T838[1];
  assign T837[0] = pageReplEn[0] & T838[0];
  assign T838[5] = idxPagesOH_7[5] | tgtPagesOH_7[5];
  assign T838[4] = idxPagesOH_7[4] | tgtPagesOH_7[4];
  assign T838[3] = idxPagesOH_7[3] | tgtPagesOH_7[3];
  assign T838[2] = idxPagesOH_7[2] | tgtPagesOH_7[2];
  assign T838[1] = idxPagesOH_7[1] | tgtPagesOH_7[1];
  assign T838[0] = idxPagesOH_7[0] | tgtPagesOH_7[0];
  assign T845[5] = pageReplEn[5] & T846[5];
  assign T845[4] = pageReplEn[4] & T846[4];
  assign T845[3] = pageReplEn[3] & T846[3];
  assign T845[2] = pageReplEn[2] & T846[2];
  assign T845[1] = pageReplEn[1] & T846[1];
  assign T845[0] = pageReplEn[0] & T846[0];
  assign T846[5] = idxPagesOH_8[5] | tgtPagesOH_8[5];
  assign T846[4] = idxPagesOH_8[4] | tgtPagesOH_8[4];
  assign T846[3] = idxPagesOH_8[3] | tgtPagesOH_8[3];
  assign T846[2] = idxPagesOH_8[2] | tgtPagesOH_8[2];
  assign T846[1] = idxPagesOH_8[1] | tgtPagesOH_8[1];
  assign T846[0] = idxPagesOH_8[0] | tgtPagesOH_8[0];
  assign T850[5] = pageReplEn[5] & T851[5];
  assign T850[4] = pageReplEn[4] & T851[4];
  assign T850[3] = pageReplEn[3] & T851[3];
  assign T850[2] = pageReplEn[2] & T851[2];
  assign T850[1] = pageReplEn[1] & T851[1];
  assign T850[0] = pageReplEn[0] & T851[0];
  assign T851[5] = idxPagesOH_9[5] | tgtPagesOH_9[5];
  assign T851[4] = idxPagesOH_9[4] | tgtPagesOH_9[4];
  assign T851[3] = idxPagesOH_9[3] | tgtPagesOH_9[3];
  assign T851[2] = idxPagesOH_9[2] | tgtPagesOH_9[2];
  assign T851[1] = idxPagesOH_9[1] | tgtPagesOH_9[1];
  assign T851[0] = idxPagesOH_9[0] | tgtPagesOH_9[0];
  assign T856[5] = pageReplEn[5] & T857[5];
  assign T856[4] = pageReplEn[4] & T857[4];
  assign T856[3] = pageReplEn[3] & T857[3];
  assign T856[2] = pageReplEn[2] & T857[2];
  assign T856[1] = pageReplEn[1] & T857[1];
  assign T856[0] = pageReplEn[0] & T857[0];
  assign T857[5] = idxPagesOH_10[5] | tgtPagesOH_10[5];
  assign T857[4] = idxPagesOH_10[4] | tgtPagesOH_10[4];
  assign T857[3] = idxPagesOH_10[3] | tgtPagesOH_10[3];
  assign T857[2] = idxPagesOH_10[2] | tgtPagesOH_10[2];
  assign T857[1] = idxPagesOH_10[1] | tgtPagesOH_10[1];
  assign T857[0] = idxPagesOH_10[0] | tgtPagesOH_10[0];
  assign T861[5] = pageReplEn[5] & T862[5];
  assign T861[4] = pageReplEn[4] & T862[4];
  assign T861[3] = pageReplEn[3] & T862[3];
  assign T861[2] = pageReplEn[2] & T862[2];
  assign T861[1] = pageReplEn[1] & T862[1];
  assign T861[0] = pageReplEn[0] & T862[0];
  assign T862[5] = idxPagesOH_11[5] | tgtPagesOH_11[5];
  assign T862[4] = idxPagesOH_11[4] | tgtPagesOH_11[4];
  assign T862[3] = idxPagesOH_11[3] | tgtPagesOH_11[3];
  assign T862[2] = idxPagesOH_11[2] | tgtPagesOH_11[2];
  assign T862[1] = idxPagesOH_11[1] | tgtPagesOH_11[1];
  assign T862[0] = idxPagesOH_11[0] | tgtPagesOH_11[0];
  assign T868[5] = pageReplEn[5] & T869[5];
  assign T868[4] = pageReplEn[4] & T869[4];
  assign T868[3] = pageReplEn[3] & T869[3];
  assign T868[2] = pageReplEn[2] & T869[2];
  assign T868[1] = pageReplEn[1] & T869[1];
  assign T868[0] = pageReplEn[0] & T869[0];
  assign T869[5] = idxPagesOH_12[5] | tgtPagesOH_12[5];
  assign T869[4] = idxPagesOH_12[4] | tgtPagesOH_12[4];
  assign T869[3] = idxPagesOH_12[3] | tgtPagesOH_12[3];
  assign T869[2] = idxPagesOH_12[2] | tgtPagesOH_12[2];
  assign T869[1] = idxPagesOH_12[1] | tgtPagesOH_12[1];
  assign T869[0] = idxPagesOH_12[0] | tgtPagesOH_12[0];
  assign T873[5] = pageReplEn[5] & T874[5];
  assign T873[4] = pageReplEn[4] & T874[4];
  assign T873[3] = pageReplEn[3] & T874[3];
  assign T873[2] = pageReplEn[2] & T874[2];
  assign T873[1] = pageReplEn[1] & T874[1];
  assign T873[0] = pageReplEn[0] & T874[0];
  assign T874[5] = idxPagesOH_13[5] | tgtPagesOH_13[5];
  assign T874[4] = idxPagesOH_13[4] | tgtPagesOH_13[4];
  assign T874[3] = idxPagesOH_13[3] | tgtPagesOH_13[3];
  assign T874[2] = idxPagesOH_13[2] | tgtPagesOH_13[2];
  assign T874[1] = idxPagesOH_13[1] | tgtPagesOH_13[1];
  assign T874[0] = idxPagesOH_13[0] | tgtPagesOH_13[0];
  assign T879[5] = pageReplEn[5] & T880[5];
  assign T879[4] = pageReplEn[4] & T880[4];
  assign T879[3] = pageReplEn[3] & T880[3];
  assign T879[2] = pageReplEn[2] & T880[2];
  assign T879[1] = pageReplEn[1] & T880[1];
  assign T879[0] = pageReplEn[0] & T880[0];
  assign T880[5] = idxPagesOH_14[5] | tgtPagesOH_14[5];
  assign T880[4] = idxPagesOH_14[4] | tgtPagesOH_14[4];
  assign T880[3] = idxPagesOH_14[3] | tgtPagesOH_14[3];
  assign T880[2] = idxPagesOH_14[2] | tgtPagesOH_14[2];
  assign T880[1] = idxPagesOH_14[1] | tgtPagesOH_14[1];
  assign T880[0] = idxPagesOH_14[0] | tgtPagesOH_14[0];
  assign T884[5] = pageReplEn[5] & T885[5];
  assign T884[4] = pageReplEn[4] & T885[4];
  assign T884[3] = pageReplEn[3] & T885[3];
  assign T884[2] = pageReplEn[2] & T885[2];
  assign T884[1] = pageReplEn[1] & T885[1];
  assign T884[0] = pageReplEn[0] & T885[0];
  assign T885[5] = idxPagesOH_15[5] | tgtPagesOH_15[5];
  assign T885[4] = idxPagesOH_15[4] | tgtPagesOH_15[4];
  assign T885[3] = idxPagesOH_15[3] | tgtPagesOH_15[3];
  assign T885[2] = idxPagesOH_15[2] | tgtPagesOH_15[2];
  assign T885[1] = idxPagesOH_15[1] | tgtPagesOH_15[1];
  assign T885[0] = idxPagesOH_15[0] | tgtPagesOH_15[0];
  assign T893[5] = pageReplEn[5] & T894[5];
  assign T893[4] = pageReplEn[4] & T894[4];
  assign T893[3] = pageReplEn[3] & T894[3];
  assign T893[2] = pageReplEn[2] & T894[2];
  assign T893[1] = pageReplEn[1] & T894[1];
  assign T893[0] = pageReplEn[0] & T894[0];
  assign T894[5] = idxPagesOH_16[5] | tgtPagesOH_16[5];
  assign T894[4] = idxPagesOH_16[4] | tgtPagesOH_16[4];
  assign T894[3] = idxPagesOH_16[3] | tgtPagesOH_16[3];
  assign T894[2] = idxPagesOH_16[2] | tgtPagesOH_16[2];
  assign T894[1] = idxPagesOH_16[1] | tgtPagesOH_16[1];
  assign T894[0] = idxPagesOH_16[0] | tgtPagesOH_16[0];
  assign T898[5] = pageReplEn[5] & T899[5];
  assign T898[4] = pageReplEn[4] & T899[4];
  assign T898[3] = pageReplEn[3] & T899[3];
  assign T898[2] = pageReplEn[2] & T899[2];
  assign T898[1] = pageReplEn[1] & T899[1];
  assign T898[0] = pageReplEn[0] & T899[0];
  assign T899[5] = idxPagesOH_17[5] | tgtPagesOH_17[5];
  assign T899[4] = idxPagesOH_17[4] | tgtPagesOH_17[4];
  assign T899[3] = idxPagesOH_17[3] | tgtPagesOH_17[3];
  assign T899[2] = idxPagesOH_17[2] | tgtPagesOH_17[2];
  assign T899[1] = idxPagesOH_17[1] | tgtPagesOH_17[1];
  assign T899[0] = idxPagesOH_17[0] | tgtPagesOH_17[0];
  assign T904[5] = pageReplEn[5] & T905[5];
  assign T904[4] = pageReplEn[4] & T905[4];
  assign T904[3] = pageReplEn[3] & T905[3];
  assign T904[2] = pageReplEn[2] & T905[2];
  assign T904[1] = pageReplEn[1] & T905[1];
  assign T904[0] = pageReplEn[0] & T905[0];
  assign T905[5] = idxPagesOH_18[5] | tgtPagesOH_18[5];
  assign T905[4] = idxPagesOH_18[4] | tgtPagesOH_18[4];
  assign T905[3] = idxPagesOH_18[3] | tgtPagesOH_18[3];
  assign T905[2] = idxPagesOH_18[2] | tgtPagesOH_18[2];
  assign T905[1] = idxPagesOH_18[1] | tgtPagesOH_18[1];
  assign T905[0] = idxPagesOH_18[0] | tgtPagesOH_18[0];
  assign T909[5] = pageReplEn[5] & T910[5];
  assign T909[4] = pageReplEn[4] & T910[4];
  assign T909[3] = pageReplEn[3] & T910[3];
  assign T909[2] = pageReplEn[2] & T910[2];
  assign T909[1] = pageReplEn[1] & T910[1];
  assign T909[0] = pageReplEn[0] & T910[0];
  assign T910[5] = idxPagesOH_19[5] | tgtPagesOH_19[5];
  assign T910[4] = idxPagesOH_19[4] | tgtPagesOH_19[4];
  assign T910[3] = idxPagesOH_19[3] | tgtPagesOH_19[3];
  assign T910[2] = idxPagesOH_19[2] | tgtPagesOH_19[2];
  assign T910[1] = idxPagesOH_19[1] | tgtPagesOH_19[1];
  assign T910[0] = idxPagesOH_19[0] | tgtPagesOH_19[0];
  assign T916[5] = pageReplEn[5] & T917[5];
  assign T916[4] = pageReplEn[4] & T917[4];
  assign T916[3] = pageReplEn[3] & T917[3];
  assign T916[2] = pageReplEn[2] & T917[2];
  assign T916[1] = pageReplEn[1] & T917[1];
  assign T916[0] = pageReplEn[0] & T917[0];
  assign T917[5] = idxPagesOH_20[5] | tgtPagesOH_20[5];
  assign T917[4] = idxPagesOH_20[4] | tgtPagesOH_20[4];
  assign T917[3] = idxPagesOH_20[3] | tgtPagesOH_20[3];
  assign T917[2] = idxPagesOH_20[2] | tgtPagesOH_20[2];
  assign T917[1] = idxPagesOH_20[1] | tgtPagesOH_20[1];
  assign T917[0] = idxPagesOH_20[0] | tgtPagesOH_20[0];
  assign T921[5] = pageReplEn[5] & T922[5];
  assign T921[4] = pageReplEn[4] & T922[4];
  assign T921[3] = pageReplEn[3] & T922[3];
  assign T921[2] = pageReplEn[2] & T922[2];
  assign T921[1] = pageReplEn[1] & T922[1];
  assign T921[0] = pageReplEn[0] & T922[0];
  assign T922[5] = idxPagesOH_21[5] | tgtPagesOH_21[5];
  assign T922[4] = idxPagesOH_21[4] | tgtPagesOH_21[4];
  assign T922[3] = idxPagesOH_21[3] | tgtPagesOH_21[3];
  assign T922[2] = idxPagesOH_21[2] | tgtPagesOH_21[2];
  assign T922[1] = idxPagesOH_21[1] | tgtPagesOH_21[1];
  assign T922[0] = idxPagesOH_21[0] | tgtPagesOH_21[0];
  assign T927[5] = pageReplEn[5] & T928[5];
  assign T927[4] = pageReplEn[4] & T928[4];
  assign T927[3] = pageReplEn[3] & T928[3];
  assign T927[2] = pageReplEn[2] & T928[2];
  assign T927[1] = pageReplEn[1] & T928[1];
  assign T927[0] = pageReplEn[0] & T928[0];
  assign T928[5] = idxPagesOH_22[5] | tgtPagesOH_22[5];
  assign T928[4] = idxPagesOH_22[4] | tgtPagesOH_22[4];
  assign T928[3] = idxPagesOH_22[3] | tgtPagesOH_22[3];
  assign T928[2] = idxPagesOH_22[2] | tgtPagesOH_22[2];
  assign T928[1] = idxPagesOH_22[1] | tgtPagesOH_22[1];
  assign T928[0] = idxPagesOH_22[0] | tgtPagesOH_22[0];
  assign T932[5] = pageReplEn[5] & T933[5];
  assign T932[4] = pageReplEn[4] & T933[4];
  assign T932[3] = pageReplEn[3] & T933[3];
  assign T932[2] = pageReplEn[2] & T933[2];
  assign T932[1] = pageReplEn[1] & T933[1];
  assign T932[0] = pageReplEn[0] & T933[0];
  assign T933[5] = idxPagesOH_23[5] | tgtPagesOH_23[5];
  assign T933[4] = idxPagesOH_23[4] | tgtPagesOH_23[4];
  assign T933[3] = idxPagesOH_23[3] | tgtPagesOH_23[3];
  assign T933[2] = idxPagesOH_23[2] | tgtPagesOH_23[2];
  assign T933[1] = idxPagesOH_23[1] | tgtPagesOH_23[1];
  assign T933[0] = idxPagesOH_23[0] | tgtPagesOH_23[0];
  assign T940[5] = pageReplEn[5] & T941[5];
  assign T940[4] = pageReplEn[4] & T941[4];
  assign T940[3] = pageReplEn[3] & T941[3];
  assign T940[2] = pageReplEn[2] & T941[2];
  assign T940[1] = pageReplEn[1] & T941[1];
  assign T940[0] = pageReplEn[0] & T941[0];
  assign T941[5] = idxPagesOH_24[5] | tgtPagesOH_24[5];
  assign T941[4] = idxPagesOH_24[4] | tgtPagesOH_24[4];
  assign T941[3] = idxPagesOH_24[3] | tgtPagesOH_24[3];
  assign T941[2] = idxPagesOH_24[2] | tgtPagesOH_24[2];
  assign T941[1] = idxPagesOH_24[1] | tgtPagesOH_24[1];
  assign T941[0] = idxPagesOH_24[0] | tgtPagesOH_24[0];
  assign T945[5] = pageReplEn[5] & T946[5];
  assign T945[4] = pageReplEn[4] & T946[4];
  assign T945[3] = pageReplEn[3] & T946[3];
  assign T945[2] = pageReplEn[2] & T946[2];
  assign T945[1] = pageReplEn[1] & T946[1];
  assign T945[0] = pageReplEn[0] & T946[0];
  assign T946[5] = idxPagesOH_25[5] | tgtPagesOH_25[5];
  assign T946[4] = idxPagesOH_25[4] | tgtPagesOH_25[4];
  assign T946[3] = idxPagesOH_25[3] | tgtPagesOH_25[3];
  assign T946[2] = idxPagesOH_25[2] | tgtPagesOH_25[2];
  assign T946[1] = idxPagesOH_25[1] | tgtPagesOH_25[1];
  assign T946[0] = idxPagesOH_25[0] | tgtPagesOH_25[0];
  assign T951[5] = pageReplEn[5] & T952[5];
  assign T951[4] = pageReplEn[4] & T952[4];
  assign T951[3] = pageReplEn[3] & T952[3];
  assign T951[2] = pageReplEn[2] & T952[2];
  assign T951[1] = pageReplEn[1] & T952[1];
  assign T951[0] = pageReplEn[0] & T952[0];
  assign T952[5] = idxPagesOH_26[5] | tgtPagesOH_26[5];
  assign T952[4] = idxPagesOH_26[4] | tgtPagesOH_26[4];
  assign T952[3] = idxPagesOH_26[3] | tgtPagesOH_26[3];
  assign T952[2] = idxPagesOH_26[2] | tgtPagesOH_26[2];
  assign T952[1] = idxPagesOH_26[1] | tgtPagesOH_26[1];
  assign T952[0] = idxPagesOH_26[0] | tgtPagesOH_26[0];
  assign T956[5] = pageReplEn[5] & T957[5];
  assign T956[4] = pageReplEn[4] & T957[4];
  assign T956[3] = pageReplEn[3] & T957[3];
  assign T956[2] = pageReplEn[2] & T957[2];
  assign T956[1] = pageReplEn[1] & T957[1];
  assign T956[0] = pageReplEn[0] & T957[0];
  assign T957[5] = idxPagesOH_27[5] | tgtPagesOH_27[5];
  assign T957[4] = idxPagesOH_27[4] | tgtPagesOH_27[4];
  assign T957[3] = idxPagesOH_27[3] | tgtPagesOH_27[3];
  assign T957[2] = idxPagesOH_27[2] | tgtPagesOH_27[2];
  assign T957[1] = idxPagesOH_27[1] | tgtPagesOH_27[1];
  assign T957[0] = idxPagesOH_27[0] | tgtPagesOH_27[0];
  assign T963[5] = pageReplEn[5] & T964[5];
  assign T963[4] = pageReplEn[4] & T964[4];
  assign T963[3] = pageReplEn[3] & T964[3];
  assign T963[2] = pageReplEn[2] & T964[2];
  assign T963[1] = pageReplEn[1] & T964[1];
  assign T963[0] = pageReplEn[0] & T964[0];
  assign T964[5] = idxPagesOH_28[5] | tgtPagesOH_28[5];
  assign T964[4] = idxPagesOH_28[4] | tgtPagesOH_28[4];
  assign T964[3] = idxPagesOH_28[3] | tgtPagesOH_28[3];
  assign T964[2] = idxPagesOH_28[2] | tgtPagesOH_28[2];
  assign T964[1] = idxPagesOH_28[1] | tgtPagesOH_28[1];
  assign T964[0] = idxPagesOH_28[0] | tgtPagesOH_28[0];
  assign T968[5] = pageReplEn[5] & T969[5];
  assign T968[4] = pageReplEn[4] & T969[4];
  assign T968[3] = pageReplEn[3] & T969[3];
  assign T968[2] = pageReplEn[2] & T969[2];
  assign T968[1] = pageReplEn[1] & T969[1];
  assign T968[0] = pageReplEn[0] & T969[0];
  assign T969[5] = idxPagesOH_29[5] | tgtPagesOH_29[5];
  assign T969[4] = idxPagesOH_29[4] | tgtPagesOH_29[4];
  assign T969[3] = idxPagesOH_29[3] | tgtPagesOH_29[3];
  assign T969[2] = idxPagesOH_29[2] | tgtPagesOH_29[2];
  assign T969[1] = idxPagesOH_29[1] | tgtPagesOH_29[1];
  assign T969[0] = idxPagesOH_29[0] | tgtPagesOH_29[0];
  assign T973[5] = pageReplEn[5] & T974[5];
  assign T973[4] = pageReplEn[4] & T974[4];
  assign T973[3] = pageReplEn[3] & T974[3];
  assign T973[2] = pageReplEn[2] & T974[2];
  assign T973[1] = pageReplEn[1] & T974[1];
  assign T973[0] = pageReplEn[0] & T974[0];
  assign T974[5] = idxPagesOH_30[5] | tgtPagesOH_30[5];
  assign T974[4] = idxPagesOH_30[4] | tgtPagesOH_30[4];
  assign T974[3] = idxPagesOH_30[3] | tgtPagesOH_30[3];
  assign T974[2] = idxPagesOH_30[2] | tgtPagesOH_30[2];
  assign T974[1] = idxPagesOH_30[1] | tgtPagesOH_30[1];
  assign T974[0] = idxPagesOH_30[0] | tgtPagesOH_30[0];
  assign T983[5] = pageReplEn[5] & T984[5];
  assign T983[4] = pageReplEn[4] & T984[4];
  assign T983[3] = pageReplEn[3] & T984[3];
  assign T983[2] = pageReplEn[2] & T984[2];
  assign T983[1] = pageReplEn[1] & T984[1];
  assign T983[0] = pageReplEn[0] & T984[0];
  assign T984[5] = idxPagesOH_31[5] | tgtPagesOH_31[5];
  assign T984[4] = idxPagesOH_31[4] | tgtPagesOH_31[4];
  assign T984[3] = idxPagesOH_31[3] | tgtPagesOH_31[3];
  assign T984[2] = idxPagesOH_31[2] | tgtPagesOH_31[2];
  assign T984[1] = idxPagesOH_31[1] | tgtPagesOH_31[1];
  assign T984[0] = idxPagesOH_31[0] | tgtPagesOH_31[0];
  assign T988[5] = pageReplEn[5] & T989[5];
  assign T988[4] = pageReplEn[4] & T989[4];
  assign T988[3] = pageReplEn[3] & T989[3];
  assign T988[2] = pageReplEn[2] & T989[2];
  assign T988[1] = pageReplEn[1] & T989[1];
  assign T988[0] = pageReplEn[0] & T989[0];
  assign T989[5] = idxPagesOH_32[5] | tgtPagesOH_32[5];
  assign T989[4] = idxPagesOH_32[4] | tgtPagesOH_32[4];
  assign T989[3] = idxPagesOH_32[3] | tgtPagesOH_32[3];
  assign T989[2] = idxPagesOH_32[2] | tgtPagesOH_32[2];
  assign T989[1] = idxPagesOH_32[1] | tgtPagesOH_32[1];
  assign T989[0] = idxPagesOH_32[0] | tgtPagesOH_32[0];
  assign T994[5] = pageReplEn[5] & T995[5];
  assign T994[4] = pageReplEn[4] & T995[4];
  assign T994[3] = pageReplEn[3] & T995[3];
  assign T994[2] = pageReplEn[2] & T995[2];
  assign T994[1] = pageReplEn[1] & T995[1];
  assign T994[0] = pageReplEn[0] & T995[0];
  assign T995[5] = idxPagesOH_33[5] | tgtPagesOH_33[5];
  assign T995[4] = idxPagesOH_33[4] | tgtPagesOH_33[4];
  assign T995[3] = idxPagesOH_33[3] | tgtPagesOH_33[3];
  assign T995[2] = idxPagesOH_33[2] | tgtPagesOH_33[2];
  assign T995[1] = idxPagesOH_33[1] | tgtPagesOH_33[1];
  assign T995[0] = idxPagesOH_33[0] | tgtPagesOH_33[0];
  assign T999[5] = pageReplEn[5] & T1000[5];
  assign T999[4] = pageReplEn[4] & T1000[4];
  assign T999[3] = pageReplEn[3] & T1000[3];
  assign T999[2] = pageReplEn[2] & T1000[2];
  assign T999[1] = pageReplEn[1] & T1000[1];
  assign T999[0] = pageReplEn[0] & T1000[0];
  assign T1000[5] = idxPagesOH_34[5] | tgtPagesOH_34[5];
  assign T1000[4] = idxPagesOH_34[4] | tgtPagesOH_34[4];
  assign T1000[3] = idxPagesOH_34[3] | tgtPagesOH_34[3];
  assign T1000[2] = idxPagesOH_34[2] | tgtPagesOH_34[2];
  assign T1000[1] = idxPagesOH_34[1] | tgtPagesOH_34[1];
  assign T1000[0] = idxPagesOH_34[0] | tgtPagesOH_34[0];
  assign T1006[5] = pageReplEn[5] & T1007[5];
  assign T1006[4] = pageReplEn[4] & T1007[4];
  assign T1006[3] = pageReplEn[3] & T1007[3];
  assign T1006[2] = pageReplEn[2] & T1007[2];
  assign T1006[1] = pageReplEn[1] & T1007[1];
  assign T1006[0] = pageReplEn[0] & T1007[0];
  assign T1007[5] = idxPagesOH_35[5] | tgtPagesOH_35[5];
  assign T1007[4] = idxPagesOH_35[4] | tgtPagesOH_35[4];
  assign T1007[3] = idxPagesOH_35[3] | tgtPagesOH_35[3];
  assign T1007[2] = idxPagesOH_35[2] | tgtPagesOH_35[2];
  assign T1007[1] = idxPagesOH_35[1] | tgtPagesOH_35[1];
  assign T1007[0] = idxPagesOH_35[0] | tgtPagesOH_35[0];
  assign T1011[5] = pageReplEn[5] & T1012[5];
  assign T1011[4] = pageReplEn[4] & T1012[4];
  assign T1011[3] = pageReplEn[3] & T1012[3];
  assign T1011[2] = pageReplEn[2] & T1012[2];
  assign T1011[1] = pageReplEn[1] & T1012[1];
  assign T1011[0] = pageReplEn[0] & T1012[0];
  assign T1012[5] = idxPagesOH_36[5] | tgtPagesOH_36[5];
  assign T1012[4] = idxPagesOH_36[4] | tgtPagesOH_36[4];
  assign T1012[3] = idxPagesOH_36[3] | tgtPagesOH_36[3];
  assign T1012[2] = idxPagesOH_36[2] | tgtPagesOH_36[2];
  assign T1012[1] = idxPagesOH_36[1] | tgtPagesOH_36[1];
  assign T1012[0] = idxPagesOH_36[0] | tgtPagesOH_36[0];
  assign T1017[5] = pageReplEn[5] & T1018[5];
  assign T1017[4] = pageReplEn[4] & T1018[4];
  assign T1017[3] = pageReplEn[3] & T1018[3];
  assign T1017[2] = pageReplEn[2] & T1018[2];
  assign T1017[1] = pageReplEn[1] & T1018[1];
  assign T1017[0] = pageReplEn[0] & T1018[0];
  assign T1018[5] = idxPagesOH_37[5] | tgtPagesOH_37[5];
  assign T1018[4] = idxPagesOH_37[4] | tgtPagesOH_37[4];
  assign T1018[3] = idxPagesOH_37[3] | tgtPagesOH_37[3];
  assign T1018[2] = idxPagesOH_37[2] | tgtPagesOH_37[2];
  assign T1018[1] = idxPagesOH_37[1] | tgtPagesOH_37[1];
  assign T1018[0] = idxPagesOH_37[0] | tgtPagesOH_37[0];
  assign T1022[5] = pageReplEn[5] & T1023[5];
  assign T1022[4] = pageReplEn[4] & T1023[4];
  assign T1022[3] = pageReplEn[3] & T1023[3];
  assign T1022[2] = pageReplEn[2] & T1023[2];
  assign T1022[1] = pageReplEn[1] & T1023[1];
  assign T1022[0] = pageReplEn[0] & T1023[0];
  assign T1023[5] = idxPagesOH_38[5] | tgtPagesOH_38[5];
  assign T1023[4] = idxPagesOH_38[4] | tgtPagesOH_38[4];
  assign T1023[3] = idxPagesOH_38[3] | tgtPagesOH_38[3];
  assign T1023[2] = idxPagesOH_38[2] | tgtPagesOH_38[2];
  assign T1023[1] = idxPagesOH_38[1] | tgtPagesOH_38[1];
  assign T1023[0] = idxPagesOH_38[0] | tgtPagesOH_38[0];
  assign T1030[5] = pageReplEn[5] & T1031[5];
  assign T1030[4] = pageReplEn[4] & T1031[4];
  assign T1030[3] = pageReplEn[3] & T1031[3];
  assign T1030[2] = pageReplEn[2] & T1031[2];
  assign T1030[1] = pageReplEn[1] & T1031[1];
  assign T1030[0] = pageReplEn[0] & T1031[0];
  assign T1031[5] = idxPagesOH_39[5] | tgtPagesOH_39[5];
  assign T1031[4] = idxPagesOH_39[4] | tgtPagesOH_39[4];
  assign T1031[3] = idxPagesOH_39[3] | tgtPagesOH_39[3];
  assign T1031[2] = idxPagesOH_39[2] | tgtPagesOH_39[2];
  assign T1031[1] = idxPagesOH_39[1] | tgtPagesOH_39[1];
  assign T1031[0] = idxPagesOH_39[0] | tgtPagesOH_39[0];
  assign T1035[5] = pageReplEn[5] & T1036[5];
  assign T1035[4] = pageReplEn[4] & T1036[4];
  assign T1035[3] = pageReplEn[3] & T1036[3];
  assign T1035[2] = pageReplEn[2] & T1036[2];
  assign T1035[1] = pageReplEn[1] & T1036[1];
  assign T1035[0] = pageReplEn[0] & T1036[0];
  assign T1036[5] = idxPagesOH_40[5] | tgtPagesOH_40[5];
  assign T1036[4] = idxPagesOH_40[4] | tgtPagesOH_40[4];
  assign T1036[3] = idxPagesOH_40[3] | tgtPagesOH_40[3];
  assign T1036[2] = idxPagesOH_40[2] | tgtPagesOH_40[2];
  assign T1036[1] = idxPagesOH_40[1] | tgtPagesOH_40[1];
  assign T1036[0] = idxPagesOH_40[0] | tgtPagesOH_40[0];
  assign T1041[5] = pageReplEn[5] & T1042[5];
  assign T1041[4] = pageReplEn[4] & T1042[4];
  assign T1041[3] = pageReplEn[3] & T1042[3];
  assign T1041[2] = pageReplEn[2] & T1042[2];
  assign T1041[1] = pageReplEn[1] & T1042[1];
  assign T1041[0] = pageReplEn[0] & T1042[0];
  assign T1042[5] = idxPagesOH_41[5] | tgtPagesOH_41[5];
  assign T1042[4] = idxPagesOH_41[4] | tgtPagesOH_41[4];
  assign T1042[3] = idxPagesOH_41[3] | tgtPagesOH_41[3];
  assign T1042[2] = idxPagesOH_41[2] | tgtPagesOH_41[2];
  assign T1042[1] = idxPagesOH_41[1] | tgtPagesOH_41[1];
  assign T1042[0] = idxPagesOH_41[0] | tgtPagesOH_41[0];
  assign T1046[5] = pageReplEn[5] & T1047[5];
  assign T1046[4] = pageReplEn[4] & T1047[4];
  assign T1046[3] = pageReplEn[3] & T1047[3];
  assign T1046[2] = pageReplEn[2] & T1047[2];
  assign T1046[1] = pageReplEn[1] & T1047[1];
  assign T1046[0] = pageReplEn[0] & T1047[0];
  assign T1047[5] = idxPagesOH_42[5] | tgtPagesOH_42[5];
  assign T1047[4] = idxPagesOH_42[4] | tgtPagesOH_42[4];
  assign T1047[3] = idxPagesOH_42[3] | tgtPagesOH_42[3];
  assign T1047[2] = idxPagesOH_42[2] | tgtPagesOH_42[2];
  assign T1047[1] = idxPagesOH_42[1] | tgtPagesOH_42[1];
  assign T1047[0] = idxPagesOH_42[0] | tgtPagesOH_42[0];
  assign T1053[5] = pageReplEn[5] & T1054[5];
  assign T1053[4] = pageReplEn[4] & T1054[4];
  assign T1053[3] = pageReplEn[3] & T1054[3];
  assign T1053[2] = pageReplEn[2] & T1054[2];
  assign T1053[1] = pageReplEn[1] & T1054[1];
  assign T1053[0] = pageReplEn[0] & T1054[0];
  assign T1054[5] = idxPagesOH_43[5] | tgtPagesOH_43[5];
  assign T1054[4] = idxPagesOH_43[4] | tgtPagesOH_43[4];
  assign T1054[3] = idxPagesOH_43[3] | tgtPagesOH_43[3];
  assign T1054[2] = idxPagesOH_43[2] | tgtPagesOH_43[2];
  assign T1054[1] = idxPagesOH_43[1] | tgtPagesOH_43[1];
  assign T1054[0] = idxPagesOH_43[0] | tgtPagesOH_43[0];
  assign T1058[5] = pageReplEn[5] & T1059[5];
  assign T1058[4] = pageReplEn[4] & T1059[4];
  assign T1058[3] = pageReplEn[3] & T1059[3];
  assign T1058[2] = pageReplEn[2] & T1059[2];
  assign T1058[1] = pageReplEn[1] & T1059[1];
  assign T1058[0] = pageReplEn[0] & T1059[0];
  assign T1059[5] = idxPagesOH_44[5] | tgtPagesOH_44[5];
  assign T1059[4] = idxPagesOH_44[4] | tgtPagesOH_44[4];
  assign T1059[3] = idxPagesOH_44[3] | tgtPagesOH_44[3];
  assign T1059[2] = idxPagesOH_44[2] | tgtPagesOH_44[2];
  assign T1059[1] = idxPagesOH_44[1] | tgtPagesOH_44[1];
  assign T1059[0] = idxPagesOH_44[0] | tgtPagesOH_44[0];
  assign T1064[5] = pageReplEn[5] & T1065[5];
  assign T1064[4] = pageReplEn[4] & T1065[4];
  assign T1064[3] = pageReplEn[3] & T1065[3];
  assign T1064[2] = pageReplEn[2] & T1065[2];
  assign T1064[1] = pageReplEn[1] & T1065[1];
  assign T1064[0] = pageReplEn[0] & T1065[0];
  assign T1065[5] = idxPagesOH_45[5] | tgtPagesOH_45[5];
  assign T1065[4] = idxPagesOH_45[4] | tgtPagesOH_45[4];
  assign T1065[3] = idxPagesOH_45[3] | tgtPagesOH_45[3];
  assign T1065[2] = idxPagesOH_45[2] | tgtPagesOH_45[2];
  assign T1065[1] = idxPagesOH_45[1] | tgtPagesOH_45[1];
  assign T1065[0] = idxPagesOH_45[0] | tgtPagesOH_45[0];
  assign T1069[5] = pageReplEn[5] & T1070[5];
  assign T1069[4] = pageReplEn[4] & T1070[4];
  assign T1069[3] = pageReplEn[3] & T1070[3];
  assign T1069[2] = pageReplEn[2] & T1070[2];
  assign T1069[1] = pageReplEn[1] & T1070[1];
  assign T1069[0] = pageReplEn[0] & T1070[0];
  assign T1070[5] = idxPagesOH_46[5] | tgtPagesOH_46[5];
  assign T1070[4] = idxPagesOH_46[4] | tgtPagesOH_46[4];
  assign T1070[3] = idxPagesOH_46[3] | tgtPagesOH_46[3];
  assign T1070[2] = idxPagesOH_46[2] | tgtPagesOH_46[2];
  assign T1070[1] = idxPagesOH_46[1] | tgtPagesOH_46[1];
  assign T1070[0] = idxPagesOH_46[0] | tgtPagesOH_46[0];
  assign T1078[5] = pageReplEn[5] & T1079[5];
  assign T1078[4] = pageReplEn[4] & T1079[4];
  assign T1078[3] = pageReplEn[3] & T1079[3];
  assign T1078[2] = pageReplEn[2] & T1079[2];
  assign T1078[1] = pageReplEn[1] & T1079[1];
  assign T1078[0] = pageReplEn[0] & T1079[0];
  assign T1079[5] = idxPagesOH_47[5] | tgtPagesOH_47[5];
  assign T1079[4] = idxPagesOH_47[4] | tgtPagesOH_47[4];
  assign T1079[3] = idxPagesOH_47[3] | tgtPagesOH_47[3];
  assign T1079[2] = idxPagesOH_47[2] | tgtPagesOH_47[2];
  assign T1079[1] = idxPagesOH_47[1] | tgtPagesOH_47[1];
  assign T1079[0] = idxPagesOH_47[0] | tgtPagesOH_47[0];
  assign T1083[5] = pageReplEn[5] & T1084[5];
  assign T1083[4] = pageReplEn[4] & T1084[4];
  assign T1083[3] = pageReplEn[3] & T1084[3];
  assign T1083[2] = pageReplEn[2] & T1084[2];
  assign T1083[1] = pageReplEn[1] & T1084[1];
  assign T1083[0] = pageReplEn[0] & T1084[0];
  assign T1084[5] = idxPagesOH_48[5] | tgtPagesOH_48[5];
  assign T1084[4] = idxPagesOH_48[4] | tgtPagesOH_48[4];
  assign T1084[3] = idxPagesOH_48[3] | tgtPagesOH_48[3];
  assign T1084[2] = idxPagesOH_48[2] | tgtPagesOH_48[2];
  assign T1084[1] = idxPagesOH_48[1] | tgtPagesOH_48[1];
  assign T1084[0] = idxPagesOH_48[0] | tgtPagesOH_48[0];
  assign T1089[5] = pageReplEn[5] & T1090[5];
  assign T1089[4] = pageReplEn[4] & T1090[4];
  assign T1089[3] = pageReplEn[3] & T1090[3];
  assign T1089[2] = pageReplEn[2] & T1090[2];
  assign T1089[1] = pageReplEn[1] & T1090[1];
  assign T1089[0] = pageReplEn[0] & T1090[0];
  assign T1090[5] = idxPagesOH_49[5] | tgtPagesOH_49[5];
  assign T1090[4] = idxPagesOH_49[4] | tgtPagesOH_49[4];
  assign T1090[3] = idxPagesOH_49[3] | tgtPagesOH_49[3];
  assign T1090[2] = idxPagesOH_49[2] | tgtPagesOH_49[2];
  assign T1090[1] = idxPagesOH_49[1] | tgtPagesOH_49[1];
  assign T1090[0] = idxPagesOH_49[0] | tgtPagesOH_49[0];
  assign T1094[5] = pageReplEn[5] & T1095[5];
  assign T1094[4] = pageReplEn[4] & T1095[4];
  assign T1094[3] = pageReplEn[3] & T1095[3];
  assign T1094[2] = pageReplEn[2] & T1095[2];
  assign T1094[1] = pageReplEn[1] & T1095[1];
  assign T1094[0] = pageReplEn[0] & T1095[0];
  assign T1095[5] = idxPagesOH_50[5] | tgtPagesOH_50[5];
  assign T1095[4] = idxPagesOH_50[4] | tgtPagesOH_50[4];
  assign T1095[3] = idxPagesOH_50[3] | tgtPagesOH_50[3];
  assign T1095[2] = idxPagesOH_50[2] | tgtPagesOH_50[2];
  assign T1095[1] = idxPagesOH_50[1] | tgtPagesOH_50[1];
  assign T1095[0] = idxPagesOH_50[0] | tgtPagesOH_50[0];
  assign T1101[5] = pageReplEn[5] & T1102[5];
  assign T1101[4] = pageReplEn[4] & T1102[4];
  assign T1101[3] = pageReplEn[3] & T1102[3];
  assign T1101[2] = pageReplEn[2] & T1102[2];
  assign T1101[1] = pageReplEn[1] & T1102[1];
  assign T1101[0] = pageReplEn[0] & T1102[0];
  assign T1102[5] = idxPagesOH_51[5] | tgtPagesOH_51[5];
  assign T1102[4] = idxPagesOH_51[4] | tgtPagesOH_51[4];
  assign T1102[3] = idxPagesOH_51[3] | tgtPagesOH_51[3];
  assign T1102[2] = idxPagesOH_51[2] | tgtPagesOH_51[2];
  assign T1102[1] = idxPagesOH_51[1] | tgtPagesOH_51[1];
  assign T1102[0] = idxPagesOH_51[0] | tgtPagesOH_51[0];
  assign T1106[5] = pageReplEn[5] & T1107[5];
  assign T1106[4] = pageReplEn[4] & T1107[4];
  assign T1106[3] = pageReplEn[3] & T1107[3];
  assign T1106[2] = pageReplEn[2] & T1107[2];
  assign T1106[1] = pageReplEn[1] & T1107[1];
  assign T1106[0] = pageReplEn[0] & T1107[0];
  assign T1107[5] = idxPagesOH_52[5] | tgtPagesOH_52[5];
  assign T1107[4] = idxPagesOH_52[4] | tgtPagesOH_52[4];
  assign T1107[3] = idxPagesOH_52[3] | tgtPagesOH_52[3];
  assign T1107[2] = idxPagesOH_52[2] | tgtPagesOH_52[2];
  assign T1107[1] = idxPagesOH_52[1] | tgtPagesOH_52[1];
  assign T1107[0] = idxPagesOH_52[0] | tgtPagesOH_52[0];
  assign T1112[5] = pageReplEn[5] & T1113[5];
  assign T1112[4] = pageReplEn[4] & T1113[4];
  assign T1112[3] = pageReplEn[3] & T1113[3];
  assign T1112[2] = pageReplEn[2] & T1113[2];
  assign T1112[1] = pageReplEn[1] & T1113[1];
  assign T1112[0] = pageReplEn[0] & T1113[0];
  assign T1113[5] = idxPagesOH_53[5] | tgtPagesOH_53[5];
  assign T1113[4] = idxPagesOH_53[4] | tgtPagesOH_53[4];
  assign T1113[3] = idxPagesOH_53[3] | tgtPagesOH_53[3];
  assign T1113[2] = idxPagesOH_53[2] | tgtPagesOH_53[2];
  assign T1113[1] = idxPagesOH_53[1] | tgtPagesOH_53[1];
  assign T1113[0] = idxPagesOH_53[0] | tgtPagesOH_53[0];
  assign T1117[5] = pageReplEn[5] & T1118[5];
  assign T1117[4] = pageReplEn[4] & T1118[4];
  assign T1117[3] = pageReplEn[3] & T1118[3];
  assign T1117[2] = pageReplEn[2] & T1118[2];
  assign T1117[1] = pageReplEn[1] & T1118[1];
  assign T1117[0] = pageReplEn[0] & T1118[0];
  assign T1118[5] = idxPagesOH_54[5] | tgtPagesOH_54[5];
  assign T1118[4] = idxPagesOH_54[4] | tgtPagesOH_54[4];
  assign T1118[3] = idxPagesOH_54[3] | tgtPagesOH_54[3];
  assign T1118[2] = idxPagesOH_54[2] | tgtPagesOH_54[2];
  assign T1118[1] = idxPagesOH_54[1] | tgtPagesOH_54[1];
  assign T1118[0] = idxPagesOH_54[0] | tgtPagesOH_54[0];
  assign T1125[5] = pageReplEn[5] & T1126[5];
  assign T1125[4] = pageReplEn[4] & T1126[4];
  assign T1125[3] = pageReplEn[3] & T1126[3];
  assign T1125[2] = pageReplEn[2] & T1126[2];
  assign T1125[1] = pageReplEn[1] & T1126[1];
  assign T1125[0] = pageReplEn[0] & T1126[0];
  assign T1126[5] = idxPagesOH_55[5] | tgtPagesOH_55[5];
  assign T1126[4] = idxPagesOH_55[4] | tgtPagesOH_55[4];
  assign T1126[3] = idxPagesOH_55[3] | tgtPagesOH_55[3];
  assign T1126[2] = idxPagesOH_55[2] | tgtPagesOH_55[2];
  assign T1126[1] = idxPagesOH_55[1] | tgtPagesOH_55[1];
  assign T1126[0] = idxPagesOH_55[0] | tgtPagesOH_55[0];
  assign T1130[5] = pageReplEn[5] & T1131[5];
  assign T1130[4] = pageReplEn[4] & T1131[4];
  assign T1130[3] = pageReplEn[3] & T1131[3];
  assign T1130[2] = pageReplEn[2] & T1131[2];
  assign T1130[1] = pageReplEn[1] & T1131[1];
  assign T1130[0] = pageReplEn[0] & T1131[0];
  assign T1131[5] = idxPagesOH_56[5] | tgtPagesOH_56[5];
  assign T1131[4] = idxPagesOH_56[4] | tgtPagesOH_56[4];
  assign T1131[3] = idxPagesOH_56[3] | tgtPagesOH_56[3];
  assign T1131[2] = idxPagesOH_56[2] | tgtPagesOH_56[2];
  assign T1131[1] = idxPagesOH_56[1] | tgtPagesOH_56[1];
  assign T1131[0] = idxPagesOH_56[0] | tgtPagesOH_56[0];
  assign T1136[5] = pageReplEn[5] & T1137[5];
  assign T1136[4] = pageReplEn[4] & T1137[4];
  assign T1136[3] = pageReplEn[3] & T1137[3];
  assign T1136[2] = pageReplEn[2] & T1137[2];
  assign T1136[1] = pageReplEn[1] & T1137[1];
  assign T1136[0] = pageReplEn[0] & T1137[0];
  assign T1137[5] = idxPagesOH_57[5] | tgtPagesOH_57[5];
  assign T1137[4] = idxPagesOH_57[4] | tgtPagesOH_57[4];
  assign T1137[3] = idxPagesOH_57[3] | tgtPagesOH_57[3];
  assign T1137[2] = idxPagesOH_57[2] | tgtPagesOH_57[2];
  assign T1137[1] = idxPagesOH_57[1] | tgtPagesOH_57[1];
  assign T1137[0] = idxPagesOH_57[0] | tgtPagesOH_57[0];
  assign T1141[5] = pageReplEn[5] & T1142[5];
  assign T1141[4] = pageReplEn[4] & T1142[4];
  assign T1141[3] = pageReplEn[3] & T1142[3];
  assign T1141[2] = pageReplEn[2] & T1142[2];
  assign T1141[1] = pageReplEn[1] & T1142[1];
  assign T1141[0] = pageReplEn[0] & T1142[0];
  assign T1142[5] = idxPagesOH_58[5] | tgtPagesOH_58[5];
  assign T1142[4] = idxPagesOH_58[4] | tgtPagesOH_58[4];
  assign T1142[3] = idxPagesOH_58[3] | tgtPagesOH_58[3];
  assign T1142[2] = idxPagesOH_58[2] | tgtPagesOH_58[2];
  assign T1142[1] = idxPagesOH_58[1] | tgtPagesOH_58[1];
  assign T1142[0] = idxPagesOH_58[0] | tgtPagesOH_58[0];
  assign T1148[5] = pageReplEn[5] & T1149[5];
  assign T1148[4] = pageReplEn[4] & T1149[4];
  assign T1148[3] = pageReplEn[3] & T1149[3];
  assign T1148[2] = pageReplEn[2] & T1149[2];
  assign T1148[1] = pageReplEn[1] & T1149[1];
  assign T1148[0] = pageReplEn[0] & T1149[0];
  assign T1149[5] = idxPagesOH_59[5] | tgtPagesOH_59[5];
  assign T1149[4] = idxPagesOH_59[4] | tgtPagesOH_59[4];
  assign T1149[3] = idxPagesOH_59[3] | tgtPagesOH_59[3];
  assign T1149[2] = idxPagesOH_59[2] | tgtPagesOH_59[2];
  assign T1149[1] = idxPagesOH_59[1] | tgtPagesOH_59[1];
  assign T1149[0] = idxPagesOH_59[0] | tgtPagesOH_59[0];
  assign T1153[5] = pageReplEn[5] & T1154[5];
  assign T1153[4] = pageReplEn[4] & T1154[4];
  assign T1153[3] = pageReplEn[3] & T1154[3];
  assign T1153[2] = pageReplEn[2] & T1154[2];
  assign T1153[1] = pageReplEn[1] & T1154[1];
  assign T1153[0] = pageReplEn[0] & T1154[0];
  assign T1154[5] = idxPagesOH_60[5] | tgtPagesOH_60[5];
  assign T1154[4] = idxPagesOH_60[4] | tgtPagesOH_60[4];
  assign T1154[3] = idxPagesOH_60[3] | tgtPagesOH_60[3];
  assign T1154[2] = idxPagesOH_60[2] | tgtPagesOH_60[2];
  assign T1154[1] = idxPagesOH_60[1] | tgtPagesOH_60[1];
  assign T1154[0] = idxPagesOH_60[0] | tgtPagesOH_60[0];
  assign T1158[5] = pageReplEn[5] & T1159[5];
  assign T1158[4] = pageReplEn[4] & T1159[4];
  assign T1158[3] = pageReplEn[3] & T1159[3];
  assign T1158[2] = pageReplEn[2] & T1159[2];
  assign T1158[1] = pageReplEn[1] & T1159[1];
  assign T1158[0] = pageReplEn[0] & T1159[0];
  assign T1159[5] = idxPagesOH_61[5] | tgtPagesOH_61[5];
  assign T1159[4] = idxPagesOH_61[4] | tgtPagesOH_61[4];
  assign T1159[3] = idxPagesOH_61[3] | tgtPagesOH_61[3];
  assign T1159[2] = idxPagesOH_61[2] | tgtPagesOH_61[2];
  assign T1159[1] = idxPagesOH_61[1] | tgtPagesOH_61[1];
  assign T1159[0] = idxPagesOH_61[0] | tgtPagesOH_61[0];
  assign T1162 = T1168 | T1163;
  assign N950 = ~hits[60];
  assign T1165 = R7 & T168[60];
  assign T1168 = T1174 | T1169;
  assign N951 = ~hits[59];
  assign T1171 = R7 & T168[59];
  assign T1174 = T1180 | T1175;
  assign N952 = ~hits[58];
  assign T1177 = R7 & T168[58];
  assign T1180 = T1186 | T1181;
  assign N953 = ~hits[57];
  assign T1183 = R7 & T168[57];
  assign T1186 = T1192 | T1187;
  assign N954 = ~hits[56];
  assign T1189 = R7 & T168[56];
  assign T1192 = T1198 | T1193;
  assign N955 = ~hits[55];
  assign T1195 = R7 & T168[55];
  assign T1198 = T1204 | T1199;
  assign N956 = ~hits[54];
  assign T1201 = R7 & T168[54];
  assign T1204 = T1210 | T1205;
  assign N957 = ~hits[53];
  assign T1207 = R7 & T168[53];
  assign T1210 = T1216 | T1211;
  assign N958 = ~hits[52];
  assign T1213 = R7 & T168[52];
  assign T1216 = T1222 | T1217;
  assign N959 = ~hits[51];
  assign T1219 = R7 & T168[51];
  assign T1222 = T1228 | T1223;
  assign N960 = ~hits[50];
  assign T1225 = R7 & T168[50];
  assign T1228 = T1234 | T1229;
  assign N961 = ~hits[49];
  assign T1231 = R7 & T168[49];
  assign T1234 = T1240 | T1235;
  assign N962 = ~hits[48];
  assign T1237 = R7 & T168[48];
  assign T1240 = T1246 | T1241;
  assign N963 = ~hits[47];
  assign T1243 = R7 & T168[47];
  assign T1246 = T1252 | T1247;
  assign N964 = ~hits[46];
  assign T1249 = R7 & T168[46];
  assign T1252 = T1258 | T1253;
  assign N965 = ~hits[45];
  assign T1255 = R7 & T168[45];
  assign T1258 = T1264 | T1259;
  assign N966 = ~hits[44];
  assign T1261 = R7 & T168[44];
  assign T1264 = T1270 | T1265;
  assign N967 = ~hits[43];
  assign T1267 = R7 & T168[43];
  assign T1270 = T1276 | T1271;
  assign N968 = ~hits[42];
  assign T1273 = R7 & T168[42];
  assign T1276 = T1282 | T1277;
  assign N969 = ~hits[41];
  assign T1279 = R7 & T168[41];
  assign T1282 = T1288 | T1283;
  assign N970 = ~hits[40];
  assign T1285 = R7 & T168[40];
  assign T1288 = T1294 | T1289;
  assign N971 = ~hits[39];
  assign T1291 = R7 & T168[39];
  assign T1294 = T1300 | T1295;
  assign N972 = ~hits[38];
  assign T1297 = R7 & T168[38];
  assign T1300 = T1306 | T1301;
  assign N973 = ~hits[37];
  assign T1303 = R7 & T168[37];
  assign T1306 = T1312 | T1307;
  assign N974 = ~hits[36];
  assign T1309 = R7 & T168[36];
  assign T1312 = T1318 | T1313;
  assign N975 = ~hits[35];
  assign T1315 = R7 & T168[35];
  assign T1318 = T1324 | T1319;
  assign N976 = ~hits[34];
  assign T1321 = R7 & T168[34];
  assign T1324 = T1330 | T1325;
  assign N977 = ~hits[33];
  assign T1327 = R7 & T168[33];
  assign T1330 = T1336 | T1331;
  assign N978 = ~hits[32];
  assign T1333 = R7 & T168[32];
  assign T1336 = T1342 | T1337;
  assign N979 = ~hits[31];
  assign T1339 = R7 & T168[31];
  assign T1342 = T1348 | T1343;
  assign N980 = ~hits[30];
  assign T1345 = R7 & T168[30];
  assign T1348 = T1354 | T1349;
  assign N981 = ~hits[29];
  assign T1351 = R7 & T168[29];
  assign T1354 = T1360 | T1355;
  assign N982 = ~hits[28];
  assign T1357 = R7 & T168[28];
  assign T1360 = T1366 | T1361;
  assign N983 = ~hits[27];
  assign T1363 = R7 & T168[27];
  assign T1366 = T1372 | T1367;
  assign N984 = ~hits[26];
  assign T1369 = R7 & T168[26];
  assign T1372 = T1378 | T1373;
  assign N985 = ~hits[25];
  assign T1375 = R7 & T168[25];
  assign T1378 = T1384 | T1379;
  assign N986 = ~hits[24];
  assign T1381 = R7 & T168[24];
  assign T1384 = T1390 | T1385;
  assign N987 = ~hits[23];
  assign T1387 = R7 & T168[23];
  assign T1390 = T1396 | T1391;
  assign N988 = ~hits[22];
  assign T1393 = R7 & T168[22];
  assign T1396 = T1402 | T1397;
  assign N989 = ~hits[21];
  assign T1399 = R7 & T168[21];
  assign T1402 = T1408 | T1403;
  assign N990 = ~hits[20];
  assign T1405 = R7 & T168[20];
  assign T1408 = T1414 | T1409;
  assign N991 = ~hits[19];
  assign T1411 = R7 & T168[19];
  assign T1414 = T1420 | T1415;
  assign N992 = ~hits[18];
  assign T1417 = R7 & T168[18];
  assign T1420 = T1426 | T1421;
  assign N993 = ~hits[17];
  assign T1423 = R7 & T168[17];
  assign T1426 = T1432 | T1427;
  assign N994 = ~hits[16];
  assign T1429 = R7 & T168[16];
  assign T1432 = T1438 | T1433;
  assign N995 = ~hits[15];
  assign T1435 = R7 & T168[15];
  assign T1438 = T1444 | T1439;
  assign N996 = ~hits[14];
  assign T1441 = R7 & T168[14];
  assign T1444 = T1450 | T1445;
  assign N997 = ~hits[13];
  assign T1447 = R7 & T168[13];
  assign T1450 = T1456 | T1451;
  assign N998 = ~hits[12];
  assign T1453 = R7 & T168[12];
  assign T1456 = T1462 | T1457;
  assign N999 = ~hits[11];
  assign T1459 = R7 & T168[11];
  assign T1462 = T1468 | T1463;
  assign N1000 = ~hits[10];
  assign T1465 = R7 & T168[10];
  assign T1468 = T1474 | T1469;
  assign N1001 = ~hits[9];
  assign T1471 = R7 & T168[9];
  assign T1474 = T1480 | T1475;
  assign N1002 = ~hits[8];
  assign T1477 = R7 & T168[8];
  assign T1480 = T1486 | T1481;
  assign N1003 = ~hits[7];
  assign T1483 = R7 & T168[7];
  assign T1486 = T1492 | T1487;
  assign N1004 = ~hits[6];
  assign T1489 = R7 & T168[6];
  assign T1492 = T1498 | T1493;
  assign N1005 = ~hits[5];
  assign T1495 = R7 & T168[5];
  assign T1498 = T1504 | T1499;
  assign N1006 = ~hits[4];
  assign T1501 = R7 & T168[4];
  assign T1504 = T1510 | T1505;
  assign N1007 = ~hits[3];
  assign T1507 = R7 & T168[3];
  assign T1510 = T1516 | T1511;
  assign N1008 = ~hits[2];
  assign T1513 = R7 & T168[2];
  assign T1516 = T1522 | T1517;
  assign N1009 = ~hits[1];
  assign T1519 = R7 & T168[1];
  assign N1010 = ~hits[0];
  assign T1524 = R7 & T168[0];
  assign T1527 = io_req_valid & io_resp_valid;
  assign T1530 = T21 & io_bht_update_bits_mispredict;
  assign io_resp_bits_entry[0] = T2458[3] | T2457[1];
  assign T2458[3] = T2460[7] | T2459[3];
  assign T2458[2] = T2460[6] | T2459[2];
  assign T2457[1] = T2460[5] | T2459[1];
  assign T2460[7] = T2462[15] | T2461[7];
  assign T2460[6] = T2462[14] | T2461[6];
  assign T2460[5] = T2462[13] | T2461[5];
  assign T2460[4] = T2462[12] | T2461[4];
  assign T2459[3] = T2462[11] | T2461[3];
  assign T2459[2] = T2462[10] | T2461[2];
  assign T2459[1] = T2462[9] | T2461[1];
  assign T2462[15] = hits[31] | T2463[15];
  assign T2462[14] = hits[30] | T2463[14];
  assign T2462[13] = T2464[29] | T2463[13];
  assign T2462[12] = T2464[28] | T2463[12];
  assign T2462[11] = T2464[27] | T2463[11];
  assign T2462[10] = T2464[26] | T2463[10];
  assign T2462[9] = T2464[25] | T2463[9];
  assign T2462[8] = T2464[24] | T2463[8];
  assign T2461[7] = T2464[23] | T2463[7];
  assign T2461[6] = T2464[22] | T2463[6];
  assign T2461[5] = T2464[21] | T2463[5];
  assign T2461[4] = T2464[20] | T2463[4];
  assign T2461[3] = T2464[19] | T2463[3];
  assign T2461[2] = T2464[18] | T2463[2];
  assign T2461[1] = T2464[17] | T2463[1];
  assign T2464[29] = hits[61] | hits[29];
  assign T2464[28] = hits[60] | hits[28];
  assign T2464[27] = hits[59] | hits[27];
  assign T2464[26] = hits[58] | hits[26];
  assign T2464[25] = hits[57] | hits[25];
  assign T2464[24] = hits[56] | hits[24];
  assign T2464[23] = hits[55] | hits[23];
  assign T2464[22] = hits[54] | hits[22];
  assign T2464[21] = hits[53] | hits[21];
  assign T2464[20] = hits[52] | hits[20];
  assign T2464[19] = hits[51] | hits[19];
  assign T2464[18] = hits[50] | hits[18];
  assign T2464[17] = hits[49] | hits[17];
  assign T2464[16] = hits[48] | hits[16];
  assign T2463[15] = hits[47] | hits[15];
  assign T2463[14] = hits[46] | hits[14];
  assign T2463[13] = hits[45] | hits[13];
  assign T2463[12] = hits[44] | hits[12];
  assign T2463[11] = hits[43] | hits[11];
  assign T2463[10] = hits[42] | hits[10];
  assign T2463[9] = hits[41] | hits[9];
  assign T2463[8] = hits[40] | hits[8];
  assign T2463[7] = hits[39] | hits[7];
  assign T2463[6] = hits[38] | hits[6];
  assign T2463[5] = hits[37] | hits[5];
  assign T2463[4] = hits[36] | hits[4];
  assign T2463[3] = hits[35] | hits[3];
  assign T2463[2] = hits[34] | hits[2];
  assign T2463[1] = hits[33] | hits[1];
  assign N1011 = ~T2406;
  assign N1012 = ~T2028;
  assign T1536[11] = T1544[11] | T1538[11];
  assign T1536[10] = T1544[10] | T1538[10];
  assign T1536[9] = T1544[9] | T1538[9];
  assign T1536[8] = T1544[8] | T1538[8];
  assign T1536[7] = T1544[7] | T1538[7];
  assign T1536[6] = T1544[6] | T1538[6];
  assign T1536[5] = T1544[5] | T1538[5];
  assign T1536[4] = T1544[4] | T1538[4];
  assign T1536[3] = T1544[3] | T1538[3];
  assign T1536[2] = T1544[2] | T1538[2];
  assign T1536[1] = T1544[1] | T1538[1];
  assign T1536[0] = T1544[0] | T1538[0];
  assign T1541 = R7 & T1542;
  assign T1544[11] = T1548[11] | T1545[11];
  assign T1544[10] = T1548[10] | T1545[10];
  assign T1544[9] = T1548[9] | T1545[9];
  assign T1544[8] = T1548[8] | T1545[8];
  assign T1544[7] = T1548[7] | T1545[7];
  assign T1544[6] = T1548[6] | T1545[6];
  assign T1544[5] = T1548[5] | T1545[5];
  assign T1544[4] = T1548[4] | T1545[4];
  assign T1544[3] = T1548[3] | T1545[3];
  assign T1544[2] = T1548[2] | T1545[2];
  assign T1544[1] = T1548[1] | T1545[1];
  assign T1544[0] = T1548[0] | T1545[0];
  assign T1548[11] = T1552[11] | T1549[11];
  assign T1548[10] = T1552[10] | T1549[10];
  assign T1548[9] = T1552[9] | T1549[9];
  assign T1548[8] = T1552[8] | T1549[8];
  assign T1548[7] = T1552[7] | T1549[7];
  assign T1548[6] = T1552[6] | T1549[6];
  assign T1548[5] = T1552[5] | T1549[5];
  assign T1548[4] = T1552[4] | T1549[4];
  assign T1548[3] = T1552[3] | T1549[3];
  assign T1548[2] = T1552[2] | T1549[2];
  assign T1548[1] = T1552[1] | T1549[1];
  assign T1548[0] = T1552[0] | T1549[0];
  assign T1552[11] = T1556[11] | T1553[11];
  assign T1552[10] = T1556[10] | T1553[10];
  assign T1552[9] = T1556[9] | T1553[9];
  assign T1552[8] = T1556[8] | T1553[8];
  assign T1552[7] = T1556[7] | T1553[7];
  assign T1552[6] = T1556[6] | T1553[6];
  assign T1552[5] = T1556[5] | T1553[5];
  assign T1552[4] = T1556[4] | T1553[4];
  assign T1552[3] = T1556[3] | T1553[3];
  assign T1552[2] = T1556[2] | T1553[2];
  assign T1552[1] = T1556[1] | T1553[1];
  assign T1552[0] = T1556[0] | T1553[0];
  assign T1556[11] = T1560[11] | T1557[11];
  assign T1556[10] = T1560[10] | T1557[10];
  assign T1556[9] = T1560[9] | T1557[9];
  assign T1556[8] = T1560[8] | T1557[8];
  assign T1556[7] = T1560[7] | T1557[7];
  assign T1556[6] = T1560[6] | T1557[6];
  assign T1556[5] = T1560[5] | T1557[5];
  assign T1556[4] = T1560[4] | T1557[4];
  assign T1556[3] = T1560[3] | T1557[3];
  assign T1556[2] = T1560[2] | T1557[2];
  assign T1556[1] = T1560[1] | T1557[1];
  assign T1556[0] = T1560[0] | T1557[0];
  assign T1560[11] = T1564[11] | T1561[11];
  assign T1560[10] = T1564[10] | T1561[10];
  assign T1560[9] = T1564[9] | T1561[9];
  assign T1560[8] = T1564[8] | T1561[8];
  assign T1560[7] = T1564[7] | T1561[7];
  assign T1560[6] = T1564[6] | T1561[6];
  assign T1560[5] = T1564[5] | T1561[5];
  assign T1560[4] = T1564[4] | T1561[4];
  assign T1560[3] = T1564[3] | T1561[3];
  assign T1560[2] = T1564[2] | T1561[2];
  assign T1560[1] = T1564[1] | T1561[1];
  assign T1560[0] = T1564[0] | T1561[0];
  assign T1564[11] = T1568[11] | T1565[11];
  assign T1564[10] = T1568[10] | T1565[10];
  assign T1564[9] = T1568[9] | T1565[9];
  assign T1564[8] = T1568[8] | T1565[8];
  assign T1564[7] = T1568[7] | T1565[7];
  assign T1564[6] = T1568[6] | T1565[6];
  assign T1564[5] = T1568[5] | T1565[5];
  assign T1564[4] = T1568[4] | T1565[4];
  assign T1564[3] = T1568[3] | T1565[3];
  assign T1564[2] = T1568[2] | T1565[2];
  assign T1564[1] = T1568[1] | T1565[1];
  assign T1564[0] = T1568[0] | T1565[0];
  assign T1568[11] = T1572[11] | T1569[11];
  assign T1568[10] = T1572[10] | T1569[10];
  assign T1568[9] = T1572[9] | T1569[9];
  assign T1568[8] = T1572[8] | T1569[8];
  assign T1568[7] = T1572[7] | T1569[7];
  assign T1568[6] = T1572[6] | T1569[6];
  assign T1568[5] = T1572[5] | T1569[5];
  assign T1568[4] = T1572[4] | T1569[4];
  assign T1568[3] = T1572[3] | T1569[3];
  assign T1568[2] = T1572[2] | T1569[2];
  assign T1568[1] = T1572[1] | T1569[1];
  assign T1568[0] = T1572[0] | T1569[0];
  assign T1572[11] = T1576[11] | T1573[11];
  assign T1572[10] = T1576[10] | T1573[10];
  assign T1572[9] = T1576[9] | T1573[9];
  assign T1572[8] = T1576[8] | T1573[8];
  assign T1572[7] = T1576[7] | T1573[7];
  assign T1572[6] = T1576[6] | T1573[6];
  assign T1572[5] = T1576[5] | T1573[5];
  assign T1572[4] = T1576[4] | T1573[4];
  assign T1572[3] = T1576[3] | T1573[3];
  assign T1572[2] = T1576[2] | T1573[2];
  assign T1572[1] = T1576[1] | T1573[1];
  assign T1572[0] = T1576[0] | T1573[0];
  assign T1576[11] = T1580[11] | T1577[11];
  assign T1576[10] = T1580[10] | T1577[10];
  assign T1576[9] = T1580[9] | T1577[9];
  assign T1576[8] = T1580[8] | T1577[8];
  assign T1576[7] = T1580[7] | T1577[7];
  assign T1576[6] = T1580[6] | T1577[6];
  assign T1576[5] = T1580[5] | T1577[5];
  assign T1576[4] = T1580[4] | T1577[4];
  assign T1576[3] = T1580[3] | T1577[3];
  assign T1576[2] = T1580[2] | T1577[2];
  assign T1576[1] = T1580[1] | T1577[1];
  assign T1576[0] = T1580[0] | T1577[0];
  assign T1580[11] = T1584[11] | T1581[11];
  assign T1580[10] = T1584[10] | T1581[10];
  assign T1580[9] = T1584[9] | T1581[9];
  assign T1580[8] = T1584[8] | T1581[8];
  assign T1580[7] = T1584[7] | T1581[7];
  assign T1580[6] = T1584[6] | T1581[6];
  assign T1580[5] = T1584[5] | T1581[5];
  assign T1580[4] = T1584[4] | T1581[4];
  assign T1580[3] = T1584[3] | T1581[3];
  assign T1580[2] = T1584[2] | T1581[2];
  assign T1580[1] = T1584[1] | T1581[1];
  assign T1580[0] = T1584[0] | T1581[0];
  assign T1584[11] = T1588[11] | T1585[11];
  assign T1584[10] = T1588[10] | T1585[10];
  assign T1584[9] = T1588[9] | T1585[9];
  assign T1584[8] = T1588[8] | T1585[8];
  assign T1584[7] = T1588[7] | T1585[7];
  assign T1584[6] = T1588[6] | T1585[6];
  assign T1584[5] = T1588[5] | T1585[5];
  assign T1584[4] = T1588[4] | T1585[4];
  assign T1584[3] = T1588[3] | T1585[3];
  assign T1584[2] = T1588[2] | T1585[2];
  assign T1584[1] = T1588[1] | T1585[1];
  assign T1584[0] = T1588[0] | T1585[0];
  assign T1588[11] = T1592[11] | T1589[11];
  assign T1588[10] = T1592[10] | T1589[10];
  assign T1588[9] = T1592[9] | T1589[9];
  assign T1588[8] = T1592[8] | T1589[8];
  assign T1588[7] = T1592[7] | T1589[7];
  assign T1588[6] = T1592[6] | T1589[6];
  assign T1588[5] = T1592[5] | T1589[5];
  assign T1588[4] = T1592[4] | T1589[4];
  assign T1588[3] = T1592[3] | T1589[3];
  assign T1588[2] = T1592[2] | T1589[2];
  assign T1588[1] = T1592[1] | T1589[1];
  assign T1588[0] = T1592[0] | T1589[0];
  assign T1592[11] = T1596[11] | T1593[11];
  assign T1592[10] = T1596[10] | T1593[10];
  assign T1592[9] = T1596[9] | T1593[9];
  assign T1592[8] = T1596[8] | T1593[8];
  assign T1592[7] = T1596[7] | T1593[7];
  assign T1592[6] = T1596[6] | T1593[6];
  assign T1592[5] = T1596[5] | T1593[5];
  assign T1592[4] = T1596[4] | T1593[4];
  assign T1592[3] = T1596[3] | T1593[3];
  assign T1592[2] = T1596[2] | T1593[2];
  assign T1592[1] = T1596[1] | T1593[1];
  assign T1592[0] = T1596[0] | T1593[0];
  assign T1596[11] = T1600[11] | T1597[11];
  assign T1596[10] = T1600[10] | T1597[10];
  assign T1596[9] = T1600[9] | T1597[9];
  assign T1596[8] = T1600[8] | T1597[8];
  assign T1596[7] = T1600[7] | T1597[7];
  assign T1596[6] = T1600[6] | T1597[6];
  assign T1596[5] = T1600[5] | T1597[5];
  assign T1596[4] = T1600[4] | T1597[4];
  assign T1596[3] = T1600[3] | T1597[3];
  assign T1596[2] = T1600[2] | T1597[2];
  assign T1596[1] = T1600[1] | T1597[1];
  assign T1596[0] = T1600[0] | T1597[0];
  assign T1600[11] = T1604[11] | T1601[11];
  assign T1600[10] = T1604[10] | T1601[10];
  assign T1600[9] = T1604[9] | T1601[9];
  assign T1600[8] = T1604[8] | T1601[8];
  assign T1600[7] = T1604[7] | T1601[7];
  assign T1600[6] = T1604[6] | T1601[6];
  assign T1600[5] = T1604[5] | T1601[5];
  assign T1600[4] = T1604[4] | T1601[4];
  assign T1600[3] = T1604[3] | T1601[3];
  assign T1600[2] = T1604[2] | T1601[2];
  assign T1600[1] = T1604[1] | T1601[1];
  assign T1600[0] = T1604[0] | T1601[0];
  assign T1604[11] = T1608[11] | T1605[11];
  assign T1604[10] = T1608[10] | T1605[10];
  assign T1604[9] = T1608[9] | T1605[9];
  assign T1604[8] = T1608[8] | T1605[8];
  assign T1604[7] = T1608[7] | T1605[7];
  assign T1604[6] = T1608[6] | T1605[6];
  assign T1604[5] = T1608[5] | T1605[5];
  assign T1604[4] = T1608[4] | T1605[4];
  assign T1604[3] = T1608[3] | T1605[3];
  assign T1604[2] = T1608[2] | T1605[2];
  assign T1604[1] = T1608[1] | T1605[1];
  assign T1604[0] = T1608[0] | T1605[0];
  assign T1608[11] = T1612[11] | T1609[11];
  assign T1608[10] = T1612[10] | T1609[10];
  assign T1608[9] = T1612[9] | T1609[9];
  assign T1608[8] = T1612[8] | T1609[8];
  assign T1608[7] = T1612[7] | T1609[7];
  assign T1608[6] = T1612[6] | T1609[6];
  assign T1608[5] = T1612[5] | T1609[5];
  assign T1608[4] = T1612[4] | T1609[4];
  assign T1608[3] = T1612[3] | T1609[3];
  assign T1608[2] = T1612[2] | T1609[2];
  assign T1608[1] = T1612[1] | T1609[1];
  assign T1608[0] = T1612[0] | T1609[0];
  assign T1612[11] = T1616[11] | T1613[11];
  assign T1612[10] = T1616[10] | T1613[10];
  assign T1612[9] = T1616[9] | T1613[9];
  assign T1612[8] = T1616[8] | T1613[8];
  assign T1612[7] = T1616[7] | T1613[7];
  assign T1612[6] = T1616[6] | T1613[6];
  assign T1612[5] = T1616[5] | T1613[5];
  assign T1612[4] = T1616[4] | T1613[4];
  assign T1612[3] = T1616[3] | T1613[3];
  assign T1612[2] = T1616[2] | T1613[2];
  assign T1612[1] = T1616[1] | T1613[1];
  assign T1612[0] = T1616[0] | T1613[0];
  assign T1616[11] = T1620[11] | T1617[11];
  assign T1616[10] = T1620[10] | T1617[10];
  assign T1616[9] = T1620[9] | T1617[9];
  assign T1616[8] = T1620[8] | T1617[8];
  assign T1616[7] = T1620[7] | T1617[7];
  assign T1616[6] = T1620[6] | T1617[6];
  assign T1616[5] = T1620[5] | T1617[5];
  assign T1616[4] = T1620[4] | T1617[4];
  assign T1616[3] = T1620[3] | T1617[3];
  assign T1616[2] = T1620[2] | T1617[2];
  assign T1616[1] = T1620[1] | T1617[1];
  assign T1616[0] = T1620[0] | T1617[0];
  assign T1620[11] = T1624[11] | T1621[11];
  assign T1620[10] = T1624[10] | T1621[10];
  assign T1620[9] = T1624[9] | T1621[9];
  assign T1620[8] = T1624[8] | T1621[8];
  assign T1620[7] = T1624[7] | T1621[7];
  assign T1620[6] = T1624[6] | T1621[6];
  assign T1620[5] = T1624[5] | T1621[5];
  assign T1620[4] = T1624[4] | T1621[4];
  assign T1620[3] = T1624[3] | T1621[3];
  assign T1620[2] = T1624[2] | T1621[2];
  assign T1620[1] = T1624[1] | T1621[1];
  assign T1620[0] = T1624[0] | T1621[0];
  assign T1624[11] = T1628[11] | T1625[11];
  assign T1624[10] = T1628[10] | T1625[10];
  assign T1624[9] = T1628[9] | T1625[9];
  assign T1624[8] = T1628[8] | T1625[8];
  assign T1624[7] = T1628[7] | T1625[7];
  assign T1624[6] = T1628[6] | T1625[6];
  assign T1624[5] = T1628[5] | T1625[5];
  assign T1624[4] = T1628[4] | T1625[4];
  assign T1624[3] = T1628[3] | T1625[3];
  assign T1624[2] = T1628[2] | T1625[2];
  assign T1624[1] = T1628[1] | T1625[1];
  assign T1624[0] = T1628[0] | T1625[0];
  assign T1628[11] = T1632[11] | T1629[11];
  assign T1628[10] = T1632[10] | T1629[10];
  assign T1628[9] = T1632[9] | T1629[9];
  assign T1628[8] = T1632[8] | T1629[8];
  assign T1628[7] = T1632[7] | T1629[7];
  assign T1628[6] = T1632[6] | T1629[6];
  assign T1628[5] = T1632[5] | T1629[5];
  assign T1628[4] = T1632[4] | T1629[4];
  assign T1628[3] = T1632[3] | T1629[3];
  assign T1628[2] = T1632[2] | T1629[2];
  assign T1628[1] = T1632[1] | T1629[1];
  assign T1628[0] = T1632[0] | T1629[0];
  assign T1632[11] = T1636[11] | T1633[11];
  assign T1632[10] = T1636[10] | T1633[10];
  assign T1632[9] = T1636[9] | T1633[9];
  assign T1632[8] = T1636[8] | T1633[8];
  assign T1632[7] = T1636[7] | T1633[7];
  assign T1632[6] = T1636[6] | T1633[6];
  assign T1632[5] = T1636[5] | T1633[5];
  assign T1632[4] = T1636[4] | T1633[4];
  assign T1632[3] = T1636[3] | T1633[3];
  assign T1632[2] = T1636[2] | T1633[2];
  assign T1632[1] = T1636[1] | T1633[1];
  assign T1632[0] = T1636[0] | T1633[0];
  assign T1636[11] = T1640[11] | T1637[11];
  assign T1636[10] = T1640[10] | T1637[10];
  assign T1636[9] = T1640[9] | T1637[9];
  assign T1636[8] = T1640[8] | T1637[8];
  assign T1636[7] = T1640[7] | T1637[7];
  assign T1636[6] = T1640[6] | T1637[6];
  assign T1636[5] = T1640[5] | T1637[5];
  assign T1636[4] = T1640[4] | T1637[4];
  assign T1636[3] = T1640[3] | T1637[3];
  assign T1636[2] = T1640[2] | T1637[2];
  assign T1636[1] = T1640[1] | T1637[1];
  assign T1636[0] = T1640[0] | T1637[0];
  assign T1640[11] = T1644[11] | T1641[11];
  assign T1640[10] = T1644[10] | T1641[10];
  assign T1640[9] = T1644[9] | T1641[9];
  assign T1640[8] = T1644[8] | T1641[8];
  assign T1640[7] = T1644[7] | T1641[7];
  assign T1640[6] = T1644[6] | T1641[6];
  assign T1640[5] = T1644[5] | T1641[5];
  assign T1640[4] = T1644[4] | T1641[4];
  assign T1640[3] = T1644[3] | T1641[3];
  assign T1640[2] = T1644[2] | T1641[2];
  assign T1640[1] = T1644[1] | T1641[1];
  assign T1640[0] = T1644[0] | T1641[0];
  assign T1644[11] = T1648[11] | T1645[11];
  assign T1644[10] = T1648[10] | T1645[10];
  assign T1644[9] = T1648[9] | T1645[9];
  assign T1644[8] = T1648[8] | T1645[8];
  assign T1644[7] = T1648[7] | T1645[7];
  assign T1644[6] = T1648[6] | T1645[6];
  assign T1644[5] = T1648[5] | T1645[5];
  assign T1644[4] = T1648[4] | T1645[4];
  assign T1644[3] = T1648[3] | T1645[3];
  assign T1644[2] = T1648[2] | T1645[2];
  assign T1644[1] = T1648[1] | T1645[1];
  assign T1644[0] = T1648[0] | T1645[0];
  assign T1648[11] = T1652[11] | T1649[11];
  assign T1648[10] = T1652[10] | T1649[10];
  assign T1648[9] = T1652[9] | T1649[9];
  assign T1648[8] = T1652[8] | T1649[8];
  assign T1648[7] = T1652[7] | T1649[7];
  assign T1648[6] = T1652[6] | T1649[6];
  assign T1648[5] = T1652[5] | T1649[5];
  assign T1648[4] = T1652[4] | T1649[4];
  assign T1648[3] = T1652[3] | T1649[3];
  assign T1648[2] = T1652[2] | T1649[2];
  assign T1648[1] = T1652[1] | T1649[1];
  assign T1648[0] = T1652[0] | T1649[0];
  assign T1652[11] = T1656[11] | T1653[11];
  assign T1652[10] = T1656[10] | T1653[10];
  assign T1652[9] = T1656[9] | T1653[9];
  assign T1652[8] = T1656[8] | T1653[8];
  assign T1652[7] = T1656[7] | T1653[7];
  assign T1652[6] = T1656[6] | T1653[6];
  assign T1652[5] = T1656[5] | T1653[5];
  assign T1652[4] = T1656[4] | T1653[4];
  assign T1652[3] = T1656[3] | T1653[3];
  assign T1652[2] = T1656[2] | T1653[2];
  assign T1652[1] = T1656[1] | T1653[1];
  assign T1652[0] = T1656[0] | T1653[0];
  assign T1656[11] = T1660[11] | T1657[11];
  assign T1656[10] = T1660[10] | T1657[10];
  assign T1656[9] = T1660[9] | T1657[9];
  assign T1656[8] = T1660[8] | T1657[8];
  assign T1656[7] = T1660[7] | T1657[7];
  assign T1656[6] = T1660[6] | T1657[6];
  assign T1656[5] = T1660[5] | T1657[5];
  assign T1656[4] = T1660[4] | T1657[4];
  assign T1656[3] = T1660[3] | T1657[3];
  assign T1656[2] = T1660[2] | T1657[2];
  assign T1656[1] = T1660[1] | T1657[1];
  assign T1656[0] = T1660[0] | T1657[0];
  assign T1660[11] = T1664[11] | T1661[11];
  assign T1660[10] = T1664[10] | T1661[10];
  assign T1660[9] = T1664[9] | T1661[9];
  assign T1660[8] = T1664[8] | T1661[8];
  assign T1660[7] = T1664[7] | T1661[7];
  assign T1660[6] = T1664[6] | T1661[6];
  assign T1660[5] = T1664[5] | T1661[5];
  assign T1660[4] = T1664[4] | T1661[4];
  assign T1660[3] = T1664[3] | T1661[3];
  assign T1660[2] = T1664[2] | T1661[2];
  assign T1660[1] = T1664[1] | T1661[1];
  assign T1660[0] = T1664[0] | T1661[0];
  assign T1664[11] = T1668[11] | T1665[11];
  assign T1664[10] = T1668[10] | T1665[10];
  assign T1664[9] = T1668[9] | T1665[9];
  assign T1664[8] = T1668[8] | T1665[8];
  assign T1664[7] = T1668[7] | T1665[7];
  assign T1664[6] = T1668[6] | T1665[6];
  assign T1664[5] = T1668[5] | T1665[5];
  assign T1664[4] = T1668[4] | T1665[4];
  assign T1664[3] = T1668[3] | T1665[3];
  assign T1664[2] = T1668[2] | T1665[2];
  assign T1664[1] = T1668[1] | T1665[1];
  assign T1664[0] = T1668[0] | T1665[0];
  assign T1668[11] = T1672[11] | T1669[11];
  assign T1668[10] = T1672[10] | T1669[10];
  assign T1668[9] = T1672[9] | T1669[9];
  assign T1668[8] = T1672[8] | T1669[8];
  assign T1668[7] = T1672[7] | T1669[7];
  assign T1668[6] = T1672[6] | T1669[6];
  assign T1668[5] = T1672[5] | T1669[5];
  assign T1668[4] = T1672[4] | T1669[4];
  assign T1668[3] = T1672[3] | T1669[3];
  assign T1668[2] = T1672[2] | T1669[2];
  assign T1668[1] = T1672[1] | T1669[1];
  assign T1668[0] = T1672[0] | T1669[0];
  assign T1672[11] = T1676[11] | T1673[11];
  assign T1672[10] = T1676[10] | T1673[10];
  assign T1672[9] = T1676[9] | T1673[9];
  assign T1672[8] = T1676[8] | T1673[8];
  assign T1672[7] = T1676[7] | T1673[7];
  assign T1672[6] = T1676[6] | T1673[6];
  assign T1672[5] = T1676[5] | T1673[5];
  assign T1672[4] = T1676[4] | T1673[4];
  assign T1672[3] = T1676[3] | T1673[3];
  assign T1672[2] = T1676[2] | T1673[2];
  assign T1672[1] = T1676[1] | T1673[1];
  assign T1672[0] = T1676[0] | T1673[0];
  assign T1676[11] = T1680[11] | T1677[11];
  assign T1676[10] = T1680[10] | T1677[10];
  assign T1676[9] = T1680[9] | T1677[9];
  assign T1676[8] = T1680[8] | T1677[8];
  assign T1676[7] = T1680[7] | T1677[7];
  assign T1676[6] = T1680[6] | T1677[6];
  assign T1676[5] = T1680[5] | T1677[5];
  assign T1676[4] = T1680[4] | T1677[4];
  assign T1676[3] = T1680[3] | T1677[3];
  assign T1676[2] = T1680[2] | T1677[2];
  assign T1676[1] = T1680[1] | T1677[1];
  assign T1676[0] = T1680[0] | T1677[0];
  assign T1680[11] = T1684[11] | T1681[11];
  assign T1680[10] = T1684[10] | T1681[10];
  assign T1680[9] = T1684[9] | T1681[9];
  assign T1680[8] = T1684[8] | T1681[8];
  assign T1680[7] = T1684[7] | T1681[7];
  assign T1680[6] = T1684[6] | T1681[6];
  assign T1680[5] = T1684[5] | T1681[5];
  assign T1680[4] = T1684[4] | T1681[4];
  assign T1680[3] = T1684[3] | T1681[3];
  assign T1680[2] = T1684[2] | T1681[2];
  assign T1680[1] = T1684[1] | T1681[1];
  assign T1680[0] = T1684[0] | T1681[0];
  assign T1684[11] = T1688[11] | T1685[11];
  assign T1684[10] = T1688[10] | T1685[10];
  assign T1684[9] = T1688[9] | T1685[9];
  assign T1684[8] = T1688[8] | T1685[8];
  assign T1684[7] = T1688[7] | T1685[7];
  assign T1684[6] = T1688[6] | T1685[6];
  assign T1684[5] = T1688[5] | T1685[5];
  assign T1684[4] = T1688[4] | T1685[4];
  assign T1684[3] = T1688[3] | T1685[3];
  assign T1684[2] = T1688[2] | T1685[2];
  assign T1684[1] = T1688[1] | T1685[1];
  assign T1684[0] = T1688[0] | T1685[0];
  assign T1688[11] = T1692[11] | T1689[11];
  assign T1688[10] = T1692[10] | T1689[10];
  assign T1688[9] = T1692[9] | T1689[9];
  assign T1688[8] = T1692[8] | T1689[8];
  assign T1688[7] = T1692[7] | T1689[7];
  assign T1688[6] = T1692[6] | T1689[6];
  assign T1688[5] = T1692[5] | T1689[5];
  assign T1688[4] = T1692[4] | T1689[4];
  assign T1688[3] = T1692[3] | T1689[3];
  assign T1688[2] = T1692[2] | T1689[2];
  assign T1688[1] = T1692[1] | T1689[1];
  assign T1688[0] = T1692[0] | T1689[0];
  assign T1692[11] = T1696[11] | T1693[11];
  assign T1692[10] = T1696[10] | T1693[10];
  assign T1692[9] = T1696[9] | T1693[9];
  assign T1692[8] = T1696[8] | T1693[8];
  assign T1692[7] = T1696[7] | T1693[7];
  assign T1692[6] = T1696[6] | T1693[6];
  assign T1692[5] = T1696[5] | T1693[5];
  assign T1692[4] = T1696[4] | T1693[4];
  assign T1692[3] = T1696[3] | T1693[3];
  assign T1692[2] = T1696[2] | T1693[2];
  assign T1692[1] = T1696[1] | T1693[1];
  assign T1692[0] = T1696[0] | T1693[0];
  assign T1696[11] = T1700[11] | T1697[11];
  assign T1696[10] = T1700[10] | T1697[10];
  assign T1696[9] = T1700[9] | T1697[9];
  assign T1696[8] = T1700[8] | T1697[8];
  assign T1696[7] = T1700[7] | T1697[7];
  assign T1696[6] = T1700[6] | T1697[6];
  assign T1696[5] = T1700[5] | T1697[5];
  assign T1696[4] = T1700[4] | T1697[4];
  assign T1696[3] = T1700[3] | T1697[3];
  assign T1696[2] = T1700[2] | T1697[2];
  assign T1696[1] = T1700[1] | T1697[1];
  assign T1696[0] = T1700[0] | T1697[0];
  assign T1700[11] = T1704[11] | T1701[11];
  assign T1700[10] = T1704[10] | T1701[10];
  assign T1700[9] = T1704[9] | T1701[9];
  assign T1700[8] = T1704[8] | T1701[8];
  assign T1700[7] = T1704[7] | T1701[7];
  assign T1700[6] = T1704[6] | T1701[6];
  assign T1700[5] = T1704[5] | T1701[5];
  assign T1700[4] = T1704[4] | T1701[4];
  assign T1700[3] = T1704[3] | T1701[3];
  assign T1700[2] = T1704[2] | T1701[2];
  assign T1700[1] = T1704[1] | T1701[1];
  assign T1700[0] = T1704[0] | T1701[0];
  assign T1704[11] = T1708[11] | T1705[11];
  assign T1704[10] = T1708[10] | T1705[10];
  assign T1704[9] = T1708[9] | T1705[9];
  assign T1704[8] = T1708[8] | T1705[8];
  assign T1704[7] = T1708[7] | T1705[7];
  assign T1704[6] = T1708[6] | T1705[6];
  assign T1704[5] = T1708[5] | T1705[5];
  assign T1704[4] = T1708[4] | T1705[4];
  assign T1704[3] = T1708[3] | T1705[3];
  assign T1704[2] = T1708[2] | T1705[2];
  assign T1704[1] = T1708[1] | T1705[1];
  assign T1704[0] = T1708[0] | T1705[0];
  assign T1708[11] = T1712[11] | T1709[11];
  assign T1708[10] = T1712[10] | T1709[10];
  assign T1708[9] = T1712[9] | T1709[9];
  assign T1708[8] = T1712[8] | T1709[8];
  assign T1708[7] = T1712[7] | T1709[7];
  assign T1708[6] = T1712[6] | T1709[6];
  assign T1708[5] = T1712[5] | T1709[5];
  assign T1708[4] = T1712[4] | T1709[4];
  assign T1708[3] = T1712[3] | T1709[3];
  assign T1708[2] = T1712[2] | T1709[2];
  assign T1708[1] = T1712[1] | T1709[1];
  assign T1708[0] = T1712[0] | T1709[0];
  assign T1712[11] = T1716[11] | T1713[11];
  assign T1712[10] = T1716[10] | T1713[10];
  assign T1712[9] = T1716[9] | T1713[9];
  assign T1712[8] = T1716[8] | T1713[8];
  assign T1712[7] = T1716[7] | T1713[7];
  assign T1712[6] = T1716[6] | T1713[6];
  assign T1712[5] = T1716[5] | T1713[5];
  assign T1712[4] = T1716[4] | T1713[4];
  assign T1712[3] = T1716[3] | T1713[3];
  assign T1712[2] = T1716[2] | T1713[2];
  assign T1712[1] = T1716[1] | T1713[1];
  assign T1712[0] = T1716[0] | T1713[0];
  assign T1716[11] = T1720[11] | T1717[11];
  assign T1716[10] = T1720[10] | T1717[10];
  assign T1716[9] = T1720[9] | T1717[9];
  assign T1716[8] = T1720[8] | T1717[8];
  assign T1716[7] = T1720[7] | T1717[7];
  assign T1716[6] = T1720[6] | T1717[6];
  assign T1716[5] = T1720[5] | T1717[5];
  assign T1716[4] = T1720[4] | T1717[4];
  assign T1716[3] = T1720[3] | T1717[3];
  assign T1716[2] = T1720[2] | T1717[2];
  assign T1716[1] = T1720[1] | T1717[1];
  assign T1716[0] = T1720[0] | T1717[0];
  assign T1720[11] = T1724[11] | T1721[11];
  assign T1720[10] = T1724[10] | T1721[10];
  assign T1720[9] = T1724[9] | T1721[9];
  assign T1720[8] = T1724[8] | T1721[8];
  assign T1720[7] = T1724[7] | T1721[7];
  assign T1720[6] = T1724[6] | T1721[6];
  assign T1720[5] = T1724[5] | T1721[5];
  assign T1720[4] = T1724[4] | T1721[4];
  assign T1720[3] = T1724[3] | T1721[3];
  assign T1720[2] = T1724[2] | T1721[2];
  assign T1720[1] = T1724[1] | T1721[1];
  assign T1720[0] = T1724[0] | T1721[0];
  assign T1724[11] = T1728[11] | T1725[11];
  assign T1724[10] = T1728[10] | T1725[10];
  assign T1724[9] = T1728[9] | T1725[9];
  assign T1724[8] = T1728[8] | T1725[8];
  assign T1724[7] = T1728[7] | T1725[7];
  assign T1724[6] = T1728[6] | T1725[6];
  assign T1724[5] = T1728[5] | T1725[5];
  assign T1724[4] = T1728[4] | T1725[4];
  assign T1724[3] = T1728[3] | T1725[3];
  assign T1724[2] = T1728[2] | T1725[2];
  assign T1724[1] = T1728[1] | T1725[1];
  assign T1724[0] = T1728[0] | T1725[0];
  assign T1728[11] = T1732[11] | T1729[11];
  assign T1728[10] = T1732[10] | T1729[10];
  assign T1728[9] = T1732[9] | T1729[9];
  assign T1728[8] = T1732[8] | T1729[8];
  assign T1728[7] = T1732[7] | T1729[7];
  assign T1728[6] = T1732[6] | T1729[6];
  assign T1728[5] = T1732[5] | T1729[5];
  assign T1728[4] = T1732[4] | T1729[4];
  assign T1728[3] = T1732[3] | T1729[3];
  assign T1728[2] = T1732[2] | T1729[2];
  assign T1728[1] = T1732[1] | T1729[1];
  assign T1728[0] = T1732[0] | T1729[0];
  assign T1732[11] = T1736[11] | T1733[11];
  assign T1732[10] = T1736[10] | T1733[10];
  assign T1732[9] = T1736[9] | T1733[9];
  assign T1732[8] = T1736[8] | T1733[8];
  assign T1732[7] = T1736[7] | T1733[7];
  assign T1732[6] = T1736[6] | T1733[6];
  assign T1732[5] = T1736[5] | T1733[5];
  assign T1732[4] = T1736[4] | T1733[4];
  assign T1732[3] = T1736[3] | T1733[3];
  assign T1732[2] = T1736[2] | T1733[2];
  assign T1732[1] = T1736[1] | T1733[1];
  assign T1732[0] = T1736[0] | T1733[0];
  assign T1736[11] = T1740[11] | T1737[11];
  assign T1736[10] = T1740[10] | T1737[10];
  assign T1736[9] = T1740[9] | T1737[9];
  assign T1736[8] = T1740[8] | T1737[8];
  assign T1736[7] = T1740[7] | T1737[7];
  assign T1736[6] = T1740[6] | T1737[6];
  assign T1736[5] = T1740[5] | T1737[5];
  assign T1736[4] = T1740[4] | T1737[4];
  assign T1736[3] = T1740[3] | T1737[3];
  assign T1736[2] = T1740[2] | T1737[2];
  assign T1736[1] = T1740[1] | T1737[1];
  assign T1736[0] = T1740[0] | T1737[0];
  assign T1740[11] = T1744[11] | T1741[11];
  assign T1740[10] = T1744[10] | T1741[10];
  assign T1740[9] = T1744[9] | T1741[9];
  assign T1740[8] = T1744[8] | T1741[8];
  assign T1740[7] = T1744[7] | T1741[7];
  assign T1740[6] = T1744[6] | T1741[6];
  assign T1740[5] = T1744[5] | T1741[5];
  assign T1740[4] = T1744[4] | T1741[4];
  assign T1740[3] = T1744[3] | T1741[3];
  assign T1740[2] = T1744[2] | T1741[2];
  assign T1740[1] = T1744[1] | T1741[1];
  assign T1740[0] = T1744[0] | T1741[0];
  assign T1744[11] = T1748[11] | T1745[11];
  assign T1744[10] = T1748[10] | T1745[10];
  assign T1744[9] = T1748[9] | T1745[9];
  assign T1744[8] = T1748[8] | T1745[8];
  assign T1744[7] = T1748[7] | T1745[7];
  assign T1744[6] = T1748[6] | T1745[6];
  assign T1744[5] = T1748[5] | T1745[5];
  assign T1744[4] = T1748[4] | T1745[4];
  assign T1744[3] = T1748[3] | T1745[3];
  assign T1744[2] = T1748[2] | T1745[2];
  assign T1744[1] = T1748[1] | T1745[1];
  assign T1744[0] = T1748[0] | T1745[0];
  assign T1748[11] = T1752[11] | T1749[11];
  assign T1748[10] = T1752[10] | T1749[10];
  assign T1748[9] = T1752[9] | T1749[9];
  assign T1748[8] = T1752[8] | T1749[8];
  assign T1748[7] = T1752[7] | T1749[7];
  assign T1748[6] = T1752[6] | T1749[6];
  assign T1748[5] = T1752[5] | T1749[5];
  assign T1748[4] = T1752[4] | T1749[4];
  assign T1748[3] = T1752[3] | T1749[3];
  assign T1748[2] = T1752[2] | T1749[2];
  assign T1748[1] = T1752[1] | T1749[1];
  assign T1748[0] = T1752[0] | T1749[0];
  assign T1752[11] = T1756[11] | T1753[11];
  assign T1752[10] = T1756[10] | T1753[10];
  assign T1752[9] = T1756[9] | T1753[9];
  assign T1752[8] = T1756[8] | T1753[8];
  assign T1752[7] = T1756[7] | T1753[7];
  assign T1752[6] = T1756[6] | T1753[6];
  assign T1752[5] = T1756[5] | T1753[5];
  assign T1752[4] = T1756[4] | T1753[4];
  assign T1752[3] = T1756[3] | T1753[3];
  assign T1752[2] = T1756[2] | T1753[2];
  assign T1752[1] = T1756[1] | T1753[1];
  assign T1752[0] = T1756[0] | T1753[0];
  assign T1756[11] = T1760[11] | T1757[11];
  assign T1756[10] = T1760[10] | T1757[10];
  assign T1756[9] = T1760[9] | T1757[9];
  assign T1756[8] = T1760[8] | T1757[8];
  assign T1756[7] = T1760[7] | T1757[7];
  assign T1756[6] = T1760[6] | T1757[6];
  assign T1756[5] = T1760[5] | T1757[5];
  assign T1756[4] = T1760[4] | T1757[4];
  assign T1756[3] = T1760[3] | T1757[3];
  assign T1756[2] = T1760[2] | T1757[2];
  assign T1756[1] = T1760[1] | T1757[1];
  assign T1756[0] = T1760[0] | T1757[0];
  assign T1760[11] = T1764[11] | T1761[11];
  assign T1760[10] = T1764[10] | T1761[10];
  assign T1760[9] = T1764[9] | T1761[9];
  assign T1760[8] = T1764[8] | T1761[8];
  assign T1760[7] = T1764[7] | T1761[7];
  assign T1760[6] = T1764[6] | T1761[6];
  assign T1760[5] = T1764[5] | T1761[5];
  assign T1760[4] = T1764[4] | T1761[4];
  assign T1760[3] = T1764[3] | T1761[3];
  assign T1760[2] = T1764[2] | T1761[2];
  assign T1760[1] = T1764[1] | T1761[1];
  assign T1760[0] = T1764[0] | T1761[0];
  assign T1764[11] = T1768[11] | T1765[11];
  assign T1764[10] = T1768[10] | T1765[10];
  assign T1764[9] = T1768[9] | T1765[9];
  assign T1764[8] = T1768[8] | T1765[8];
  assign T1764[7] = T1768[7] | T1765[7];
  assign T1764[6] = T1768[6] | T1765[6];
  assign T1764[5] = T1768[5] | T1765[5];
  assign T1764[4] = T1768[4] | T1765[4];
  assign T1764[3] = T1768[3] | T1765[3];
  assign T1764[2] = T1768[2] | T1765[2];
  assign T1764[1] = T1768[1] | T1765[1];
  assign T1764[0] = T1768[0] | T1765[0];
  assign T1768[11] = T1772[11] | T1769[11];
  assign T1768[10] = T1772[10] | T1769[10];
  assign T1768[9] = T1772[9] | T1769[9];
  assign T1768[8] = T1772[8] | T1769[8];
  assign T1768[7] = T1772[7] | T1769[7];
  assign T1768[6] = T1772[6] | T1769[6];
  assign T1768[5] = T1772[5] | T1769[5];
  assign T1768[4] = T1772[4] | T1769[4];
  assign T1768[3] = T1772[3] | T1769[3];
  assign T1768[2] = T1772[2] | T1769[2];
  assign T1768[1] = T1772[1] | T1769[1];
  assign T1768[0] = T1772[0] | T1769[0];
  assign T1772[11] = T1776[11] | T1773[11];
  assign T1772[10] = T1776[10] | T1773[10];
  assign T1772[9] = T1776[9] | T1773[9];
  assign T1772[8] = T1776[8] | T1773[8];
  assign T1772[7] = T1776[7] | T1773[7];
  assign T1772[6] = T1776[6] | T1773[6];
  assign T1772[5] = T1776[5] | T1773[5];
  assign T1772[4] = T1776[4] | T1773[4];
  assign T1772[3] = T1776[3] | T1773[3];
  assign T1772[2] = T1776[2] | T1773[2];
  assign T1772[1] = T1776[1] | T1773[1];
  assign T1772[0] = T1776[0] | T1773[0];
  assign T1776[11] = T1780[11] | T1777[11];
  assign T1776[10] = T1780[10] | T1777[10];
  assign T1776[9] = T1780[9] | T1777[9];
  assign T1776[8] = T1780[8] | T1777[8];
  assign T1776[7] = T1780[7] | T1777[7];
  assign T1776[6] = T1780[6] | T1777[6];
  assign T1776[5] = T1780[5] | T1777[5];
  assign T1776[4] = T1780[4] | T1777[4];
  assign T1776[3] = T1780[3] | T1777[3];
  assign T1776[2] = T1780[2] | T1777[2];
  assign T1776[1] = T1780[1] | T1777[1];
  assign T1776[0] = T1780[0] | T1777[0];
  assign T1780[11] = T1784[11] | T1781[11];
  assign T1780[10] = T1784[10] | T1781[10];
  assign T1780[9] = T1784[9] | T1781[9];
  assign T1780[8] = T1784[8] | T1781[8];
  assign T1780[7] = T1784[7] | T1781[7];
  assign T1780[6] = T1784[6] | T1781[6];
  assign T1780[5] = T1784[5] | T1781[5];
  assign T1780[4] = T1784[4] | T1781[4];
  assign T1780[3] = T1784[3] | T1781[3];
  assign T1780[2] = T1784[2] | T1781[2];
  assign T1780[1] = T1784[1] | T1781[1];
  assign T1780[0] = T1784[0] | T1781[0];
  assign T1536[38] = T1976[26] | T1788[26];
  assign T1536[37] = T1976[25] | T1788[25];
  assign T1536[36] = T1976[24] | T1788[24];
  assign T1536[35] = T1976[23] | T1788[23];
  assign T1536[34] = T1976[22] | T1788[22];
  assign T1536[33] = T1976[21] | T1788[21];
  assign T1536[32] = T1976[20] | T1788[20];
  assign T1536[31] = T1976[19] | T1788[19];
  assign T1536[30] = T1976[18] | T1788[18];
  assign T1536[29] = T1976[17] | T1788[17];
  assign T1536[28] = T1976[16] | T1788[16];
  assign T1536[27] = T1976[15] | T1788[15];
  assign T1536[26] = T1976[14] | T1788[14];
  assign T1536[25] = T1976[13] | T1788[13];
  assign T1536[24] = T1976[12] | T1788[12];
  assign T1536[23] = T1976[11] | T1788[11];
  assign T1536[22] = T1976[10] | T1788[10];
  assign T1536[21] = T1976[9] | T1788[9];
  assign T1536[20] = T1976[8] | T1788[8];
  assign T1536[19] = T1976[7] | T1788[7];
  assign T1536[18] = T1976[6] | T1788[6];
  assign T1536[17] = T1976[5] | T1788[5];
  assign T1536[16] = T1976[4] | T1788[4];
  assign T1536[15] = T1976[3] | T1788[3];
  assign T1536[14] = T1976[2] | T1788[2];
  assign T1536[13] = T1976[1] | T1788[1];
  assign T1536[12] = T1976[0] | T1788[0];
  assign N1013 = ~T1791[5];
  assign T1791[5] = T1794[5] | T1792[5];
  assign T1791[4] = T1794[4] | T1792[4];
  assign T1791[3] = T1794[3] | T1792[3];
  assign T1791[2] = T1794[2] | T1792[2];
  assign T1791[1] = T1794[1] | T1792[1];
  assign T1791[0] = T1794[0] | T1792[0];
  assign T1794[5] = T1797[5] | T1795[5];
  assign T1794[4] = T1797[4] | T1795[4];
  assign T1794[3] = T1797[3] | T1795[3];
  assign T1794[2] = T1797[2] | T1795[2];
  assign T1794[1] = T1797[1] | T1795[1];
  assign T1794[0] = T1797[0] | T1795[0];
  assign T1797[5] = T1800[5] | T1798[5];
  assign T1797[4] = T1800[4] | T1798[4];
  assign T1797[3] = T1800[3] | T1798[3];
  assign T1797[2] = T1800[2] | T1798[2];
  assign T1797[1] = T1800[1] | T1798[1];
  assign T1797[0] = T1800[0] | T1798[0];
  assign T1800[5] = T1803[5] | T1801[5];
  assign T1800[4] = T1803[4] | T1801[4];
  assign T1800[3] = T1803[3] | T1801[3];
  assign T1800[2] = T1803[2] | T1801[2];
  assign T1800[1] = T1803[1] | T1801[1];
  assign T1800[0] = T1803[0] | T1801[0];
  assign T1803[5] = T1806[5] | T1804[5];
  assign T1803[4] = T1806[4] | T1804[4];
  assign T1803[3] = T1806[3] | T1804[3];
  assign T1803[2] = T1806[2] | T1804[2];
  assign T1803[1] = T1806[1] | T1804[1];
  assign T1803[0] = T1806[0] | T1804[0];
  assign T1806[5] = T1809[5] | T1807[5];
  assign T1806[4] = T1809[4] | T1807[4];
  assign T1806[3] = T1809[3] | T1807[3];
  assign T1806[2] = T1809[2] | T1807[2];
  assign T1806[1] = T1809[1] | T1807[1];
  assign T1806[0] = T1809[0] | T1807[0];
  assign T1809[5] = T1812[5] | T1810[5];
  assign T1809[4] = T1812[4] | T1810[4];
  assign T1809[3] = T1812[3] | T1810[3];
  assign T1809[2] = T1812[2] | T1810[2];
  assign T1809[1] = T1812[1] | T1810[1];
  assign T1809[0] = T1812[0] | T1810[0];
  assign T1812[5] = T1815[5] | T1813[5];
  assign T1812[4] = T1815[4] | T1813[4];
  assign T1812[3] = T1815[3] | T1813[3];
  assign T1812[2] = T1815[2] | T1813[2];
  assign T1812[1] = T1815[1] | T1813[1];
  assign T1812[0] = T1815[0] | T1813[0];
  assign T1815[5] = T1818[5] | T1816[5];
  assign T1815[4] = T1818[4] | T1816[4];
  assign T1815[3] = T1818[3] | T1816[3];
  assign T1815[2] = T1818[2] | T1816[2];
  assign T1815[1] = T1818[1] | T1816[1];
  assign T1815[0] = T1818[0] | T1816[0];
  assign T1818[5] = T1821[5] | T1819[5];
  assign T1818[4] = T1821[4] | T1819[4];
  assign T1818[3] = T1821[3] | T1819[3];
  assign T1818[2] = T1821[2] | T1819[2];
  assign T1818[1] = T1821[1] | T1819[1];
  assign T1818[0] = T1821[0] | T1819[0];
  assign T1821[5] = T1824[5] | T1822[5];
  assign T1821[4] = T1824[4] | T1822[4];
  assign T1821[3] = T1824[3] | T1822[3];
  assign T1821[2] = T1824[2] | T1822[2];
  assign T1821[1] = T1824[1] | T1822[1];
  assign T1821[0] = T1824[0] | T1822[0];
  assign T1824[5] = T1827[5] | T1825[5];
  assign T1824[4] = T1827[4] | T1825[4];
  assign T1824[3] = T1827[3] | T1825[3];
  assign T1824[2] = T1827[2] | T1825[2];
  assign T1824[1] = T1827[1] | T1825[1];
  assign T1824[0] = T1827[0] | T1825[0];
  assign T1827[5] = T1830[5] | T1828[5];
  assign T1827[4] = T1830[4] | T1828[4];
  assign T1827[3] = T1830[3] | T1828[3];
  assign T1827[2] = T1830[2] | T1828[2];
  assign T1827[1] = T1830[1] | T1828[1];
  assign T1827[0] = T1830[0] | T1828[0];
  assign T1830[5] = T1833[5] | T1831[5];
  assign T1830[4] = T1833[4] | T1831[4];
  assign T1830[3] = T1833[3] | T1831[3];
  assign T1830[2] = T1833[2] | T1831[2];
  assign T1830[1] = T1833[1] | T1831[1];
  assign T1830[0] = T1833[0] | T1831[0];
  assign T1833[5] = T1836[5] | T1834[5];
  assign T1833[4] = T1836[4] | T1834[4];
  assign T1833[3] = T1836[3] | T1834[3];
  assign T1833[2] = T1836[2] | T1834[2];
  assign T1833[1] = T1836[1] | T1834[1];
  assign T1833[0] = T1836[0] | T1834[0];
  assign T1836[5] = T1839[5] | T1837[5];
  assign T1836[4] = T1839[4] | T1837[4];
  assign T1836[3] = T1839[3] | T1837[3];
  assign T1836[2] = T1839[2] | T1837[2];
  assign T1836[1] = T1839[1] | T1837[1];
  assign T1836[0] = T1839[0] | T1837[0];
  assign T1839[5] = T1842[5] | T1840[5];
  assign T1839[4] = T1842[4] | T1840[4];
  assign T1839[3] = T1842[3] | T1840[3];
  assign T1839[2] = T1842[2] | T1840[2];
  assign T1839[1] = T1842[1] | T1840[1];
  assign T1839[0] = T1842[0] | T1840[0];
  assign T1842[5] = T1845[5] | T1843[5];
  assign T1842[4] = T1845[4] | T1843[4];
  assign T1842[3] = T1845[3] | T1843[3];
  assign T1842[2] = T1845[2] | T1843[2];
  assign T1842[1] = T1845[1] | T1843[1];
  assign T1842[0] = T1845[0] | T1843[0];
  assign T1845[5] = T1848[5] | T1846[5];
  assign T1845[4] = T1848[4] | T1846[4];
  assign T1845[3] = T1848[3] | T1846[3];
  assign T1845[2] = T1848[2] | T1846[2];
  assign T1845[1] = T1848[1] | T1846[1];
  assign T1845[0] = T1848[0] | T1846[0];
  assign T1848[5] = T1851[5] | T1849[5];
  assign T1848[4] = T1851[4] | T1849[4];
  assign T1848[3] = T1851[3] | T1849[3];
  assign T1848[2] = T1851[2] | T1849[2];
  assign T1848[1] = T1851[1] | T1849[1];
  assign T1848[0] = T1851[0] | T1849[0];
  assign T1851[5] = T1854[5] | T1852[5];
  assign T1851[4] = T1854[4] | T1852[4];
  assign T1851[3] = T1854[3] | T1852[3];
  assign T1851[2] = T1854[2] | T1852[2];
  assign T1851[1] = T1854[1] | T1852[1];
  assign T1851[0] = T1854[0] | T1852[0];
  assign T1854[5] = T1857[5] | T1855[5];
  assign T1854[4] = T1857[4] | T1855[4];
  assign T1854[3] = T1857[3] | T1855[3];
  assign T1854[2] = T1857[2] | T1855[2];
  assign T1854[1] = T1857[1] | T1855[1];
  assign T1854[0] = T1857[0] | T1855[0];
  assign T1857[5] = T1860[5] | T1858[5];
  assign T1857[4] = T1860[4] | T1858[4];
  assign T1857[3] = T1860[3] | T1858[3];
  assign T1857[2] = T1860[2] | T1858[2];
  assign T1857[1] = T1860[1] | T1858[1];
  assign T1857[0] = T1860[0] | T1858[0];
  assign T1860[5] = T1863[5] | T1861[5];
  assign T1860[4] = T1863[4] | T1861[4];
  assign T1860[3] = T1863[3] | T1861[3];
  assign T1860[2] = T1863[2] | T1861[2];
  assign T1860[1] = T1863[1] | T1861[1];
  assign T1860[0] = T1863[0] | T1861[0];
  assign T1863[5] = T1866[5] | T1864[5];
  assign T1863[4] = T1866[4] | T1864[4];
  assign T1863[3] = T1866[3] | T1864[3];
  assign T1863[2] = T1866[2] | T1864[2];
  assign T1863[1] = T1866[1] | T1864[1];
  assign T1863[0] = T1866[0] | T1864[0];
  assign T1866[5] = T1869[5] | T1867[5];
  assign T1866[4] = T1869[4] | T1867[4];
  assign T1866[3] = T1869[3] | T1867[3];
  assign T1866[2] = T1869[2] | T1867[2];
  assign T1866[1] = T1869[1] | T1867[1];
  assign T1866[0] = T1869[0] | T1867[0];
  assign T1869[5] = T1872[5] | T1870[5];
  assign T1869[4] = T1872[4] | T1870[4];
  assign T1869[3] = T1872[3] | T1870[3];
  assign T1869[2] = T1872[2] | T1870[2];
  assign T1869[1] = T1872[1] | T1870[1];
  assign T1869[0] = T1872[0] | T1870[0];
  assign T1872[5] = T1875[5] | T1873[5];
  assign T1872[4] = T1875[4] | T1873[4];
  assign T1872[3] = T1875[3] | T1873[3];
  assign T1872[2] = T1875[2] | T1873[2];
  assign T1872[1] = T1875[1] | T1873[1];
  assign T1872[0] = T1875[0] | T1873[0];
  assign T1875[5] = T1878[5] | T1876[5];
  assign T1875[4] = T1878[4] | T1876[4];
  assign T1875[3] = T1878[3] | T1876[3];
  assign T1875[2] = T1878[2] | T1876[2];
  assign T1875[1] = T1878[1] | T1876[1];
  assign T1875[0] = T1878[0] | T1876[0];
  assign T1878[5] = T1881[5] | T1879[5];
  assign T1878[4] = T1881[4] | T1879[4];
  assign T1878[3] = T1881[3] | T1879[3];
  assign T1878[2] = T1881[2] | T1879[2];
  assign T1878[1] = T1881[1] | T1879[1];
  assign T1878[0] = T1881[0] | T1879[0];
  assign T1881[5] = T1884[5] | T1882[5];
  assign T1881[4] = T1884[4] | T1882[4];
  assign T1881[3] = T1884[3] | T1882[3];
  assign T1881[2] = T1884[2] | T1882[2];
  assign T1881[1] = T1884[1] | T1882[1];
  assign T1881[0] = T1884[0] | T1882[0];
  assign T1884[5] = T1887[5] | T1885[5];
  assign T1884[4] = T1887[4] | T1885[4];
  assign T1884[3] = T1887[3] | T1885[3];
  assign T1884[2] = T1887[2] | T1885[2];
  assign T1884[1] = T1887[1] | T1885[1];
  assign T1884[0] = T1887[0] | T1885[0];
  assign T1887[5] = T1890[5] | T1888[5];
  assign T1887[4] = T1890[4] | T1888[4];
  assign T1887[3] = T1890[3] | T1888[3];
  assign T1887[2] = T1890[2] | T1888[2];
  assign T1887[1] = T1890[1] | T1888[1];
  assign T1887[0] = T1890[0] | T1888[0];
  assign T1890[5] = T1893[5] | T1891[5];
  assign T1890[4] = T1893[4] | T1891[4];
  assign T1890[3] = T1893[3] | T1891[3];
  assign T1890[2] = T1893[2] | T1891[2];
  assign T1890[1] = T1893[1] | T1891[1];
  assign T1890[0] = T1893[0] | T1891[0];
  assign T1893[5] = T1896[5] | T1894[5];
  assign T1893[4] = T1896[4] | T1894[4];
  assign T1893[3] = T1896[3] | T1894[3];
  assign T1893[2] = T1896[2] | T1894[2];
  assign T1893[1] = T1896[1] | T1894[1];
  assign T1893[0] = T1896[0] | T1894[0];
  assign T1896[5] = T1899[5] | T1897[5];
  assign T1896[4] = T1899[4] | T1897[4];
  assign T1896[3] = T1899[3] | T1897[3];
  assign T1896[2] = T1899[2] | T1897[2];
  assign T1896[1] = T1899[1] | T1897[1];
  assign T1896[0] = T1899[0] | T1897[0];
  assign T1899[5] = T1902[5] | T1900[5];
  assign T1899[4] = T1902[4] | T1900[4];
  assign T1899[3] = T1902[3] | T1900[3];
  assign T1899[2] = T1902[2] | T1900[2];
  assign T1899[1] = T1902[1] | T1900[1];
  assign T1899[0] = T1902[0] | T1900[0];
  assign T1902[5] = T1905[5] | T1903[5];
  assign T1902[4] = T1905[4] | T1903[4];
  assign T1902[3] = T1905[3] | T1903[3];
  assign T1902[2] = T1905[2] | T1903[2];
  assign T1902[1] = T1905[1] | T1903[1];
  assign T1902[0] = T1905[0] | T1903[0];
  assign T1905[5] = T1908[5] | T1906[5];
  assign T1905[4] = T1908[4] | T1906[4];
  assign T1905[3] = T1908[3] | T1906[3];
  assign T1905[2] = T1908[2] | T1906[2];
  assign T1905[1] = T1908[1] | T1906[1];
  assign T1905[0] = T1908[0] | T1906[0];
  assign T1908[5] = T1911[5] | T1909[5];
  assign T1908[4] = T1911[4] | T1909[4];
  assign T1908[3] = T1911[3] | T1909[3];
  assign T1908[2] = T1911[2] | T1909[2];
  assign T1908[1] = T1911[1] | T1909[1];
  assign T1908[0] = T1911[0] | T1909[0];
  assign T1911[5] = T1914[5] | T1912[5];
  assign T1911[4] = T1914[4] | T1912[4];
  assign T1911[3] = T1914[3] | T1912[3];
  assign T1911[2] = T1914[2] | T1912[2];
  assign T1911[1] = T1914[1] | T1912[1];
  assign T1911[0] = T1914[0] | T1912[0];
  assign T1914[5] = T1917[5] | T1915[5];
  assign T1914[4] = T1917[4] | T1915[4];
  assign T1914[3] = T1917[3] | T1915[3];
  assign T1914[2] = T1917[2] | T1915[2];
  assign T1914[1] = T1917[1] | T1915[1];
  assign T1914[0] = T1917[0] | T1915[0];
  assign T1917[5] = T1920[5] | T1918[5];
  assign T1917[4] = T1920[4] | T1918[4];
  assign T1917[3] = T1920[3] | T1918[3];
  assign T1917[2] = T1920[2] | T1918[2];
  assign T1917[1] = T1920[1] | T1918[1];
  assign T1917[0] = T1920[0] | T1918[0];
  assign T1920[5] = T1923[5] | T1921[5];
  assign T1920[4] = T1923[4] | T1921[4];
  assign T1920[3] = T1923[3] | T1921[3];
  assign T1920[2] = T1923[2] | T1921[2];
  assign T1920[1] = T1923[1] | T1921[1];
  assign T1920[0] = T1923[0] | T1921[0];
  assign T1923[5] = T1926[5] | T1924[5];
  assign T1923[4] = T1926[4] | T1924[4];
  assign T1923[3] = T1926[3] | T1924[3];
  assign T1923[2] = T1926[2] | T1924[2];
  assign T1923[1] = T1926[1] | T1924[1];
  assign T1923[0] = T1926[0] | T1924[0];
  assign T1926[5] = T1929[5] | T1927[5];
  assign T1926[4] = T1929[4] | T1927[4];
  assign T1926[3] = T1929[3] | T1927[3];
  assign T1926[2] = T1929[2] | T1927[2];
  assign T1926[1] = T1929[1] | T1927[1];
  assign T1926[0] = T1929[0] | T1927[0];
  assign T1929[5] = T1932[5] | T1930[5];
  assign T1929[4] = T1932[4] | T1930[4];
  assign T1929[3] = T1932[3] | T1930[3];
  assign T1929[2] = T1932[2] | T1930[2];
  assign T1929[1] = T1932[1] | T1930[1];
  assign T1929[0] = T1932[0] | T1930[0];
  assign T1932[5] = T1935[5] | T1933[5];
  assign T1932[4] = T1935[4] | T1933[4];
  assign T1932[3] = T1935[3] | T1933[3];
  assign T1932[2] = T1935[2] | T1933[2];
  assign T1932[1] = T1935[1] | T1933[1];
  assign T1932[0] = T1935[0] | T1933[0];
  assign T1935[5] = T1938[5] | T1936[5];
  assign T1935[4] = T1938[4] | T1936[4];
  assign T1935[3] = T1938[3] | T1936[3];
  assign T1935[2] = T1938[2] | T1936[2];
  assign T1935[1] = T1938[1] | T1936[1];
  assign T1935[0] = T1938[0] | T1936[0];
  assign T1938[5] = T1941[5] | T1939[5];
  assign T1938[4] = T1941[4] | T1939[4];
  assign T1938[3] = T1941[3] | T1939[3];
  assign T1938[2] = T1941[2] | T1939[2];
  assign T1938[1] = T1941[1] | T1939[1];
  assign T1938[0] = T1941[0] | T1939[0];
  assign T1941[5] = T1944[5] | T1942[5];
  assign T1941[4] = T1944[4] | T1942[4];
  assign T1941[3] = T1944[3] | T1942[3];
  assign T1941[2] = T1944[2] | T1942[2];
  assign T1941[1] = T1944[1] | T1942[1];
  assign T1941[0] = T1944[0] | T1942[0];
  assign T1944[5] = T1947[5] | T1945[5];
  assign T1944[4] = T1947[4] | T1945[4];
  assign T1944[3] = T1947[3] | T1945[3];
  assign T1944[2] = T1947[2] | T1945[2];
  assign T1944[1] = T1947[1] | T1945[1];
  assign T1944[0] = T1947[0] | T1945[0];
  assign T1947[5] = T1950[5] | T1948[5];
  assign T1947[4] = T1950[4] | T1948[4];
  assign T1947[3] = T1950[3] | T1948[3];
  assign T1947[2] = T1950[2] | T1948[2];
  assign T1947[1] = T1950[1] | T1948[1];
  assign T1947[0] = T1950[0] | T1948[0];
  assign T1950[5] = T1953[5] | T1951[5];
  assign T1950[4] = T1953[4] | T1951[4];
  assign T1950[3] = T1953[3] | T1951[3];
  assign T1950[2] = T1953[2] | T1951[2];
  assign T1950[1] = T1953[1] | T1951[1];
  assign T1950[0] = T1953[0] | T1951[0];
  assign T1953[5] = T1956[5] | T1954[5];
  assign T1953[4] = T1956[4] | T1954[4];
  assign T1953[3] = T1956[3] | T1954[3];
  assign T1953[2] = T1956[2] | T1954[2];
  assign T1953[1] = T1956[1] | T1954[1];
  assign T1953[0] = T1956[0] | T1954[0];
  assign T1956[5] = T1959[5] | T1957[5];
  assign T1956[4] = T1959[4] | T1957[4];
  assign T1956[3] = T1959[3] | T1957[3];
  assign T1956[2] = T1959[2] | T1957[2];
  assign T1956[1] = T1959[1] | T1957[1];
  assign T1956[0] = T1959[0] | T1957[0];
  assign T1959[5] = T1962[5] | T1960[5];
  assign T1959[4] = T1962[4] | T1960[4];
  assign T1959[3] = T1962[3] | T1960[3];
  assign T1959[2] = T1962[2] | T1960[2];
  assign T1959[1] = T1962[1] | T1960[1];
  assign T1959[0] = T1962[0] | T1960[0];
  assign T1962[5] = T1965[5] | T1963[5];
  assign T1962[4] = T1965[4] | T1963[4];
  assign T1962[3] = T1965[3] | T1963[3];
  assign T1962[2] = T1965[2] | T1963[2];
  assign T1962[1] = T1965[1] | T1963[1];
  assign T1962[0] = T1965[0] | T1963[0];
  assign T1965[5] = T1968[5] | T1966[5];
  assign T1965[4] = T1968[4] | T1966[4];
  assign T1965[3] = T1968[3] | T1966[3];
  assign T1965[2] = T1968[2] | T1966[2];
  assign T1965[1] = T1968[1] | T1966[1];
  assign T1965[0] = T1968[0] | T1966[0];
  assign T1968[5] = T1971[5] | T1969[5];
  assign T1968[4] = T1971[4] | T1969[4];
  assign T1968[3] = T1971[3] | T1969[3];
  assign T1968[2] = T1971[2] | T1969[2];
  assign T1968[1] = T1971[1] | T1969[1];
  assign T1968[0] = T1971[0] | T1969[0];
  assign T1971[5] = T1974[5] | T1972[5];
  assign T1971[4] = T1974[4] | T1972[4];
  assign T1971[3] = T1974[3] | T1972[3];
  assign T1971[2] = T1974[2] | T1972[2];
  assign T1971[1] = T1974[1] | T1972[1];
  assign T1971[0] = T1974[0] | T1972[0];
  assign T1976[26] = T1980[26] | T1977[26];
  assign T1976[25] = T1980[25] | T1977[25];
  assign T1976[24] = T1980[24] | T1977[24];
  assign T1976[23] = T1980[23] | T1977[23];
  assign T1976[22] = T1980[22] | T1977[22];
  assign T1976[21] = T1980[21] | T1977[21];
  assign T1976[20] = T1980[20] | T1977[20];
  assign T1976[19] = T1980[19] | T1977[19];
  assign T1976[18] = T1980[18] | T1977[18];
  assign T1976[17] = T1980[17] | T1977[17];
  assign T1976[16] = T1980[16] | T1977[16];
  assign T1976[15] = T1980[15] | T1977[15];
  assign T1976[14] = T1980[14] | T1977[14];
  assign T1976[13] = T1980[13] | T1977[13];
  assign T1976[12] = T1980[12] | T1977[12];
  assign T1976[11] = T1980[11] | T1977[11];
  assign T1976[10] = T1980[10] | T1977[10];
  assign T1976[9] = T1980[9] | T1977[9];
  assign T1976[8] = T1980[8] | T1977[8];
  assign T1976[7] = T1980[7] | T1977[7];
  assign T1976[6] = T1980[6] | T1977[6];
  assign T1976[5] = T1980[5] | T1977[5];
  assign T1976[4] = T1980[4] | T1977[4];
  assign T1976[3] = T1980[3] | T1977[3];
  assign T1976[2] = T1980[2] | T1977[2];
  assign T1976[1] = T1980[1] | T1977[1];
  assign T1976[0] = T1980[0] | T1977[0];
  assign N1014 = ~T1791[4];
  assign T1980[26] = T1984[26] | T1981[26];
  assign T1980[25] = T1984[25] | T1981[25];
  assign T1980[24] = T1984[24] | T1981[24];
  assign T1980[23] = T1984[23] | T1981[23];
  assign T1980[22] = T1984[22] | T1981[22];
  assign T1980[21] = T1984[21] | T1981[21];
  assign T1980[20] = T1984[20] | T1981[20];
  assign T1980[19] = T1984[19] | T1981[19];
  assign T1980[18] = T1984[18] | T1981[18];
  assign T1980[17] = T1984[17] | T1981[17];
  assign T1980[16] = T1984[16] | T1981[16];
  assign T1980[15] = T1984[15] | T1981[15];
  assign T1980[14] = T1984[14] | T1981[14];
  assign T1980[13] = T1984[13] | T1981[13];
  assign T1980[12] = T1984[12] | T1981[12];
  assign T1980[11] = T1984[11] | T1981[11];
  assign T1980[10] = T1984[10] | T1981[10];
  assign T1980[9] = T1984[9] | T1981[9];
  assign T1980[8] = T1984[8] | T1981[8];
  assign T1980[7] = T1984[7] | T1981[7];
  assign T1980[6] = T1984[6] | T1981[6];
  assign T1980[5] = T1984[5] | T1981[5];
  assign T1980[4] = T1984[4] | T1981[4];
  assign T1980[3] = T1984[3] | T1981[3];
  assign T1980[2] = T1984[2] | T1981[2];
  assign T1980[1] = T1984[1] | T1981[1];
  assign T1980[0] = T1984[0] | T1981[0];
  assign N1015 = ~T1791[3];
  assign T1984[26] = T1988[26] | T1985[26];
  assign T1984[25] = T1988[25] | T1985[25];
  assign T1984[24] = T1988[24] | T1985[24];
  assign T1984[23] = T1988[23] | T1985[23];
  assign T1984[22] = T1988[22] | T1985[22];
  assign T1984[21] = T1988[21] | T1985[21];
  assign T1984[20] = T1988[20] | T1985[20];
  assign T1984[19] = T1988[19] | T1985[19];
  assign T1984[18] = T1988[18] | T1985[18];
  assign T1984[17] = T1988[17] | T1985[17];
  assign T1984[16] = T1988[16] | T1985[16];
  assign T1984[15] = T1988[15] | T1985[15];
  assign T1984[14] = T1988[14] | T1985[14];
  assign T1984[13] = T1988[13] | T1985[13];
  assign T1984[12] = T1988[12] | T1985[12];
  assign T1984[11] = T1988[11] | T1985[11];
  assign T1984[10] = T1988[10] | T1985[10];
  assign T1984[9] = T1988[9] | T1985[9];
  assign T1984[8] = T1988[8] | T1985[8];
  assign T1984[7] = T1988[7] | T1985[7];
  assign T1984[6] = T1988[6] | T1985[6];
  assign T1984[5] = T1988[5] | T1985[5];
  assign T1984[4] = T1988[4] | T1985[4];
  assign T1984[3] = T1988[3] | T1985[3];
  assign T1984[2] = T1988[2] | T1985[2];
  assign T1984[1] = T1988[1] | T1985[1];
  assign T1984[0] = T1988[0] | T1985[0];
  assign N1016 = ~T1791[2];
  assign T1988[26] = T1992[26] | T1989[26];
  assign T1988[25] = T1992[25] | T1989[25];
  assign T1988[24] = T1992[24] | T1989[24];
  assign T1988[23] = T1992[23] | T1989[23];
  assign T1988[22] = T1992[22] | T1989[22];
  assign T1988[21] = T1992[21] | T1989[21];
  assign T1988[20] = T1992[20] | T1989[20];
  assign T1988[19] = T1992[19] | T1989[19];
  assign T1988[18] = T1992[18] | T1989[18];
  assign T1988[17] = T1992[17] | T1989[17];
  assign T1988[16] = T1992[16] | T1989[16];
  assign T1988[15] = T1992[15] | T1989[15];
  assign T1988[14] = T1992[14] | T1989[14];
  assign T1988[13] = T1992[13] | T1989[13];
  assign T1988[12] = T1992[12] | T1989[12];
  assign T1988[11] = T1992[11] | T1989[11];
  assign T1988[10] = T1992[10] | T1989[10];
  assign T1988[9] = T1992[9] | T1989[9];
  assign T1988[8] = T1992[8] | T1989[8];
  assign T1988[7] = T1992[7] | T1989[7];
  assign T1988[6] = T1992[6] | T1989[6];
  assign T1988[5] = T1992[5] | T1989[5];
  assign T1988[4] = T1992[4] | T1989[4];
  assign T1988[3] = T1992[3] | T1989[3];
  assign T1988[2] = T1992[2] | T1989[2];
  assign T1988[1] = T1992[1] | T1989[1];
  assign T1988[0] = T1992[0] | T1989[0];
  assign N1017 = ~T1791[1];
  assign N1018 = ~T1791[0];
  assign N1019 = ~T2027;
  assign T1998 = T2022 & T2000[0];
  assign T2007 = T2018 & T2008;
  assign T2008 = ~N2777;
  assign T2015 = T2022 & T2016;
  assign T2016 = ~R2010[1];
  assign T2018 = io_ras_update_valid & T2019;
  assign T2019 = T2021 & T2020;
  assign T2020 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T2021 = ~io_ras_update_bits_isCall;
  assign T2022 = io_ras_update_valid & io_ras_update_bits_isCall;
  assign T2025 = T2022 & T2000[1];
  assign T2028 = T2404 & T2029;
  assign T2029 = T2039 | T2030;
  assign T2034 = R7 & T2036[61];
  assign T2039 = T2045 | T2040;
  assign T2042 = R7 & T2036[60];
  assign T2045 = T2051 | T2046;
  assign T2048 = R7 & T2036[59];
  assign T2051 = T2057 | T2052;
  assign T2054 = R7 & T2036[58];
  assign T2057 = T2063 | T2058;
  assign T2060 = R7 & T2036[57];
  assign T2063 = T2069 | T2064;
  assign T2066 = R7 & T2036[56];
  assign T2069 = T2075 | T2070;
  assign T2072 = R7 & T2036[55];
  assign T2075 = T2081 | T2076;
  assign T2078 = R7 & T2036[54];
  assign T2081 = T2087 | T2082;
  assign T2084 = R7 & T2036[53];
  assign T2087 = T2093 | T2088;
  assign T2090 = R7 & T2036[52];
  assign T2093 = T2099 | T2094;
  assign T2096 = R7 & T2036[51];
  assign T2099 = T2105 | T2100;
  assign T2102 = R7 & T2036[50];
  assign T2105 = T2111 | T2106;
  assign T2108 = R7 & T2036[49];
  assign T2111 = T2117 | T2112;
  assign T2114 = R7 & T2036[48];
  assign T2117 = T2123 | T2118;
  assign T2120 = R7 & T2036[47];
  assign T2123 = T2129 | T2124;
  assign T2126 = R7 & T2036[46];
  assign T2129 = T2135 | T2130;
  assign T2132 = R7 & T2036[45];
  assign T2135 = T2141 | T2136;
  assign T2138 = R7 & T2036[44];
  assign T2141 = T2147 | T2142;
  assign T2144 = R7 & T2036[43];
  assign T2147 = T2153 | T2148;
  assign T2150 = R7 & T2036[42];
  assign T2153 = T2159 | T2154;
  assign T2156 = R7 & T2036[41];
  assign T2159 = T2165 | T2160;
  assign T2162 = R7 & T2036[40];
  assign T2165 = T2171 | T2166;
  assign T2168 = R7 & T2036[39];
  assign T2171 = T2177 | T2172;
  assign T2174 = R7 & T2036[38];
  assign T2177 = T2183 | T2178;
  assign T2180 = R7 & T2036[37];
  assign T2183 = T2189 | T2184;
  assign T2186 = R7 & T2036[36];
  assign T2189 = T2195 | T2190;
  assign T2192 = R7 & T2036[35];
  assign T2195 = T2201 | T2196;
  assign T2198 = R7 & T2036[34];
  assign T2201 = T2207 | T2202;
  assign T2204 = R7 & T2036[33];
  assign T2207 = T2213 | T2208;
  assign T2210 = R7 & T2036[32];
  assign T2213 = T2219 | T2214;
  assign T2216 = R7 & T2036[31];
  assign T2219 = T2225 | T2220;
  assign T2222 = R7 & T2036[30];
  assign T2225 = T2231 | T2226;
  assign T2228 = R7 & T2036[29];
  assign T2231 = T2237 | T2232;
  assign T2234 = R7 & T2036[28];
  assign T2237 = T2243 | T2238;
  assign T2240 = R7 & T2036[27];
  assign T2243 = T2249 | T2244;
  assign T2246 = R7 & T2036[26];
  assign T2249 = T2255 | T2250;
  assign T2252 = R7 & T2036[25];
  assign T2255 = T2261 | T2256;
  assign T2258 = R7 & T2036[24];
  assign T2261 = T2267 | T2262;
  assign T2264 = R7 & T2036[23];
  assign T2267 = T2273 | T2268;
  assign T2270 = R7 & T2036[22];
  assign T2273 = T2279 | T2274;
  assign T2276 = R7 & T2036[21];
  assign T2279 = T2285 | T2280;
  assign T2282 = R7 & T2036[20];
  assign T2285 = T2291 | T2286;
  assign T2288 = R7 & T2036[19];
  assign T2291 = T2297 | T2292;
  assign T2294 = R7 & T2036[18];
  assign T2297 = T2303 | T2298;
  assign T2300 = R7 & T2036[17];
  assign T2303 = T2309 | T2304;
  assign T2306 = R7 & T2036[16];
  assign T2309 = T2315 | T2310;
  assign T2312 = R7 & T2036[15];
  assign T2315 = T2321 | T2316;
  assign T2318 = R7 & T2036[14];
  assign T2321 = T2327 | T2322;
  assign T2324 = R7 & T2036[13];
  assign T2327 = T2333 | T2328;
  assign T2330 = R7 & T2036[12];
  assign T2333 = T2339 | T2334;
  assign T2336 = R7 & T2036[11];
  assign T2339 = T2345 | T2340;
  assign T2342 = R7 & T2036[10];
  assign T2345 = T2351 | T2346;
  assign T2348 = R7 & T2036[9];
  assign T2351 = T2357 | T2352;
  assign T2354 = R7 & T2036[8];
  assign T2357 = T2363 | T2358;
  assign T2360 = R7 & T2036[7];
  assign T2363 = T2369 | T2364;
  assign T2366 = R7 & T2036[6];
  assign T2369 = T2375 | T2370;
  assign T2372 = R7 & T2036[5];
  assign T2375 = T2381 | T2376;
  assign T2378 = R7 & T2036[4];
  assign T2381 = T2387 | T2382;
  assign T2384 = R7 & T2036[3];
  assign T2387 = T2393 | T2388;
  assign T2390 = R7 & T2036[2];
  assign T2393 = T2399 | T2394;
  assign T2396 = R7 & T2036[1];
  assign T2401 = R7 & T2036[0];
  assign T2404 = ~N2403;
  assign T2406 = T2022 & T2029;
  assign T2409 = R7 & T2410;
  assign N1082 = ~T2412;
  assign T2412 = T2413 & T160;
  assign T2413 = ~io_resp_bits_bht_value[0];
  assign N1083 = ~reset;
  assign N1085 = ~T21;
  assign N1635 = T1530 | reset;
  assign N1636 = T159 | N1635;
  assign N1637 = ~N1636;
  assign N1646 = T175 | reset;
  assign N1647 = ~N1646;
  assign N1655 = io_invalidate | reset;
  assign N1656 = T265 | N1655;
  assign N1657 = ~N1656;
  assign N1665 = T203 | reset;
  assign N1666 = ~N1665;
  assign N1671 = ~T288;
  assign N1796 = ~T601;
  assign N1921 = ~T800;
  assign N2046 = ~T1541;
  assign N2171 = T2007 | reset;
  assign N2172 = T2022 | N2171;
  assign N2173 = ~N2172;
  assign N2176 = T2007 | N1655;
  assign N2177 = T2015 | N2176;
  assign N2178 = ~N2177;
  assign N2182 = ~T2409;
  assign N2307 = T1530 & N2311;
  assign N2308 = ~T1530;
  assign N2309 = N2311 & N2308;
  assign N2310 = T159 & N2309;
  assign N2311 = ~reset;
  assign N2312 = T175 & N2311;
  assign N2313 = io_invalidate & N2311;
  assign N2314 = ~io_invalidate;
  assign N2315 = N2311 & N2314;
  assign N2316 = T265 & N2315;
  assign N2317 = T203 & N2311;
  assign N2318 = T2007 & N2311;
  assign N2319 = ~T2007;
  assign N2320 = N2311 & N2319;
  assign N2321 = T2022 & N2320;
  assign N2322 = T2007 & N2315;
  assign N2323 = N2315 & N2319;
  assign N2324 = T2015 & N2323;
  assign N2325 = N947 & N1083;
  assign N2326 = N948 & N2325;
  assign N2327 = ~N2326;

endmodule