module commit_stage
(
  clk_i,
  rst_ni,
  halt_i,
  flush_dcache_i,
  exception_o,
  dirty_fp_state_o,
  debug_mode_i,
  debug_req_i,
  single_step_i,
  commit_instr_i,
  commit_ack_o,
  waddr_o,
  wdata_o,
  we_gpr_o,
  we_fpr_o,
  amo_resp_i,
  pc_o,
  csr_op_o,
  csr_wdata_o,
  csr_rdata_i,
  csr_exception_i,
  csr_write_fflags_o,
  commit_lsu_o,
  commit_lsu_ready_i,
  amo_valid_commit_o,
  no_st_pending_i,
  commit_csr_o,
  fence_i_o,
  fence_o,
  flush_commit_o,
  sfence_vma_o
);

  output [128:0] exception_o;
  input [723:0] commit_instr_i;
  output [1:0] commit_ack_o;
  output [9:0] waddr_o;
  output [127:0] wdata_o;
  output [1:0] we_gpr_o;
  output [1:0] we_fpr_o;
  input [64:0] amo_resp_i;
  output [63:0] pc_o;
  output [6:0] csr_op_o;
  output [63:0] csr_wdata_o;
  input [63:0] csr_rdata_i;
  input [128:0] csr_exception_i;
  input clk_i;
  input rst_ni;
  input halt_i;
  input flush_dcache_i;
  input debug_mode_i;
  input debug_req_i;
  input single_step_i;
  input commit_lsu_ready_i;
  input no_st_pending_i;
  output dirty_fp_state_o;
  output csr_write_fflags_o;
  output commit_lsu_o;
  output amo_valid_commit_o;
  output commit_csr_o;
  output fence_i_o;
  output fence_o;
  output flush_commit_o;
  output sfence_vma_o;
  wire [128:0] exception_o;
  wire [1:0] commit_ack_o,we_gpr_o,we_fpr_o;
  wire [9:0] waddr_o;
  wire [127:0] wdata_o;
  wire [63:0] pc_o,csr_wdata_o;
  wire [6:0] csr_op_o;
  wire dirty_fp_state_o,csr_write_fflags_o,commit_lsu_o,amo_valid_commit_o,
  commit_csr_o,fence_i_o,fence_o,flush_commit_o,sfence_vma_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,
  N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,
  N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,
  N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,
  N70,N71,N72,N73,N74,instr_0_is_amo,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,
  N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,
  N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,
  N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,
  N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,
  N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,
  N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,
  N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,
  N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,
  N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,
  N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,
  N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,
  N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,
  N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,
  N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,
  N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,
  N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,
  N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,
  N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,
  N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,
  N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
  N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,
  N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,
  N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,
  N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,
  N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,
  N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,
  N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,
  N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,
  N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,
  N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,
  N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,
  N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,
  N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,
  N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,
  N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,
  N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,
  N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,
  N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,
  N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,
  N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,
  N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,
  N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,
  N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,
  N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,
  N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,
  N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,
  N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,
  N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,
  N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,
  N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,
  N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,
  N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,
  N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,
  N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,
  N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,
  N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,
  N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,
  N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,
  N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,
  N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,
  N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,
  N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,
  N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,
  N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,
  N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,
  N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,
  N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,
  N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,
  N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,
  N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,
  N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187;
  assign we_fpr_o[0] = 1'b0;
  assign we_fpr_o[1] = 1'b0;
  assign pc_o[63] = commit_instr_i[361];
  assign pc_o[62] = commit_instr_i[360];
  assign pc_o[61] = commit_instr_i[359];
  assign pc_o[60] = commit_instr_i[358];
  assign pc_o[59] = commit_instr_i[357];
  assign pc_o[58] = commit_instr_i[356];
  assign pc_o[57] = commit_instr_i[355];
  assign pc_o[56] = commit_instr_i[354];
  assign pc_o[55] = commit_instr_i[353];
  assign pc_o[54] = commit_instr_i[352];
  assign pc_o[53] = commit_instr_i[351];
  assign pc_o[52] = commit_instr_i[350];
  assign pc_o[51] = commit_instr_i[349];
  assign pc_o[50] = commit_instr_i[348];
  assign pc_o[49] = commit_instr_i[347];
  assign pc_o[48] = commit_instr_i[346];
  assign pc_o[47] = commit_instr_i[345];
  assign pc_o[46] = commit_instr_i[344];
  assign pc_o[45] = commit_instr_i[343];
  assign pc_o[44] = commit_instr_i[342];
  assign pc_o[43] = commit_instr_i[341];
  assign pc_o[42] = commit_instr_i[340];
  assign pc_o[41] = commit_instr_i[339];
  assign pc_o[40] = commit_instr_i[338];
  assign pc_o[39] = commit_instr_i[337];
  assign pc_o[38] = commit_instr_i[336];
  assign pc_o[37] = commit_instr_i[335];
  assign pc_o[36] = commit_instr_i[334];
  assign pc_o[35] = commit_instr_i[333];
  assign pc_o[34] = commit_instr_i[332];
  assign pc_o[33] = commit_instr_i[331];
  assign pc_o[32] = commit_instr_i[330];
  assign pc_o[31] = commit_instr_i[329];
  assign pc_o[30] = commit_instr_i[328];
  assign pc_o[29] = commit_instr_i[327];
  assign pc_o[28] = commit_instr_i[326];
  assign pc_o[27] = commit_instr_i[325];
  assign pc_o[26] = commit_instr_i[324];
  assign pc_o[25] = commit_instr_i[323];
  assign pc_o[24] = commit_instr_i[322];
  assign pc_o[23] = commit_instr_i[321];
  assign pc_o[22] = commit_instr_i[320];
  assign pc_o[21] = commit_instr_i[319];
  assign pc_o[20] = commit_instr_i[318];
  assign pc_o[19] = commit_instr_i[317];
  assign pc_o[18] = commit_instr_i[316];
  assign pc_o[17] = commit_instr_i[315];
  assign pc_o[16] = commit_instr_i[314];
  assign pc_o[15] = commit_instr_i[313];
  assign pc_o[14] = commit_instr_i[312];
  assign pc_o[13] = commit_instr_i[311];
  assign pc_o[12] = commit_instr_i[310];
  assign pc_o[11] = commit_instr_i[309];
  assign pc_o[10] = commit_instr_i[308];
  assign pc_o[9] = commit_instr_i[307];
  assign pc_o[8] = commit_instr_i[306];
  assign pc_o[7] = commit_instr_i[305];
  assign pc_o[6] = commit_instr_i[304];
  assign pc_o[5] = commit_instr_i[303];
  assign pc_o[4] = commit_instr_i[302];
  assign pc_o[3] = commit_instr_i[301];
  assign pc_o[2] = commit_instr_i[300];
  assign pc_o[1] = commit_instr_i[299];
  assign pc_o[0] = commit_instr_i[298];
  assign waddr_o[9] = commit_instr_i[632];
  assign waddr_o[8] = commit_instr_i[631];
  assign waddr_o[7] = commit_instr_i[630];
  assign waddr_o[6] = commit_instr_i[629];
  assign waddr_o[5] = commit_instr_i[628];
  assign waddr_o[4] = commit_instr_i[270];
  assign waddr_o[3] = commit_instr_i[269];
  assign waddr_o[2] = commit_instr_i[268];
  assign waddr_o[1] = commit_instr_i[267];
  assign waddr_o[0] = commit_instr_i[266];
  assign wdata_o[127] = commit_instr_i[627];
  assign wdata_o[126] = commit_instr_i[626];
  assign wdata_o[125] = commit_instr_i[625];
  assign wdata_o[124] = commit_instr_i[624];
  assign wdata_o[123] = commit_instr_i[623];
  assign wdata_o[122] = commit_instr_i[622];
  assign wdata_o[121] = commit_instr_i[621];
  assign wdata_o[120] = commit_instr_i[620];
  assign wdata_o[119] = commit_instr_i[619];
  assign wdata_o[118] = commit_instr_i[618];
  assign wdata_o[117] = commit_instr_i[617];
  assign wdata_o[116] = commit_instr_i[616];
  assign wdata_o[115] = commit_instr_i[615];
  assign wdata_o[114] = commit_instr_i[614];
  assign wdata_o[113] = commit_instr_i[613];
  assign wdata_o[112] = commit_instr_i[612];
  assign wdata_o[111] = commit_instr_i[611];
  assign wdata_o[110] = commit_instr_i[610];
  assign wdata_o[109] = commit_instr_i[609];
  assign wdata_o[108] = commit_instr_i[608];
  assign wdata_o[107] = commit_instr_i[607];
  assign wdata_o[106] = commit_instr_i[606];
  assign wdata_o[105] = commit_instr_i[605];
  assign wdata_o[104] = commit_instr_i[604];
  assign wdata_o[103] = commit_instr_i[603];
  assign wdata_o[102] = commit_instr_i[602];
  assign wdata_o[101] = commit_instr_i[601];
  assign wdata_o[100] = commit_instr_i[600];
  assign wdata_o[99] = commit_instr_i[599];
  assign wdata_o[98] = commit_instr_i[598];
  assign wdata_o[97] = commit_instr_i[597];
  assign wdata_o[96] = commit_instr_i[596];
  assign wdata_o[95] = commit_instr_i[595];
  assign wdata_o[94] = commit_instr_i[594];
  assign wdata_o[93] = commit_instr_i[593];
  assign wdata_o[92] = commit_instr_i[592];
  assign wdata_o[91] = commit_instr_i[591];
  assign wdata_o[90] = commit_instr_i[590];
  assign wdata_o[89] = commit_instr_i[589];
  assign wdata_o[88] = commit_instr_i[588];
  assign wdata_o[87] = commit_instr_i[587];
  assign wdata_o[86] = commit_instr_i[586];
  assign wdata_o[85] = commit_instr_i[585];
  assign wdata_o[84] = commit_instr_i[584];
  assign wdata_o[83] = commit_instr_i[583];
  assign wdata_o[82] = commit_instr_i[582];
  assign wdata_o[81] = commit_instr_i[581];
  assign wdata_o[80] = commit_instr_i[580];
  assign wdata_o[79] = commit_instr_i[579];
  assign wdata_o[78] = commit_instr_i[578];
  assign wdata_o[77] = commit_instr_i[577];
  assign wdata_o[76] = commit_instr_i[576];
  assign wdata_o[75] = commit_instr_i[575];
  assign wdata_o[74] = commit_instr_i[574];
  assign wdata_o[73] = commit_instr_i[573];
  assign wdata_o[72] = commit_instr_i[572];
  assign wdata_o[71] = commit_instr_i[571];
  assign wdata_o[70] = commit_instr_i[570];
  assign wdata_o[69] = commit_instr_i[569];
  assign wdata_o[68] = commit_instr_i[568];
  assign wdata_o[67] = commit_instr_i[567];
  assign wdata_o[66] = commit_instr_i[566];
  assign wdata_o[65] = commit_instr_i[565];
  assign wdata_o[64] = commit_instr_i[564];
  assign N28 = commit_instr_i[290] | N74;
  assign N29 = commit_instr_i[288] | N1097;
  assign N30 = N1107 | commit_instr_i[285];
  assign N31 = N28 | N29;
  assign N32 = N30 | N1099;
  assign N33 = N31 | N32;
  assign N34 = N1107 | N1098;
  assign N35 = N34 | commit_instr_i[284];
  assign N36 = N31 | N35;
  assign N37 = N34 | N1099;
  assign N38 = N31 | N37;
  assign N39 = N1096 | commit_instr_i[287];
  assign N40 = commit_instr_i[286] | commit_instr_i[285];
  assign N41 = N28 | N39;
  assign N42 = N40 | commit_instr_i[284];
  assign N43 = N41 | N42;
  assign N44 = N40 | N1099;
  assign N45 = N41 | N44;
  assign N46 = commit_instr_i[286] | N1098;
  assign N47 = N46 | commit_instr_i[284];
  assign N48 = N41 | N47;
  assign N49 = N46 | N1099;
  assign N50 = N41 | N49;
  assign N51 = N30 | commit_instr_i[284];
  assign N52 = N41 | N51;
  assign N53 = N41 | N32;
  assign N54 = N41 | N35;
  assign N55 = N41 | N37;
  assign N56 = N1096 | N1097;
  assign N57 = N28 | N56;
  assign N58 = N57 | N42;
  assign N59 = N57 | N44;
  assign N60 = N57 | N47;
  assign N61 = N57 | N49;
  assign N62 = N57 | N51;
  assign N63 = N57 | N32;
  assign N64 = N57 | N35;
  assign N65 = N57 | N37;
  assign N66 = N73 | commit_instr_i[289];
  assign N67 = commit_instr_i[288] | commit_instr_i[287];
  assign N68 = N66 | N67;
  assign N69 = N68 | N42;
  assign N70 = N68 | N44;
  assign N71 = N68 | N47;
  assign N151 = N1091 | N150;
  assign N152 = N528 | N151;
  assign N154 = N153 | commit_instr_i[293];
  assign N155 = commit_instr_i[292] | commit_instr_i[291];
  assign N156 = N154 | N155;
  assign N528 = commit_instr_i[294] | N1090;
  assign N529 = N1091 | commit_instr_i[291];
  assign N530 = N528 | N529;
  assign N533 = commit_instr_i[656] | commit_instr_i[655];
  assign N534 = N533 | N546;
  assign N535 = commit_instr_i[654] | N544;
  assign N536 = N533 | N535;
  assign N537 = N545 | N550;
  assign N538 = N545 | N535;
  assign N545 = commit_instr_i[656] | N542;
  assign N546 = N543 | N544;
  assign N547 = N545 | N546;
  assign N549 = N548 | commit_instr_i[655];
  assign N550 = commit_instr_i[654] | commit_instr_i[653];
  assign N551 = N549 | N550;
  assign N1090 = ~commit_instr_i[293];
  assign N1091 = ~commit_instr_i[292];
  assign N1092 = N1090 | commit_instr_i[294];
  assign N1093 = N1091 | N1092;
  assign N1094 = commit_instr_i[291] | N1093;
  assign N1095 = ~N1094;
  assign N1096 = ~commit_instr_i[288];
  assign N1097 = ~commit_instr_i[287];
  assign N1098 = ~commit_instr_i[285];
  assign N1099 = ~commit_instr_i[284];
  assign N1100 = commit_instr_i[289] | commit_instr_i[290];
  assign N1101 = N1096 | N1100;
  assign N1102 = N1097 | N1101;
  assign N1103 = commit_instr_i[286] | N1102;
  assign N1104 = N1098 | N1103;
  assign N1105 = N1099 | N1104;
  assign N1106 = ~N1105;
  assign N1107 = ~commit_instr_i[286];
  assign N1108 = N1107 | N1102;
  assign N1109 = commit_instr_i[285] | N1108;
  assign N1110 = N1099 | N1109;
  assign N1111 = ~N1110;
  assign N1112 = commit_instr_i[284] | N1109;
  assign N1113 = ~N1112;
  assign N1114 = commit_instr_i[293] | commit_instr_i[294];
  assign N1115 = N1091 | N1114;
  assign N1116 = commit_instr_i[291] | N1115;
  assign N1117 = ~N1116;
  assign { N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78 } = (N0)? amo_resp_i[63:0] : 
                                                                                                                                                                                                                                                                                                                                                                                        (N77)? commit_instr_i[265:202] : 1'b0;
  assign N0 = amo_resp_i[64];
  assign N148 = (N1)? commit_lsu_ready_i : 
                (N147)? 1'b1 : 1'b0;
  assign N1 = N146;
  assign N149 = (N1)? commit_lsu_ready_i : 
                (N147)? 1'b0 : 1'b0;
  assign { N163, N162, N161, N160, N159 } = (N2)? commit_instr_i[138:134] : 
                                            (N3)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N2 = N157;
  assign N3 = N158;
  assign N164 = (N4)? N149 : 
                (N5)? 1'b0 : 1'b0;
  assign N4 = N76;
  assign N5 = exception_o[0];
  assign N165 = (N4)? N148 : 
                (N5)? 1'b1 : 1'b0;
  assign { N170, N169, N168, N167, N166 } = (N4)? { N163, N162, N161, N160, N159 } : 
                                            (N5)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N171 = (N4)? N157 : 
                (N5)? 1'b0 : 1'b0;
  assign { N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } = (N6)? csr_rdata_i : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? { N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78 } : 1'b0;
  assign N6 = N1095;
  assign N7 = N1094;
  assign { N242, N241, N240, N239, N238, N237, N236 } = (N6)? commit_instr_i[290:284] : 
                                                        (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243 } = (N6)? commit_instr_i[265:202] : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N7)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N170, N169, N168, N167, N166 } : 1'b0;
  assign N307 = (N8)? no_st_pending_i : 
                (N9)? 1'b0 : 1'b0;
  assign N8 = N1111;
  assign N9 = N1110;
  assign N308 = (N8)? no_st_pending_i : 
                (N9)? N165 : 1'b0;
  assign N311 = (N10)? no_st_pending_i : 
                (N310)? N308 : 1'b0;
  assign N10 = N309;
  assign N312 = (N10)? no_st_pending_i : 
                (N310)? 1'b0 : 1'b0;
  assign N313 = (N11)? no_st_pending_i : 
                (N12)? N311 : 1'b0;
  assign N11 = N1106;
  assign N12 = N1105;
  assign N314 = (N11)? no_st_pending_i : 
                (N12)? 1'b0 : 1'b0;
  assign N315 = (N13)? N313 : 
                (N145)? 1'b0 : 1'b0;
  assign N13 = N144;
  assign N316 = (N13)? N171 : 
                (N145)? 1'b0 : 1'b0;
  assign N317 = (N13)? N76 : 
                (N145)? 1'b0 : 1'b0;
  assign N318 = (N13)? N164 : 
                (N145)? 1'b0 : 1'b0;
  assign { N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319 } = (N13)? { N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N145)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign { N389, N388, N387, N386, N385, N384, N383 } = (N13)? { N242, N241, N240, N239, N238, N237, N236 } : 
                                                        (N145)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N390 = (N13)? N1095 : 
                (N145)? 1'b0 : 1'b0;
  assign { N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391 } = (N13)? { N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N145)? { N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78 } : 1'b0;
  assign N455 = (N13)? N307 : 
                (N145)? 1'b0 : 1'b0;
  assign N456 = (N13)? N312 : 
                (N145)? 1'b0 : 1'b0;
  assign N457 = (N13)? N314 : 
                (N145)? 1'b0 : 1'b0;
  assign N460 = (N14)? amo_resp_i[64] : 
                (N459)? N315 : 1'b0;
  assign N14 = N458;
  assign N461 = (N14)? amo_resp_i[64] : 
                (N459)? 1'b0 : 1'b0;
  assign N462 = (N14)? amo_resp_i[64] : 
                (N459)? N317 : 1'b0;
  assign fence_o = (N15)? N457 : 
                   (N143)? 1'b0 : 1'b0;
  assign N15 = N142;
  assign commit_ack_o[0] = (N15)? N460 : 
                           (N143)? 1'b0 : 1'b0;
  assign N463 = (N15)? N316 : 
                (N143)? 1'b0 : 1'b0;
  assign we_gpr_o[0] = (N15)? N462 : 
                       (N143)? 1'b0 : 1'b0;
  assign commit_lsu_o = (N15)? N318 : 
                        (N143)? 1'b0 : 1'b0;
  assign { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } = (N15)? { N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N143)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign csr_op_o = (N15)? { N389, N388, N387, N386, N385, N384, N383 } : 
                    (N143)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign commit_csr_o = (N15)? N390 : 
                        (N143)? 1'b0 : 1'b0;
  assign wdata_o[63:0] = (N15)? { N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391 } : 
                         (N143)? { N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78 } : 1'b0;
  assign sfence_vma_o = (N15)? N455 : 
                        (N143)? 1'b0 : 1'b0;
  assign fence_i_o = (N15)? N456 : 
                     (N143)? 1'b0 : 1'b0;
  assign amo_valid_commit_o = (N15)? N458 : 
                              (N143)? 1'b0 : 1'b0;
  assign flush_commit_o = (N15)? N461 : 
                          (N143)? 1'b0 : 1'b0;
  assign { N564, N563, N562, N561, N560 } = (N16)? { N555, N556, N557, N558, N559 } : 
                                            (N17)? commit_instr_i[500:496] : 1'b0;
  assign N16 = N463;
  assign N17 = N554;
  assign { N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565 } = (N18)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N564, N563, N562, N561, N560 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } : 1'b0;
  assign N18 = N552;
  assign N19 = N553;
  assign N629 = (N18)? 1'b1 : 
                (N19)? N463 : 1'b0;
  assign { N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630 } = (N20)? { N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565 } : 
                                                                                                                                                                                                                                                                                                                                                                                                              (N541)? { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } : 1'b0;
  assign N20 = N540;
  assign N694 = (N20)? N629 : 
                (N541)? N463 : 1'b0;
  assign csr_wdata_o = (N21)? { N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630 } : 
                       (N532)? { N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464 } : 1'b0;
  assign N21 = N531;
  assign csr_write_fflags_o = (N21)? N694 : 
                              (N532)? N463 : 1'b0;
  assign we_gpr_o[1] = (N21)? N540 : 
                       (N532)? 1'b0 : 1'b0;
  assign commit_ack_o[1] = (N21)? N540 : 
                           (N532)? 1'b0 : 1'b0;
  assign { N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698 } = (N22)? { csr_exception_i[128:65], commit_instr_i[133:70], csr_exception_i[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N697)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N22 = N696;
  assign { N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828 } = (N23)? commit_instr_i[197:69] : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N827)? { N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698 } : 1'b0;
  assign N23 = commit_instr_i[69];
  assign { N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959 } = (N24)? { csr_exception_i[128:65], commit_instr_i[133:70], csr_exception_i[0:0] } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            (N958)? { N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828 } : 1'b0;
  assign N24 = N957;
  assign { exception_o[128:1], N1088 } = (N25)? { N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959 } : 
                                         (N695)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N25 = commit_instr_i[201];
  assign exception_o[0] = (N26)? 1'b0 : 
                          (N27)? N1088 : 1'b0;
  assign N26 = halt_i;
  assign N27 = N1089;
  assign dirty_fp_state_o = 1'b0 | 1'b0;
  assign N72 = N1158 | N1159;
  assign N1158 = N1156 | N1157;
  assign N1156 = N1154 | N1155;
  assign N1154 = N1152 | N1153;
  assign N1152 = N1150 | N1151;
  assign N1150 = N1148 | N1149;
  assign N1148 = N1146 | N1147;
  assign N1146 = N1144 | N1145;
  assign N1144 = N1142 | N1143;
  assign N1142 = N1140 | N1141;
  assign N1140 = N1138 | N1139;
  assign N1138 = N1136 | N1137;
  assign N1136 = N1134 | N1135;
  assign N1134 = N1132 | N1133;
  assign N1132 = N1130 | N1131;
  assign N1130 = N1128 | N1129;
  assign N1128 = N1126 | N1127;
  assign N1126 = N1124 | N1125;
  assign N1124 = N1122 | N1123;
  assign N1122 = N1120 | N1121;
  assign N1120 = N1118 | N1119;
  assign N1118 = ~N33;
  assign N1119 = ~N36;
  assign N1121 = ~N38;
  assign N1123 = ~N43;
  assign N1125 = ~N45;
  assign N1127 = ~N48;
  assign N1129 = ~N50;
  assign N1131 = ~N52;
  assign N1133 = ~N53;
  assign N1135 = ~N54;
  assign N1137 = ~N55;
  assign N1139 = ~N58;
  assign N1141 = ~N59;
  assign N1143 = ~N60;
  assign N1145 = ~N61;
  assign N1147 = ~N62;
  assign N1149 = ~N63;
  assign N1151 = ~N64;
  assign N1153 = ~N65;
  assign N1155 = ~N69;
  assign N1157 = ~N70;
  assign N1159 = ~N71;
  assign N73 = ~commit_instr_i[290];
  assign N74 = ~commit_instr_i[289];
  assign instr_0_is_amo = N72;
  assign N75 = ~instr_0_is_amo;
  assign N76 = ~exception_o[0];
  assign N77 = ~amo_resp_i[64];
  assign N142 = commit_instr_i[201] & N1089;
  assign N143 = ~N142;
  assign N144 = N1160 | debug_mode_i;
  assign N1160 = ~debug_req_i;
  assign N145 = ~N144;
  assign N146 = N1117 & N75;
  assign N147 = ~N146;
  assign N150 = ~commit_instr_i[291];
  assign N153 = ~commit_instr_i[294];
  assign N157 = N1161 | N1162;
  assign N1161 = ~N152;
  assign N1162 = ~N156;
  assign N158 = ~N157;
  assign N309 = N1113 | N1163;
  assign N1163 = flush_dcache_i & N1116;
  assign N310 = ~N309;
  assign N458 = instr_0_is_amo & N1164;
  assign N1164 = ~commit_instr_i[69];
  assign N459 = ~N458;
  assign N531 = N1170 & N1171;
  assign N1170 = N1169 & N75;
  assign N1169 = N1167 & N1168;
  assign N1167 = N1166 & N530;
  assign N1166 = N1165 & N1089;
  assign N1165 = commit_ack_o[0] & commit_instr_i[563];
  assign N1168 = ~flush_dcache_i;
  assign N1171 = ~single_step_i;
  assign N532 = ~N531;
  assign N539 = N1180 | N1181;
  assign N1180 = N1178 | N1179;
  assign N1178 = N1176 | N1177;
  assign N1176 = N1174 | N1175;
  assign N1174 = N1172 | N1173;
  assign N1172 = ~N534;
  assign N1173 = ~N536;
  assign N1175 = ~N537;
  assign N1177 = ~N538;
  assign N1179 = ~N547;
  assign N1181 = ~N551;
  assign N540 = N1183 & N539;
  assign N1183 = N76 & N1182;
  assign N1182 = ~commit_instr_i[431];
  assign N541 = ~N540;
  assign N542 = ~commit_instr_i[655];
  assign N543 = ~commit_instr_i[654];
  assign N544 = ~commit_instr_i[653];
  assign N548 = ~commit_instr_i[656];
  assign N552 = N1179 | N1181;
  assign N553 = ~N552;
  assign N554 = ~N463;
  assign N555 = commit_instr_i[138] | commit_instr_i[500];
  assign N556 = commit_instr_i[137] | commit_instr_i[499];
  assign N557 = commit_instr_i[136] | commit_instr_i[498];
  assign N558 = commit_instr_i[135] | commit_instr_i[497];
  assign N559 = commit_instr_i[134] | commit_instr_i[496];
  assign N695 = ~commit_instr_i[201];
  assign N696 = csr_exception_i[0] & N1184;
  assign N1184 = ~csr_exception_i[128];
  assign N697 = ~N696;
  assign N827 = ~commit_instr_i[69];
  assign N957 = N1187 & N1094;
  assign N1187 = N1185 & N1186;
  assign N1185 = csr_exception_i[0] & csr_exception_i[128];
  assign N1186 = ~amo_valid_commit_o;
  assign N958 = ~N957;
  assign N1089 = ~halt_i;

endmodule